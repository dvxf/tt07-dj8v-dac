magic
tech sky130A
magscale 1 2
timestamp 1717153468
<< viali >>
rect 7021 21641 7055 21675
rect 10241 21641 10275 21675
rect 12541 21641 12575 21675
rect 14105 21641 14139 21675
rect 14381 21641 14415 21675
rect 16589 21641 16623 21675
rect 20637 21641 20671 21675
rect 26709 21641 26743 21675
rect 29837 21641 29871 21675
rect 8217 21573 8251 21607
rect 8769 21573 8803 21607
rect 13553 21573 13587 21607
rect 14841 21573 14875 21607
rect 17049 21573 17083 21607
rect 18981 21573 19015 21607
rect 21557 21573 21591 21607
rect 24501 21573 24535 21607
rect 25513 21573 25547 21607
rect 26433 21573 26467 21607
rect 26893 21573 26927 21607
rect 27537 21573 27571 21607
rect 29561 21573 29595 21607
rect 1317 21505 1351 21539
rect 3617 21505 3651 21539
rect 5641 21505 5675 21539
rect 6377 21505 6411 21539
rect 7573 21505 7607 21539
rect 9413 21505 9447 21539
rect 9505 21505 9539 21539
rect 11161 21505 11195 21539
rect 29285 21505 29319 21539
rect 2697 21437 2731 21471
rect 3065 21437 3099 21471
rect 3525 21437 3559 21471
rect 6653 21437 6687 21471
rect 7849 21437 7883 21471
rect 9137 21437 9171 21471
rect 12449 21437 12483 21471
rect 12909 21437 12943 21471
rect 13737 21437 13771 21471
rect 14657 21437 14691 21471
rect 16497 21437 16531 21471
rect 16865 21437 16899 21471
rect 18705 21437 18739 21471
rect 18889 21437 18923 21471
rect 19073 21437 19107 21471
rect 19165 21437 19199 21471
rect 19349 21437 19383 21471
rect 20453 21437 20487 21471
rect 20637 21437 20671 21471
rect 21833 21437 21867 21471
rect 24041 21437 24075 21471
rect 24685 21437 24719 21471
rect 25789 21437 25823 21471
rect 26065 21437 26099 21471
rect 26617 21437 26651 21471
rect 27445 21437 27479 21471
rect 27721 21437 27755 21471
rect 28089 21437 28123 21471
rect 29009 21437 29043 21471
rect 29147 21437 29181 21471
rect 29469 21437 29503 21471
rect 29745 21437 29779 21471
rect 30021 21437 30055 21471
rect 30481 21437 30515 21471
rect 3893 21369 3927 21403
rect 7297 21369 7331 21403
rect 8493 21369 8527 21403
rect 10149 21369 10183 21403
rect 11437 21369 11471 21403
rect 11897 21369 11931 21403
rect 13093 21369 13127 21403
rect 13277 21369 13311 21403
rect 14565 21369 14599 21403
rect 24409 21369 24443 21403
rect 27169 21369 27203 21403
rect 3341 21301 3375 21335
rect 5825 21301 5859 21335
rect 6193 21301 6227 21335
rect 6285 21301 6319 21335
rect 6837 21301 6871 21335
rect 7757 21301 7791 21335
rect 8953 21301 8987 21335
rect 9597 21301 9631 21335
rect 9965 21301 9999 21335
rect 12173 21301 12207 21335
rect 13829 21301 13863 21335
rect 13921 21301 13955 21335
rect 14197 21301 14231 21335
rect 14365 21301 14399 21335
rect 21373 21301 21407 21335
rect 23949 21301 23983 21335
rect 24133 21301 24167 21335
rect 24225 21301 24259 21335
rect 25329 21301 25363 21335
rect 25881 21301 25915 21335
rect 27261 21301 27295 21335
rect 28273 21301 28307 21335
rect 29377 21301 29411 21335
rect 30297 21301 30331 21335
rect 3525 21097 3559 21131
rect 3985 21097 4019 21131
rect 4077 21097 4111 21131
rect 4629 21097 4663 21131
rect 4997 21097 5031 21131
rect 5089 21097 5123 21131
rect 6469 21097 6503 21131
rect 6837 21097 6871 21131
rect 10057 21097 10091 21131
rect 13753 21097 13787 21131
rect 13921 21097 13955 21131
rect 15761 21097 15795 21131
rect 18521 21097 18555 21131
rect 19073 21097 19107 21131
rect 19241 21097 19275 21131
rect 21557 21097 21591 21131
rect 24317 21097 24351 21131
rect 28089 21097 28123 21131
rect 30113 21097 30147 21131
rect 30849 21097 30883 21131
rect 2881 21029 2915 21063
rect 7021 21029 7055 21063
rect 8769 21029 8803 21063
rect 9597 21029 9631 21063
rect 9689 21029 9723 21063
rect 13553 21029 13587 21063
rect 16405 21029 16439 21063
rect 16681 21029 16715 21063
rect 19441 21029 19475 21063
rect 21465 21029 21499 21063
rect 27629 21029 27663 21063
rect 27721 21029 27755 21063
rect 3065 20961 3099 20995
rect 3341 20961 3375 20995
rect 5457 20961 5491 20995
rect 5825 20961 5859 20995
rect 6377 20961 6411 20995
rect 10425 20961 10459 20995
rect 10517 20961 10551 20995
rect 11345 20961 11379 20995
rect 12449 20961 12483 20995
rect 12541 20961 12575 20995
rect 13277 20961 13311 20995
rect 14197 20961 14231 20995
rect 15117 20961 15151 20995
rect 15210 20961 15244 20995
rect 15393 20961 15427 20995
rect 15485 20961 15519 20995
rect 15623 20961 15657 20995
rect 16129 20961 16163 20995
rect 16313 20961 16347 20995
rect 16497 20961 16531 20995
rect 18735 20961 18769 20995
rect 20177 20961 20211 20995
rect 20269 20961 20303 20995
rect 20361 20961 20395 20995
rect 21649 20961 21683 20995
rect 22569 20961 22603 20995
rect 22753 20961 22787 20995
rect 22845 20961 22879 20995
rect 22937 20961 22971 20995
rect 23305 20961 23339 20995
rect 23489 20961 23523 20995
rect 23581 20961 23615 20995
rect 24501 20961 24535 20995
rect 24593 20961 24627 20995
rect 24961 20961 24995 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 25421 20961 25455 20995
rect 25513 20961 25547 20995
rect 25697 20961 25731 20995
rect 25789 20961 25823 20995
rect 26525 20961 26559 20995
rect 26709 20961 26743 20995
rect 27491 20961 27525 20995
rect 27904 20961 27938 20995
rect 27997 20961 28031 20995
rect 28457 20961 28491 20995
rect 30297 20961 30331 20995
rect 30757 20961 30791 20995
rect 857 20893 891 20927
rect 1133 20893 1167 20927
rect 4169 20893 4203 20927
rect 5181 20893 5215 20927
rect 6193 20893 6227 20927
rect 9045 20893 9079 20927
rect 9873 20893 9907 20927
rect 10701 20893 10735 20927
rect 11437 20893 11471 20927
rect 11529 20893 11563 20927
rect 12633 20893 12667 20927
rect 14473 20893 14507 20927
rect 18889 20893 18923 20927
rect 18981 20893 19015 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 26617 20893 26651 20927
rect 28365 20893 28399 20927
rect 30573 20893 30607 20927
rect 3617 20825 3651 20859
rect 9229 20825 9263 20859
rect 21833 20825 21867 20859
rect 23765 20825 23799 20859
rect 25513 20825 25547 20859
rect 3249 20757 3283 20791
rect 5641 20757 5675 20791
rect 6009 20757 6043 20791
rect 10977 20757 11011 20791
rect 12081 20757 12115 20791
rect 13001 20757 13035 20791
rect 13737 20757 13771 20791
rect 19257 20757 19291 20791
rect 21281 20757 21315 20791
rect 23213 20757 23247 20791
rect 23305 20757 23339 20791
rect 27353 20757 27387 20791
rect 28273 20757 28307 20791
rect 30481 20757 30515 20791
rect 2881 20553 2915 20587
rect 8677 20553 8711 20587
rect 10517 20553 10551 20587
rect 11069 20553 11103 20587
rect 14105 20553 14139 20587
rect 15577 20553 15611 20587
rect 16313 20553 16347 20587
rect 17877 20553 17911 20587
rect 22661 20553 22695 20587
rect 24685 20553 24719 20587
rect 24777 20553 24811 20587
rect 29377 20553 29411 20587
rect 29469 20553 29503 20587
rect 31125 20553 31159 20587
rect 8953 20485 8987 20519
rect 16865 20485 16899 20519
rect 17693 20485 17727 20519
rect 20361 20485 20395 20519
rect 30573 20485 30607 20519
rect 1869 20417 1903 20451
rect 2605 20417 2639 20451
rect 3249 20417 3283 20451
rect 5273 20417 5307 20451
rect 7297 20417 7331 20451
rect 7849 20417 7883 20451
rect 9597 20417 9631 20451
rect 9965 20417 9999 20451
rect 10057 20417 10091 20451
rect 11391 20417 11425 20451
rect 15761 20417 15795 20451
rect 17233 20417 17267 20451
rect 17509 20417 17543 20451
rect 22569 20417 22603 20451
rect 24869 20417 24903 20451
rect 27629 20417 27663 20451
rect 949 20349 983 20383
rect 1593 20349 1627 20383
rect 1685 20349 1719 20383
rect 3065 20349 3099 20383
rect 7573 20349 7607 20383
rect 8769 20349 8803 20383
rect 11161 20349 11195 20383
rect 12817 20349 12851 20383
rect 13185 20349 13219 20383
rect 13553 20349 13587 20383
rect 14289 20349 14323 20383
rect 14381 20349 14415 20383
rect 14749 20349 14783 20383
rect 14841 20349 14875 20383
rect 15025 20349 15059 20383
rect 15485 20349 15519 20383
rect 15669 20349 15703 20383
rect 15945 20349 15979 20383
rect 16405 20349 16439 20383
rect 16589 20349 16623 20383
rect 16773 20349 16807 20383
rect 16957 20349 16991 20383
rect 17325 20349 17359 20383
rect 17417 20349 17451 20383
rect 20177 20349 20211 20383
rect 20269 20349 20303 20383
rect 20453 20349 20487 20383
rect 21189 20349 21223 20383
rect 21281 20349 21315 20383
rect 21373 20349 21407 20383
rect 21557 20349 21591 20383
rect 22477 20349 22511 20383
rect 24594 20327 24628 20361
rect 27167 20349 27201 20383
rect 27491 20349 27525 20383
rect 29009 20323 29043 20357
rect 29469 20349 29503 20383
rect 30573 20349 30607 20383
rect 30757 20349 30791 20383
rect 31033 20349 31067 20383
rect 31217 20349 31251 20383
rect 2421 20281 2455 20315
rect 3525 20281 3559 20315
rect 5549 20281 5583 20315
rect 8125 20281 8159 20315
rect 9321 20281 9355 20315
rect 13645 20281 13679 20315
rect 17861 20281 17895 20315
rect 18061 20281 18095 20315
rect 20913 20281 20947 20315
rect 22201 20281 22235 20315
rect 29219 20281 29253 20315
rect 29745 20281 29779 20315
rect 1133 20213 1167 20247
rect 1225 20213 1259 20247
rect 2053 20213 2087 20247
rect 2513 20213 2547 20247
rect 9413 20213 9447 20247
rect 10149 20213 10183 20247
rect 14565 20213 14599 20247
rect 14657 20213 14691 20247
rect 14841 20213 14875 20247
rect 16037 20213 16071 20247
rect 16129 20213 16163 20247
rect 16497 20213 16531 20247
rect 17049 20213 17083 20247
rect 19993 20213 20027 20247
rect 22293 20213 22327 20247
rect 26985 20213 27019 20247
rect 27169 20213 27203 20247
rect 29101 20213 29135 20247
rect 29837 20213 29871 20247
rect 10425 20009 10459 20043
rect 12541 20009 12575 20043
rect 17969 20009 18003 20043
rect 25145 20009 25179 20043
rect 27077 20009 27111 20043
rect 1225 19941 1259 19975
rect 2973 19941 3007 19975
rect 6193 19941 6227 19975
rect 22937 19941 22971 19975
rect 23029 19941 23063 19975
rect 24133 19941 24167 19975
rect 24501 19941 24535 19975
rect 30665 19941 30699 19975
rect 3617 19873 3651 19907
rect 5917 19873 5951 19907
rect 8033 19873 8067 19907
rect 10241 19873 10275 19907
rect 10701 19873 10735 19907
rect 11345 19873 11379 19907
rect 11897 19873 11931 19907
rect 12265 19873 12299 19907
rect 12449 19873 12483 19907
rect 17601 19873 17635 19907
rect 18277 19873 18311 19907
rect 18613 19873 18647 19907
rect 18797 19873 18831 19907
rect 18889 19873 18923 19907
rect 18981 19873 19015 19907
rect 19625 19873 19659 19907
rect 19901 19873 19935 19907
rect 20085 19873 20119 19907
rect 22385 19873 22419 19907
rect 23397 19873 23431 19907
rect 23673 19873 23707 19907
rect 23857 19873 23891 19907
rect 24317 19873 24351 19907
rect 24593 19873 24627 19907
rect 24777 19873 24811 19907
rect 24961 19873 24995 19907
rect 25237 19873 25271 19907
rect 25329 19873 25363 19907
rect 26433 19873 26467 19907
rect 26617 19873 26651 19907
rect 26893 19873 26927 19907
rect 27905 19873 27939 19907
rect 28089 19873 28123 19907
rect 28181 19873 28215 19907
rect 30389 19873 30423 19907
rect 30481 19873 30515 19907
rect 949 19805 983 19839
rect 3985 19805 4019 19839
rect 7941 19805 7975 19839
rect 8309 19805 8343 19839
rect 11437 19805 11471 19839
rect 11529 19805 11563 19839
rect 17693 19805 17727 19839
rect 18061 19805 18095 19839
rect 18521 19805 18555 19839
rect 22108 19805 22142 19839
rect 22201 19805 22235 19839
rect 22293 19805 22327 19839
rect 22569 19805 22603 19839
rect 22661 19805 22695 19839
rect 23146 19805 23180 19839
rect 24869 19805 24903 19839
rect 26801 19805 26835 19839
rect 9781 19737 9815 19771
rect 19717 19737 19751 19771
rect 19809 19737 19843 19771
rect 23305 19737 23339 19771
rect 26709 19737 26743 19771
rect 27997 19737 28031 19771
rect 5411 19669 5445 19703
rect 10057 19669 10091 19703
rect 10977 19669 11011 19703
rect 17601 19669 17635 19703
rect 18153 19669 18187 19703
rect 19257 19669 19291 19703
rect 19349 19669 19383 19703
rect 23581 19669 23615 19703
rect 24041 19669 24075 19703
rect 27721 19669 27755 19703
rect 3065 19465 3099 19499
rect 3433 19465 3467 19499
rect 10149 19465 10183 19499
rect 10701 19465 10735 19499
rect 14289 19465 14323 19499
rect 14565 19465 14599 19499
rect 14657 19465 14691 19499
rect 15301 19465 15335 19499
rect 16221 19465 16255 19499
rect 18981 19465 19015 19499
rect 19165 19465 19199 19499
rect 19349 19465 19383 19499
rect 24409 19465 24443 19499
rect 24869 19465 24903 19499
rect 26157 19465 26191 19499
rect 26709 19465 26743 19499
rect 29929 19465 29963 19499
rect 30849 19465 30883 19499
rect 6101 19397 6135 19431
rect 7941 19397 7975 19431
rect 9597 19397 9631 19431
rect 13185 19397 13219 19431
rect 29009 19397 29043 19431
rect 857 19329 891 19363
rect 4169 19329 4203 19363
rect 4353 19329 4387 19363
rect 4721 19329 4755 19363
rect 5549 19329 5583 19363
rect 6837 19329 6871 19363
rect 8585 19329 8619 19363
rect 14841 19329 14875 19363
rect 16405 19329 16439 19363
rect 21465 19329 21499 19363
rect 21649 19329 21683 19363
rect 21925 19329 21959 19363
rect 22293 19329 22327 19363
rect 22385 19329 22419 19363
rect 23121 19329 23155 19363
rect 2881 19261 2915 19295
rect 8125 19261 8159 19295
rect 8769 19261 8803 19295
rect 10793 19261 10827 19295
rect 11437 19261 11471 19295
rect 11529 19261 11563 19295
rect 11897 19261 11931 19295
rect 12449 19261 12483 19295
rect 12725 19261 12759 19295
rect 13001 19261 13035 19295
rect 13185 19261 13219 19295
rect 13921 19261 13955 19295
rect 14013 19261 14047 19295
rect 14381 19261 14415 19295
rect 14933 19261 14967 19295
rect 15025 19261 15059 19295
rect 15117 19261 15151 19295
rect 15485 19261 15519 19295
rect 15577 19261 15611 19295
rect 15669 19261 15703 19295
rect 15761 19261 15795 19295
rect 16497 19261 16531 19295
rect 16589 19261 16623 19295
rect 16681 19261 16715 19295
rect 16957 19261 16991 19295
rect 17049 19261 17083 19295
rect 17233 19261 17267 19295
rect 17325 19261 17359 19295
rect 17417 19261 17451 19295
rect 19257 19261 19291 19295
rect 19441 19261 19475 19295
rect 20269 19261 20303 19295
rect 20361 19261 20395 19295
rect 20453 19261 20487 19295
rect 20545 19261 20579 19295
rect 20730 19239 20764 19273
rect 20821 19261 20855 19295
rect 21005 19261 21039 19295
rect 21189 19261 21223 19295
rect 21741 19261 21775 19295
rect 21833 19261 21867 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 23029 19261 23063 19295
rect 23489 19261 23523 19295
rect 23857 19261 23891 19295
rect 24041 19261 24075 19295
rect 24593 19261 24627 19295
rect 24685 19261 24719 19295
rect 24961 19261 24995 19295
rect 26341 19261 26375 19295
rect 26433 19261 26467 19295
rect 26893 19261 26927 19295
rect 27169 19261 27203 19295
rect 29193 19261 29227 19295
rect 29285 19261 29319 19295
rect 29377 19261 29411 19295
rect 29469 19261 29503 19295
rect 29653 19261 29687 19295
rect 30113 19261 30147 19295
rect 30382 19261 30416 19295
rect 30490 19261 30524 19295
rect 1133 19193 1167 19227
rect 3249 19193 3283 19227
rect 6653 19193 6687 19227
rect 7573 19193 7607 19227
rect 9321 19193 9355 19227
rect 9873 19193 9907 19227
rect 11621 19193 11655 19227
rect 11759 19193 11793 19227
rect 12265 19193 12299 19227
rect 12633 19193 12667 19227
rect 18797 19193 18831 19227
rect 21097 19193 21131 19227
rect 26157 19193 26191 19227
rect 27077 19193 27111 19227
rect 30817 19193 30851 19227
rect 31033 19193 31067 19227
rect 2605 19125 2639 19159
rect 3449 19125 3483 19159
rect 3617 19125 3651 19159
rect 3709 19125 3743 19159
rect 4077 19125 4111 19159
rect 4813 19125 4847 19159
rect 4905 19125 4939 19159
rect 5273 19125 5307 19159
rect 5641 19125 5675 19159
rect 5733 19125 5767 19159
rect 6285 19125 6319 19159
rect 6745 19125 6779 19159
rect 7481 19125 7515 19159
rect 8677 19125 8711 19159
rect 9137 19125 9171 19159
rect 11253 19125 11287 19159
rect 17601 19125 17635 19159
rect 19007 19125 19041 19159
rect 20085 19125 20119 19159
rect 21373 19125 21407 19159
rect 22109 19125 22143 19159
rect 22845 19125 22879 19159
rect 23213 19125 23247 19159
rect 23397 19125 23431 19159
rect 23857 19125 23891 19159
rect 26617 19125 26651 19159
rect 30665 19125 30699 19159
rect 1225 18921 1259 18955
rect 1501 18921 1535 18955
rect 3157 18921 3191 18955
rect 3985 18921 4019 18955
rect 4353 18921 4387 18955
rect 4813 18921 4847 18955
rect 8493 18921 8527 18955
rect 10057 18921 10091 18955
rect 17601 18921 17635 18955
rect 17785 18921 17819 18955
rect 22477 18921 22511 18955
rect 22937 18921 22971 18955
rect 24777 18921 24811 18955
rect 26893 18921 26927 18955
rect 29377 18921 29411 18955
rect 1869 18853 1903 18887
rect 3617 18853 3651 18887
rect 5181 18853 5215 18887
rect 6193 18853 6227 18887
rect 8953 18853 8987 18887
rect 9597 18853 9631 18887
rect 11529 18853 11563 18887
rect 21741 18853 21775 18887
rect 949 18785 983 18819
rect 1409 18785 1443 18819
rect 2697 18785 2731 18819
rect 3525 18785 3559 18819
rect 4445 18785 4479 18819
rect 5825 18785 5859 18819
rect 6009 18785 6043 18819
rect 8401 18785 8435 18819
rect 8861 18785 8895 18819
rect 9689 18785 9723 18819
rect 11253 18785 11287 18819
rect 11621 18785 11655 18819
rect 11805 18785 11839 18819
rect 13645 18785 13679 18819
rect 13737 18785 13771 18819
rect 13921 18785 13955 18819
rect 16957 18785 16991 18819
rect 17141 18785 17175 18819
rect 17233 18785 17267 18819
rect 17325 18785 17359 18819
rect 17969 18785 18003 18819
rect 19073 18785 19107 18819
rect 19257 18785 19291 18819
rect 19349 18785 19383 18819
rect 19441 18785 19475 18819
rect 19993 18785 20027 18819
rect 20085 18785 20119 18819
rect 20453 18785 20487 18819
rect 20545 18785 20579 18819
rect 21649 18785 21683 18819
rect 21833 18785 21867 18819
rect 22109 18785 22143 18819
rect 22753 18785 22787 18819
rect 26709 18785 26743 18819
rect 26893 18785 26927 18819
rect 26985 18785 27019 18819
rect 27077 18785 27111 18819
rect 28917 18785 28951 18819
rect 29009 18785 29043 18819
rect 29193 18785 29227 18819
rect 1961 18717 1995 18751
rect 2145 18717 2179 18751
rect 2513 18717 2547 18751
rect 2605 18717 2639 18751
rect 3801 18717 3835 18751
rect 4537 18717 4571 18751
rect 5273 18717 5307 18751
rect 5457 18717 5491 18751
rect 8125 18717 8159 18751
rect 9045 18717 9079 18751
rect 9505 18717 9539 18751
rect 10701 18717 10735 18751
rect 11437 18717 11471 18751
rect 11713 18717 11747 18751
rect 18061 18717 18095 18751
rect 18153 18717 18187 18751
rect 18245 18717 18279 18751
rect 20177 18717 20211 18751
rect 20269 18717 20303 18751
rect 20637 18717 20671 18751
rect 22017 18717 22051 18751
rect 22201 18717 22235 18751
rect 22293 18717 22327 18751
rect 22569 18717 22603 18751
rect 24961 18717 24995 18751
rect 25053 18717 25087 18751
rect 25145 18717 25179 18751
rect 25237 18717 25271 18751
rect 27261 18717 27295 18751
rect 5825 18649 5859 18683
rect 11069 18649 11103 18683
rect 19717 18649 19751 18683
rect 20913 18649 20947 18683
rect 27169 18649 27203 18683
rect 29101 18649 29135 18683
rect 1133 18581 1167 18615
rect 3065 18581 3099 18615
rect 6469 18581 6503 18615
rect 6653 18581 6687 18615
rect 10149 18581 10183 18615
rect 11529 18581 11563 18615
rect 19809 18581 19843 18615
rect 20545 18581 20579 18615
rect 2789 18377 2823 18411
rect 3801 18377 3835 18411
rect 5641 18377 5675 18411
rect 5733 18377 5767 18411
rect 8217 18377 8251 18411
rect 10977 18377 11011 18411
rect 11253 18377 11287 18411
rect 17049 18377 17083 18411
rect 17417 18377 17451 18411
rect 19533 18377 19567 18411
rect 19625 18377 19659 18411
rect 20453 18377 20487 18411
rect 24041 18377 24075 18411
rect 24777 18377 24811 18411
rect 24961 18377 24995 18411
rect 27537 18377 27571 18411
rect 29377 18377 29411 18411
rect 2881 18309 2915 18343
rect 4169 18309 4203 18343
rect 10333 18309 10367 18343
rect 11805 18309 11839 18343
rect 14841 18309 14875 18343
rect 20821 18309 20855 18343
rect 23213 18309 23247 18343
rect 1041 18241 1075 18275
rect 1317 18241 1351 18275
rect 3525 18241 3559 18275
rect 5089 18241 5123 18275
rect 8585 18241 8619 18275
rect 12173 18241 12207 18275
rect 12265 18241 12299 18275
rect 12541 18241 12575 18275
rect 13185 18241 13219 18275
rect 14105 18241 14139 18275
rect 14381 18241 14415 18275
rect 15853 18241 15887 18275
rect 19349 18241 19383 18275
rect 19437 18241 19471 18275
rect 20453 18241 20487 18275
rect 22753 18241 22787 18275
rect 24685 18241 24719 18275
rect 25053 18241 25087 18275
rect 26709 18241 26743 18275
rect 30389 18241 30423 18275
rect 30573 18241 30607 18275
rect 3065 18173 3099 18207
rect 3433 18173 3467 18207
rect 3893 18173 3927 18207
rect 4261 18173 4295 18207
rect 5917 18173 5951 18207
rect 6009 18173 6043 18207
rect 6193 18173 6227 18207
rect 8033 18173 8067 18207
rect 8217 18173 8251 18207
rect 10609 18173 10643 18207
rect 10885 18173 10919 18207
rect 11161 18173 11195 18207
rect 11437 18173 11471 18207
rect 11621 18173 11655 18207
rect 11713 18173 11747 18207
rect 11989 18173 12023 18207
rect 12633 18173 12667 18207
rect 12909 18173 12943 18207
rect 13001 18173 13035 18207
rect 13921 18173 13955 18207
rect 14013 18173 14047 18207
rect 14197 18173 14231 18207
rect 14473 18173 14507 18207
rect 14657 18173 14691 18207
rect 14749 18173 14783 18207
rect 14933 18173 14967 18207
rect 15209 18173 15243 18207
rect 15393 18173 15427 18207
rect 15485 18173 15519 18207
rect 15577 18173 15611 18207
rect 15945 18173 15979 18207
rect 16037 18173 16071 18207
rect 16221 18173 16255 18207
rect 16865 18173 16899 18207
rect 17141 18173 17175 18207
rect 18797 18173 18831 18207
rect 18889 18173 18923 18207
rect 19073 18173 19107 18207
rect 19165 18173 19199 18207
rect 19717 18173 19751 18207
rect 20637 18173 20671 18207
rect 22661 18173 22695 18207
rect 22937 18173 22971 18207
rect 23029 18173 23063 18207
rect 23949 18173 23983 18207
rect 24409 18173 24443 18207
rect 24961 18173 24995 18207
rect 25237 18173 25271 18207
rect 30481 18173 30515 18207
rect 30665 18173 30699 18207
rect 27491 18139 27525 18173
rect 3985 18105 4019 18139
rect 4169 18105 4203 18139
rect 4445 18105 4479 18139
rect 5723 18105 5757 18139
rect 6469 18105 6503 18139
rect 8861 18105 8895 18139
rect 10793 18105 10827 18139
rect 20361 18105 20395 18139
rect 24225 18105 24259 18139
rect 26709 18105 26743 18139
rect 26801 18105 26835 18139
rect 27721 18105 27755 18139
rect 29101 18105 29135 18139
rect 4629 18037 4663 18071
rect 5181 18037 5215 18071
rect 5273 18037 5307 18071
rect 7941 18037 7975 18071
rect 10425 18037 10459 18071
rect 12725 18037 12759 18071
rect 15945 18037 15979 18071
rect 24317 18037 24351 18071
rect 26231 18037 26265 18071
rect 27353 18037 27387 18071
rect 30205 18037 30239 18071
rect 6285 17833 6319 17867
rect 7849 17833 7883 17867
rect 9965 17833 9999 17867
rect 11897 17833 11931 17867
rect 12350 17833 12384 17867
rect 16957 17833 16991 17867
rect 17325 17833 17359 17867
rect 17877 17833 17911 17867
rect 19809 17833 19843 17867
rect 23965 17833 23999 17867
rect 24133 17833 24167 17867
rect 25145 17833 25179 17867
rect 28917 17833 28951 17867
rect 29929 17833 29963 17867
rect 6653 17765 6687 17799
rect 8201 17765 8235 17799
rect 8401 17765 8435 17799
rect 8861 17765 8895 17799
rect 9505 17765 9539 17799
rect 10333 17765 10367 17799
rect 11129 17765 11163 17799
rect 11345 17765 11379 17799
rect 12265 17765 12299 17799
rect 19441 17765 19475 17799
rect 19533 17765 19567 17799
rect 20177 17765 20211 17799
rect 21649 17765 21683 17799
rect 23765 17765 23799 17799
rect 24225 17765 24259 17799
rect 24409 17765 24443 17799
rect 24685 17765 24719 17799
rect 28549 17765 28583 17799
rect 29101 17765 29135 17799
rect 29285 17765 29319 17799
rect 857 17697 891 17731
rect 2697 17697 2731 17731
rect 4813 17697 4847 17731
rect 4905 17697 4939 17731
rect 5089 17697 5123 17731
rect 6101 17697 6135 17731
rect 6745 17697 6779 17731
rect 7389 17697 7423 17731
rect 7481 17697 7515 17731
rect 8493 17697 8527 17731
rect 8586 17697 8620 17731
rect 8769 17697 8803 17731
rect 8999 17697 9033 17731
rect 9229 17697 9263 17731
rect 9322 17697 9356 17731
rect 9597 17697 9631 17731
rect 9694 17697 9728 17731
rect 10144 17697 10178 17731
rect 10241 17697 10275 17731
rect 10516 17697 10550 17731
rect 10609 17697 10643 17731
rect 11713 17697 11747 17731
rect 11805 17697 11839 17731
rect 12081 17697 12115 17731
rect 12173 17697 12207 17731
rect 12449 17697 12483 17731
rect 17233 17697 17267 17731
rect 17417 17697 17451 17731
rect 17601 17697 17635 17731
rect 17693 17697 17727 17731
rect 17969 17697 18003 17731
rect 18153 17697 18187 17731
rect 19165 17697 19199 17731
rect 19257 17697 19291 17731
rect 19625 17697 19659 17731
rect 19901 17697 19935 17731
rect 19993 17697 20027 17731
rect 21465 17697 21499 17731
rect 21557 17697 21591 17731
rect 21833 17697 21867 17731
rect 21925 17697 21959 17731
rect 24501 17697 24535 17731
rect 24593 17697 24627 17731
rect 24869 17697 24903 17731
rect 25697 17697 25731 17731
rect 25973 17697 26007 17731
rect 26617 17697 26651 17731
rect 28365 17697 28399 17731
rect 28641 17697 28675 17731
rect 28733 17697 28767 17731
rect 29009 17697 29043 17731
rect 30205 17697 30239 17731
rect 30297 17697 30331 17731
rect 30389 17697 30423 17731
rect 30573 17697 30607 17731
rect 1133 17629 1167 17663
rect 2973 17629 3007 17663
rect 5549 17629 5583 17663
rect 6837 17629 6871 17663
rect 7297 17629 7331 17663
rect 25145 17629 25179 17663
rect 25513 17629 25547 17663
rect 26893 17629 26927 17663
rect 9137 17561 9171 17595
rect 11529 17561 11563 17595
rect 12081 17561 12115 17595
rect 20177 17561 20211 17595
rect 24225 17561 24259 17595
rect 24961 17561 24995 17595
rect 25789 17561 25823 17595
rect 25881 17561 25915 17595
rect 26433 17561 26467 17595
rect 29285 17561 29319 17595
rect 2605 17493 2639 17527
rect 4445 17493 4479 17527
rect 5917 17493 5951 17527
rect 8033 17493 8067 17527
rect 8217 17493 8251 17527
rect 9873 17493 9907 17527
rect 10977 17493 11011 17527
rect 11161 17493 11195 17527
rect 21281 17493 21315 17527
rect 23949 17493 23983 17527
rect 26801 17493 26835 17527
rect 1225 17289 1259 17323
rect 3249 17289 3283 17323
rect 4905 17289 4939 17323
rect 5365 17289 5399 17323
rect 5812 17289 5846 17323
rect 8125 17289 8159 17323
rect 8769 17289 8803 17323
rect 8861 17289 8895 17323
rect 9689 17289 9723 17323
rect 14381 17289 14415 17323
rect 16129 17289 16163 17323
rect 17049 17289 17083 17323
rect 19073 17289 19107 17323
rect 19257 17289 19291 17323
rect 20913 17289 20947 17323
rect 27077 17289 27111 17323
rect 27813 17289 27847 17323
rect 30757 17289 30791 17323
rect 22293 17221 22327 17255
rect 25329 17221 25363 17255
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 4077 17153 4111 17187
rect 7573 17153 7607 17187
rect 9229 17153 9263 17187
rect 10517 17153 10551 17187
rect 14473 17153 14507 17187
rect 17417 17153 17451 17187
rect 18797 17153 18831 17187
rect 21005 17153 21039 17187
rect 1409 17085 1443 17119
rect 2697 17085 2731 17119
rect 3433 17085 3467 17119
rect 4353 17085 4387 17119
rect 4721 17085 4755 17119
rect 5089 17085 5123 17119
rect 5549 17085 5583 17119
rect 8401 17085 8435 17119
rect 9045 17085 9079 17119
rect 9321 17085 9355 17119
rect 9413 17085 9447 17119
rect 9597 17085 9631 17119
rect 9873 17085 9907 17119
rect 10057 17085 10091 17119
rect 10149 17085 10183 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 11161 17085 11195 17119
rect 11345 17085 11379 17119
rect 11713 17085 11747 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 12725 17085 12759 17119
rect 13093 17085 13127 17119
rect 13185 17085 13219 17119
rect 13737 17085 13771 17119
rect 13830 17085 13864 17119
rect 14013 17085 14047 17119
rect 14243 17085 14277 17119
rect 14657 17085 14691 17119
rect 14933 17085 14967 17119
rect 15485 17085 15519 17119
rect 15648 17085 15682 17119
rect 15764 17085 15798 17119
rect 15899 17085 15933 17119
rect 17233 17085 17267 17119
rect 17325 17085 17359 17119
rect 17509 17085 17543 17119
rect 18061 17085 18095 17119
rect 18245 17085 18279 17119
rect 18705 17095 18739 17129
rect 18889 17085 18923 17119
rect 20729 17085 20763 17119
rect 20821 17085 20855 17119
rect 21649 17085 21683 17119
rect 22109 17085 22143 17119
rect 22201 17085 22235 17119
rect 22385 17085 22419 17119
rect 26434 17085 26468 17119
rect 26525 17085 26559 17119
rect 26709 17085 26743 17119
rect 26893 17085 26927 17119
rect 27261 17095 27295 17129
rect 27353 17085 27387 17119
rect 27537 17085 27571 17119
rect 27629 17085 27663 17119
rect 27905 17085 27939 17119
rect 28089 17085 28123 17119
rect 30113 17085 30147 17119
rect 30206 17085 30240 17119
rect 30578 17085 30612 17119
rect 1869 17017 1903 17051
rect 3985 17017 4019 17051
rect 4537 17017 4571 17051
rect 4629 17017 4663 17051
rect 7665 17017 7699 17051
rect 8585 17017 8619 17051
rect 10701 17017 10735 17051
rect 10885 17017 10919 17051
rect 10977 17017 11011 17051
rect 11989 17017 12023 17051
rect 12817 17017 12851 17051
rect 12909 17017 12943 17051
rect 14105 17017 14139 17051
rect 19241 17017 19275 17051
rect 19441 17017 19475 17051
rect 21097 17017 21131 17051
rect 21281 17017 21315 17051
rect 25145 17017 25179 17051
rect 26801 17017 26835 17051
rect 27997 17017 28031 17051
rect 30389 17017 30423 17051
rect 30481 17017 30515 17051
rect 1501 16949 1535 16983
rect 1961 16949 1995 16983
rect 2605 16949 2639 16983
rect 3065 16949 3099 16983
rect 3525 16949 3559 16983
rect 3893 16949 3927 16983
rect 7297 16949 7331 16983
rect 7757 16949 7791 16983
rect 11529 16949 11563 16983
rect 12357 16949 12391 16983
rect 12541 16949 12575 16983
rect 14841 16949 14875 16983
rect 18061 16949 18095 16983
rect 21373 16949 21407 16983
rect 21465 16949 21499 16983
rect 21925 16949 21959 16983
rect 7665 16745 7699 16779
rect 10149 16745 10183 16779
rect 14381 16745 14415 16779
rect 19717 16745 19751 16779
rect 20177 16745 20211 16779
rect 25329 16745 25363 16779
rect 26433 16745 26467 16779
rect 27169 16745 27203 16779
rect 28181 16745 28215 16779
rect 5273 16677 5307 16711
rect 16589 16677 16623 16711
rect 22385 16677 22419 16711
rect 24409 16677 24443 16711
rect 24961 16677 24995 16711
rect 25145 16677 25179 16711
rect 25697 16677 25731 16711
rect 857 16609 891 16643
rect 3065 16609 3099 16643
rect 4905 16609 4939 16643
rect 5457 16609 5491 16643
rect 8033 16609 8067 16643
rect 8125 16609 8159 16643
rect 9505 16609 9539 16643
rect 9873 16609 9907 16643
rect 10057 16609 10091 16643
rect 10328 16609 10362 16643
rect 10425 16609 10459 16643
rect 10517 16609 10551 16643
rect 10645 16609 10679 16643
rect 10793 16609 10827 16643
rect 10977 16609 11011 16643
rect 11529 16609 11563 16643
rect 11713 16609 11747 16643
rect 11805 16609 11839 16643
rect 11989 16609 12023 16643
rect 12081 16609 12115 16643
rect 12357 16609 12391 16643
rect 12541 16609 12575 16643
rect 14105 16609 14139 16643
rect 14289 16609 14323 16643
rect 14565 16609 14599 16643
rect 14841 16609 14875 16643
rect 16313 16609 16347 16643
rect 16773 16609 16807 16643
rect 16957 16609 16991 16643
rect 17233 16609 17267 16643
rect 17417 16609 17451 16643
rect 19533 16609 19567 16643
rect 19809 16609 19843 16643
rect 19901 16609 19935 16643
rect 20085 16609 20119 16643
rect 20177 16609 20211 16643
rect 20361 16609 20395 16643
rect 22017 16609 22051 16643
rect 23029 16609 23063 16643
rect 23121 16609 23155 16643
rect 23213 16609 23247 16643
rect 23397 16609 23431 16643
rect 23489 16609 23523 16643
rect 24317 16599 24351 16633
rect 24501 16609 24535 16643
rect 25973 16609 26007 16643
rect 26709 16609 26743 16643
rect 26801 16609 26835 16643
rect 26893 16609 26927 16643
rect 27077 16609 27111 16643
rect 27169 16609 27203 16643
rect 27353 16609 27387 16643
rect 27997 16609 28031 16643
rect 28641 16609 28675 16643
rect 28825 16609 28859 16643
rect 29101 16609 29135 16643
rect 29285 16609 29319 16643
rect 29377 16609 29411 16643
rect 29561 16609 29595 16643
rect 1133 16541 1167 16575
rect 3341 16541 3375 16575
rect 5825 16541 5859 16575
rect 6101 16541 6135 16575
rect 7573 16541 7607 16575
rect 8217 16541 8251 16575
rect 8585 16541 8619 16575
rect 9689 16541 9723 16575
rect 9781 16541 9815 16575
rect 12725 16541 12759 16575
rect 12909 16541 12943 16575
rect 13001 16541 13035 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 16129 16541 16163 16575
rect 16681 16541 16715 16575
rect 19993 16541 20027 16575
rect 25697 16541 25731 16575
rect 5641 16473 5675 16507
rect 12449 16473 12483 16507
rect 14657 16473 14691 16507
rect 14749 16473 14783 16507
rect 19349 16473 19383 16507
rect 25513 16473 25547 16507
rect 25881 16473 25915 16507
rect 28825 16473 28859 16507
rect 28917 16473 28951 16507
rect 29193 16473 29227 16507
rect 2605 16405 2639 16439
rect 4813 16405 4847 16439
rect 9137 16405 9171 16439
rect 9321 16405 9355 16439
rect 12265 16405 12299 16439
rect 14289 16405 14323 16439
rect 16865 16405 16899 16439
rect 17417 16405 17451 16439
rect 22385 16405 22419 16439
rect 22569 16405 22603 16439
rect 22845 16405 22879 16439
rect 24685 16405 24719 16439
rect 25329 16405 25363 16439
rect 1225 16201 1259 16235
rect 7573 16201 7607 16235
rect 9321 16201 9355 16235
rect 11437 16201 11471 16235
rect 12265 16201 12299 16235
rect 14657 16201 14691 16235
rect 14841 16201 14875 16235
rect 17877 16201 17911 16235
rect 19441 16201 19475 16235
rect 21189 16201 21223 16235
rect 22937 16201 22971 16235
rect 24225 16201 24259 16235
rect 30205 16201 30239 16235
rect 30389 16201 30423 16235
rect 2329 16133 2363 16167
rect 8401 16133 8435 16167
rect 17601 16133 17635 16167
rect 19349 16133 19383 16167
rect 21649 16133 21683 16167
rect 27077 16133 27111 16167
rect 2145 16065 2179 16099
rect 2973 16065 3007 16099
rect 3985 16065 4019 16099
rect 4353 16065 4387 16099
rect 5181 16065 5215 16099
rect 5273 16065 5307 16099
rect 5825 16065 5859 16099
rect 7849 16065 7883 16099
rect 9045 16065 9079 16099
rect 9873 16065 9907 16099
rect 11345 16065 11379 16099
rect 11989 16065 12023 16099
rect 13093 16065 13127 16099
rect 13369 16065 13403 16099
rect 20085 16065 20119 16099
rect 20821 16065 20855 16099
rect 21281 16065 21315 16099
rect 22753 16065 22787 16099
rect 27537 16065 27571 16099
rect 27629 16065 27663 16099
rect 1409 15997 1443 16031
rect 1869 15997 1903 16031
rect 2697 15997 2731 16031
rect 3709 15997 3743 16031
rect 5365 15997 5399 16031
rect 8033 15997 8067 16031
rect 8217 15997 8251 16031
rect 9597 15997 9631 16031
rect 11805 15997 11839 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 14565 15997 14599 16031
rect 14749 15997 14783 16031
rect 14841 15997 14875 16031
rect 15025 15997 15059 16031
rect 17233 15997 17267 16031
rect 17417 15997 17451 16031
rect 17509 15997 17543 16031
rect 17693 15997 17727 16031
rect 18705 15997 18739 16031
rect 18889 15997 18923 16031
rect 18981 15997 19015 16031
rect 19073 15997 19107 16031
rect 19626 15975 19660 16009
rect 19717 15997 19751 16031
rect 19809 15997 19843 16031
rect 20545 15997 20579 16031
rect 20637 15997 20671 16031
rect 21465 15997 21499 16031
rect 22569 15997 22603 16031
rect 22949 15997 22983 16031
rect 24041 15997 24075 16031
rect 24133 15997 24167 16031
rect 30389 15997 30423 16031
rect 30481 15997 30515 16031
rect 1961 15929 1995 15963
rect 3801 15929 3835 15963
rect 4445 15929 4479 15963
rect 6101 15929 6135 15963
rect 9413 15929 9447 15963
rect 11897 15929 11931 15963
rect 12884 15929 12918 15963
rect 19947 15929 19981 15963
rect 21189 15929 21223 15963
rect 22661 15929 22695 15963
rect 24317 15929 24351 15963
rect 30665 15929 30699 15963
rect 1501 15861 1535 15895
rect 2789 15861 2823 15895
rect 3341 15861 3375 15895
rect 4537 15861 4571 15895
rect 4905 15861 4939 15895
rect 5733 15861 5767 15895
rect 8769 15861 8803 15895
rect 8861 15861 8895 15895
rect 12725 15861 12759 15895
rect 13001 15861 13035 15895
rect 23857 15861 23891 15895
rect 27537 15861 27571 15895
rect 1133 15657 1167 15691
rect 5181 15657 5215 15691
rect 6561 15657 6595 15691
rect 11989 15657 12023 15691
rect 12541 15657 12575 15691
rect 13645 15657 13679 15691
rect 15301 15657 15335 15691
rect 17233 15657 17267 15691
rect 18245 15657 18279 15691
rect 18337 15657 18371 15691
rect 18797 15657 18831 15691
rect 22569 15657 22603 15691
rect 24501 15657 24535 15691
rect 24961 15657 24995 15691
rect 27997 15657 28031 15691
rect 29929 15657 29963 15691
rect 1501 15589 1535 15623
rect 7297 15589 7331 15623
rect 12233 15589 12267 15623
rect 12449 15589 12483 15623
rect 16865 15589 16899 15623
rect 17081 15589 17115 15623
rect 18889 15589 18923 15623
rect 22845 15589 22879 15623
rect 24133 15589 24167 15623
rect 24225 15589 24259 15623
rect 25237 15589 25271 15623
rect 25697 15589 25731 15623
rect 27353 15589 27387 15623
rect 27629 15589 27663 15623
rect 27721 15589 27755 15623
rect 28181 15589 28215 15623
rect 949 15521 983 15555
rect 3157 15521 3191 15555
rect 6469 15521 6503 15555
rect 6653 15521 6687 15555
rect 6929 15521 6963 15555
rect 9045 15521 9079 15555
rect 9321 15521 9355 15555
rect 9689 15521 9723 15555
rect 9873 15521 9907 15555
rect 10977 15521 11011 15555
rect 11161 15521 11195 15555
rect 11621 15521 11655 15555
rect 12728 15521 12762 15555
rect 12817 15521 12851 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14197 15521 14231 15555
rect 14749 15521 14783 15555
rect 14933 15521 14967 15555
rect 15393 15521 15427 15555
rect 15577 15521 15611 15555
rect 16313 15521 16347 15555
rect 16497 15521 16531 15555
rect 16589 15521 16623 15555
rect 16773 15521 16807 15555
rect 18521 15521 18555 15555
rect 19073 15521 19107 15555
rect 19165 15521 19199 15555
rect 19262 15521 19296 15555
rect 19441 15521 19475 15555
rect 19625 15521 19659 15555
rect 20729 15521 20763 15555
rect 21005 15521 21039 15555
rect 22201 15521 22235 15555
rect 22753 15521 22787 15555
rect 22937 15521 22971 15555
rect 23857 15521 23891 15555
rect 23950 15521 23984 15555
rect 24363 15521 24397 15555
rect 25422 15543 25456 15577
rect 25789 15521 25823 15555
rect 25881 15521 25915 15555
rect 26065 15521 26099 15555
rect 26249 15521 26283 15555
rect 26617 15521 26651 15555
rect 26801 15521 26835 15555
rect 27169 15521 27203 15555
rect 27445 15521 27479 15555
rect 27813 15521 27847 15555
rect 28089 15521 28123 15555
rect 28365 15521 28399 15555
rect 29285 15521 29319 15555
rect 29377 15521 29411 15555
rect 29469 15521 29503 15555
rect 29653 15521 29687 15555
rect 30113 15521 30147 15555
rect 30205 15521 30239 15555
rect 30297 15521 30331 15555
rect 1225 15453 1259 15487
rect 3433 15453 3467 15487
rect 3709 15453 3743 15487
rect 9505 15453 9539 15487
rect 9597 15453 9631 15487
rect 10241 15453 10275 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 16129 15453 16163 15487
rect 18153 15453 18187 15487
rect 18609 15453 18643 15487
rect 18981 15453 19015 15487
rect 22293 15453 22327 15487
rect 25697 15453 25731 15487
rect 26893 15453 26927 15487
rect 26985 15453 27019 15487
rect 29009 15453 29043 15487
rect 30389 15453 30423 15487
rect 3341 15385 3375 15419
rect 9137 15385 9171 15419
rect 10977 15385 11011 15419
rect 16405 15385 16439 15419
rect 19533 15385 19567 15419
rect 20913 15385 20947 15419
rect 2973 15317 3007 15351
rect 6837 15317 6871 15351
rect 10793 15317 10827 15351
rect 12081 15317 12115 15351
rect 12265 15317 12299 15351
rect 13093 15317 13127 15351
rect 14381 15317 14415 15351
rect 15117 15317 15151 15351
rect 17049 15317 17083 15351
rect 22385 15317 22419 15351
rect 25513 15317 25547 15351
rect 28549 15317 28583 15351
rect 3341 15113 3375 15147
rect 6653 15113 6687 15147
rect 8401 15113 8435 15147
rect 10241 15113 10275 15147
rect 16129 15113 16163 15147
rect 16681 15113 16715 15147
rect 18797 15113 18831 15147
rect 19717 15113 19751 15147
rect 19901 15113 19935 15147
rect 22661 15113 22695 15147
rect 22845 15113 22879 15147
rect 25605 15113 25639 15147
rect 28273 15113 28307 15147
rect 28457 15113 28491 15147
rect 30849 15113 30883 15147
rect 12449 15045 12483 15079
rect 22937 15045 22971 15079
rect 4261 14977 4295 15011
rect 4537 14977 4571 15011
rect 8861 14977 8895 15011
rect 9045 14977 9079 15011
rect 10333 14977 10367 15011
rect 10609 14977 10643 15011
rect 12081 14977 12115 15011
rect 14841 14977 14875 15011
rect 15301 14977 15335 15011
rect 22569 14977 22603 15011
rect 24225 14977 24259 15011
rect 24777 14977 24811 15011
rect 25237 14977 25271 15011
rect 857 14909 891 14943
rect 1225 14909 1259 14943
rect 3525 14885 3559 14919
rect 4169 14909 4203 14943
rect 8769 14909 8803 14943
rect 9229 14909 9263 14943
rect 9413 14909 9447 14943
rect 9505 14909 9539 14943
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 9873 14909 9907 14943
rect 10057 14909 10091 14943
rect 12449 14909 12483 14943
rect 12817 14909 12851 14943
rect 13185 14909 13219 14943
rect 13553 14909 13587 14943
rect 13737 14909 13771 14943
rect 14013 14909 14047 14943
rect 14565 14909 14599 14943
rect 14657 14909 14691 14943
rect 15485 14909 15519 14943
rect 15669 14909 15703 14943
rect 15853 14909 15887 14943
rect 16405 14909 16439 14943
rect 20177 14909 20211 14943
rect 20361 14909 20395 14943
rect 20453 14909 20487 14943
rect 21005 14909 21039 14943
rect 21097 14909 21131 14943
rect 22385 14909 22419 14943
rect 22661 14909 22695 14943
rect 23121 14909 23155 14943
rect 23213 14909 23247 14943
rect 23305 14909 23339 14943
rect 23489 14909 23523 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 25329 14909 25363 14943
rect 25421 14909 25455 14943
rect 26801 14909 26835 14943
rect 26893 14909 26927 14943
rect 26985 14909 27019 14943
rect 30573 14909 30607 14943
rect 4813 14841 4847 14875
rect 8125 14841 8159 14875
rect 19073 14841 19107 14875
rect 19533 14841 19567 14875
rect 21281 14841 21315 14875
rect 22937 14841 22971 14875
rect 23397 14841 23431 14875
rect 28089 14841 28123 14875
rect 2651 14773 2685 14807
rect 3709 14773 3743 14807
rect 4077 14773 4111 14807
rect 6285 14773 6319 14807
rect 9321 14773 9355 14807
rect 19743 14773 19777 14807
rect 19993 14773 20027 14807
rect 21182 14773 21216 14807
rect 24501 14773 24535 14807
rect 28299 14773 28333 14807
rect 1409 14569 1443 14603
rect 1685 14569 1719 14603
rect 3249 14569 3283 14603
rect 5457 14569 5491 14603
rect 6285 14569 6319 14603
rect 7021 14569 7055 14603
rect 7389 14569 7423 14603
rect 8677 14569 8711 14603
rect 9413 14569 9447 14603
rect 10149 14569 10183 14603
rect 16221 14569 16255 14603
rect 16497 14569 16531 14603
rect 16957 14569 16991 14603
rect 18153 14569 18187 14603
rect 19349 14569 19383 14603
rect 19441 14569 19475 14603
rect 19809 14569 19843 14603
rect 21465 14569 21499 14603
rect 21925 14569 21959 14603
rect 23857 14569 23891 14603
rect 24593 14569 24627 14603
rect 25237 14569 25271 14603
rect 26617 14569 26651 14603
rect 30021 14569 30055 14603
rect 31033 14569 31067 14603
rect 7757 14501 7791 14535
rect 9873 14501 9907 14535
rect 17969 14501 18003 14535
rect 18429 14501 18463 14535
rect 24961 14501 24995 14535
rect 30757 14501 30791 14535
rect 1593 14433 1627 14467
rect 2053 14433 2087 14467
rect 2881 14433 2915 14467
rect 5181 14433 5215 14467
rect 5641 14433 5675 14467
rect 6193 14433 6227 14467
rect 6929 14433 6963 14467
rect 7849 14433 7883 14467
rect 8493 14433 8527 14467
rect 8769 14433 8803 14467
rect 8917 14433 8951 14467
rect 9045 14433 9079 14467
rect 9137 14433 9171 14467
rect 9275 14433 9309 14467
rect 11161 14433 11195 14467
rect 11345 14433 11379 14467
rect 11437 14433 11471 14467
rect 11529 14433 11563 14467
rect 11713 14433 11747 14467
rect 12173 14433 12207 14467
rect 12633 14433 12667 14467
rect 13001 14433 13035 14467
rect 13553 14433 13587 14467
rect 14657 14433 14691 14467
rect 14749 14433 14783 14467
rect 15025 14433 15059 14467
rect 15576 14433 15610 14467
rect 15669 14433 15703 14467
rect 15761 14433 15795 14467
rect 15945 14433 15979 14467
rect 16129 14433 16163 14467
rect 16313 14433 16347 14467
rect 17417 14433 17451 14467
rect 17877 14433 17911 14467
rect 18061 14433 18095 14467
rect 18337 14433 18371 14467
rect 18521 14433 18555 14467
rect 18659 14433 18693 14467
rect 19533 14433 19567 14467
rect 20545 14433 20579 14467
rect 24133 14433 24167 14467
rect 24501 14433 24535 14467
rect 24777 14433 24811 14467
rect 25145 14433 25179 14467
rect 25421 14433 25455 14467
rect 25881 14433 25915 14467
rect 25973 14433 26007 14467
rect 26249 14433 26283 14467
rect 26801 14433 26835 14467
rect 27629 14433 27663 14467
rect 27721 14433 27755 14467
rect 27905 14433 27939 14467
rect 27997 14433 28031 14467
rect 28549 14433 28583 14467
rect 28641 14433 28675 14467
rect 28825 14433 28859 14467
rect 29745 14433 29779 14467
rect 29929 14433 29963 14467
rect 30481 14433 30515 14467
rect 2145 14365 2179 14399
rect 2237 14365 2271 14399
rect 2697 14365 2731 14399
rect 2789 14365 2823 14399
rect 4905 14365 4939 14399
rect 6377 14365 6411 14399
rect 6837 14365 6871 14399
rect 7665 14365 7699 14399
rect 8309 14365 8343 14399
rect 10701 14365 10735 14399
rect 11897 14365 11931 14399
rect 12449 14365 12483 14399
rect 13093 14365 13127 14399
rect 13737 14365 13771 14399
rect 15117 14365 15151 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 17141 14365 17175 14399
rect 17233 14365 17267 14399
rect 18797 14365 18831 14399
rect 19073 14365 19107 14399
rect 19165 14365 19199 14399
rect 20637 14365 20671 14399
rect 21649 14365 21683 14399
rect 21741 14365 21775 14399
rect 22017 14365 22051 14399
rect 22109 14365 22143 14399
rect 23765 14365 23799 14399
rect 24317 14365 24351 14399
rect 26065 14365 26099 14399
rect 27077 14365 27111 14399
rect 30205 14365 30239 14399
rect 30297 14365 30331 14399
rect 30389 14365 30423 14399
rect 5825 14297 5859 14331
rect 8217 14297 8251 14331
rect 9505 14297 9539 14331
rect 12265 14297 12299 14331
rect 15301 14297 15335 14331
rect 17601 14297 17635 14331
rect 26249 14297 26283 14331
rect 3433 14229 3467 14263
rect 9873 14229 9907 14263
rect 10057 14229 10091 14263
rect 14105 14229 14139 14263
rect 20545 14229 20579 14263
rect 20913 14229 20947 14263
rect 25421 14229 25455 14263
rect 26985 14229 27019 14263
rect 27445 14229 27479 14263
rect 29837 14229 29871 14263
rect 3295 14025 3329 14059
rect 5181 14025 5215 14059
rect 10425 14025 10459 14059
rect 11516 14025 11550 14059
rect 13829 14025 13863 14059
rect 14013 14025 14047 14059
rect 14749 14025 14783 14059
rect 19809 14025 19843 14059
rect 20453 14025 20487 14059
rect 20637 14025 20671 14059
rect 20821 14025 20855 14059
rect 22661 14025 22695 14059
rect 23121 14025 23155 14059
rect 24409 14025 24443 14059
rect 27445 14025 27479 14059
rect 3065 13957 3099 13991
rect 4721 13889 4755 13923
rect 5089 13889 5123 13923
rect 5549 13889 5583 13923
rect 8033 13889 8067 13923
rect 11253 13889 11287 13923
rect 13277 13889 13311 13923
rect 14841 13889 14875 13923
rect 17969 13889 18003 13923
rect 18705 13889 18739 13923
rect 27997 13889 28031 13923
rect 857 13821 891 13855
rect 1225 13821 1259 13855
rect 2881 13821 2915 13855
rect 5365 13821 5399 13855
rect 8401 13821 8435 13855
rect 8769 13821 8803 13855
rect 9229 13821 9263 13855
rect 9505 13821 9539 13855
rect 9781 13821 9815 13855
rect 9874 13821 9908 13855
rect 10149 13821 10183 13855
rect 10287 13821 10321 13855
rect 10701 13821 10735 13855
rect 10977 13821 11011 13855
rect 13553 13821 13587 13855
rect 13737 13821 13771 13855
rect 13829 13821 13863 13855
rect 14379 13821 14413 13855
rect 16957 13821 16991 13855
rect 17049 13821 17083 13855
rect 17601 13821 17635 13855
rect 17785 13821 17819 13855
rect 18245 13821 18279 13855
rect 19349 13821 19383 13855
rect 19533 13821 19567 13855
rect 22109 13821 22143 13855
rect 22529 13821 22563 13855
rect 22845 13821 22879 13855
rect 23857 13821 23891 13855
rect 24225 13821 24259 13855
rect 24593 13821 24627 13855
rect 24869 13821 24903 13855
rect 25421 13821 25455 13855
rect 25605 13821 25639 13855
rect 25789 13821 25823 13855
rect 30205 13821 30239 13855
rect 30481 13821 30515 13855
rect 5825 13753 5859 13787
rect 7849 13753 7883 13787
rect 8677 13753 8711 13787
rect 9321 13753 9355 13787
rect 9689 13753 9723 13787
rect 10057 13753 10091 13787
rect 20177 13753 20211 13787
rect 20805 13753 20839 13787
rect 21005 13753 21039 13787
rect 22293 13753 22327 13787
rect 22385 13753 22419 13787
rect 23305 13753 23339 13787
rect 24133 13753 24167 13787
rect 25053 13753 25087 13787
rect 27813 13753 27847 13787
rect 2651 13685 2685 13719
rect 7297 13685 7331 13719
rect 7389 13685 7423 13719
rect 7757 13685 7791 13719
rect 10517 13685 10551 13719
rect 10885 13685 10919 13719
rect 14197 13685 14231 13719
rect 14381 13685 14415 13719
rect 15669 13685 15703 13719
rect 23121 13685 23155 13719
rect 24041 13685 24075 13719
rect 24685 13685 24719 13719
rect 27905 13685 27939 13719
rect 1225 13481 1259 13515
rect 1869 13481 1903 13515
rect 2237 13481 2271 13515
rect 3065 13481 3099 13515
rect 3433 13481 3467 13515
rect 6009 13481 6043 13515
rect 9305 13481 9339 13515
rect 11529 13481 11563 13515
rect 21833 13481 21867 13515
rect 22201 13481 22235 13515
rect 23857 13481 23891 13515
rect 24225 13481 24259 13515
rect 25881 13481 25915 13515
rect 27077 13481 27111 13515
rect 8677 13413 8711 13447
rect 8861 13413 8895 13447
rect 9505 13413 9539 13447
rect 9873 13413 9907 13447
rect 13737 13413 13771 13447
rect 16681 13413 16715 13447
rect 17095 13413 17129 13447
rect 18705 13413 18739 13447
rect 26801 13413 26835 13447
rect 1409 13345 1443 13379
rect 2329 13345 2363 13379
rect 3525 13345 3559 13379
rect 3893 13345 3927 13379
rect 6193 13345 6227 13379
rect 6285 13345 6319 13379
rect 6561 13345 6595 13379
rect 8401 13345 8435 13379
rect 8585 13345 8619 13379
rect 9045 13345 9079 13379
rect 9597 13345 9631 13379
rect 9735 13345 9769 13379
rect 9965 13345 9999 13379
rect 10062 13345 10096 13379
rect 10425 13345 10459 13379
rect 11069 13345 11103 13379
rect 11253 13345 11287 13379
rect 11345 13345 11379 13379
rect 14657 13345 14691 13379
rect 15025 13345 15059 13379
rect 15209 13345 15243 13379
rect 15485 13345 15519 13379
rect 16313 13345 16347 13379
rect 16405 13345 16439 13379
rect 16957 13345 16991 13379
rect 17233 13345 17267 13379
rect 17325 13345 17359 13379
rect 17417 13345 17451 13379
rect 17969 13345 18003 13379
rect 18153 13345 18187 13379
rect 18245 13345 18279 13379
rect 18337 13345 18371 13379
rect 19349 13345 19383 13379
rect 19717 13345 19751 13379
rect 19901 13345 19935 13379
rect 19993 13345 20027 13379
rect 20269 13345 20303 13379
rect 21281 13345 21315 13379
rect 21373 13345 21407 13379
rect 21557 13345 21591 13379
rect 21649 13345 21683 13379
rect 22109 13345 22143 13379
rect 22753 13345 22787 13379
rect 22937 13345 22971 13379
rect 23673 13345 23707 13379
rect 24041 13355 24075 13389
rect 24225 13345 24259 13379
rect 24777 13345 24811 13379
rect 25053 13345 25087 13379
rect 26157 13345 26191 13379
rect 26433 13345 26467 13379
rect 26525 13345 26559 13379
rect 26709 13345 26743 13379
rect 26893 13345 26927 13379
rect 27537 13345 27571 13379
rect 27905 13345 27939 13379
rect 27997 13345 28031 13379
rect 28549 13345 28583 13379
rect 29009 13345 29043 13379
rect 29469 13345 29503 13379
rect 29745 13345 29779 13379
rect 30021 13345 30055 13379
rect 30481 13345 30515 13379
rect 30665 13345 30699 13379
rect 30757 13345 30791 13379
rect 30941 13345 30975 13379
rect 31033 13345 31067 13379
rect 23121 13311 23155 13345
rect 2513 13277 2547 13311
rect 3709 13277 3743 13311
rect 4169 13277 4203 13311
rect 5641 13277 5675 13311
rect 6837 13277 6871 13311
rect 8493 13277 8527 13311
rect 11713 13277 11747 13311
rect 11989 13277 12023 13311
rect 16773 13277 16807 13311
rect 17601 13277 17635 13311
rect 19257 13277 19291 13311
rect 20545 13277 20579 13311
rect 27721 13277 27755 13311
rect 27813 13277 27847 13311
rect 28181 13277 28215 13311
rect 6469 13209 6503 13243
rect 9137 13209 9171 13243
rect 15117 13209 15151 13243
rect 18521 13209 18555 13243
rect 20085 13209 20119 13243
rect 23305 13209 23339 13243
rect 28641 13209 28675 13243
rect 8309 13141 8343 13175
rect 9321 13141 9355 13175
rect 10241 13141 10275 13175
rect 10517 13141 10551 13175
rect 11345 13141 11379 13175
rect 16129 13141 16163 13175
rect 17785 13141 17819 13175
rect 24961 13141 24995 13175
rect 3709 12937 3743 12971
rect 7205 12937 7239 12971
rect 17509 12937 17543 12971
rect 18429 12937 18463 12971
rect 19625 12937 19659 12971
rect 20453 12937 20487 12971
rect 20545 12937 20579 12971
rect 21097 12937 21131 12971
rect 21465 12937 21499 12971
rect 23305 12937 23339 12971
rect 23489 12937 23523 12971
rect 24501 12937 24535 12971
rect 24961 12937 24995 12971
rect 25145 12937 25179 12971
rect 25789 12937 25823 12971
rect 27445 12937 27479 12971
rect 27721 12937 27755 12971
rect 29929 12937 29963 12971
rect 30297 12937 30331 12971
rect 2789 12869 2823 12903
rect 9965 12869 9999 12903
rect 13093 12869 13127 12903
rect 15669 12869 15703 12903
rect 19349 12869 19383 12903
rect 20085 12869 20119 12903
rect 21005 12869 21039 12903
rect 21741 12869 21775 12903
rect 1041 12801 1075 12835
rect 4629 12801 4663 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 9045 12801 9079 12835
rect 10057 12801 10091 12835
rect 10885 12801 10919 12835
rect 11345 12801 11379 12835
rect 14473 12801 14507 12835
rect 14933 12801 14967 12835
rect 18153 12801 18187 12835
rect 20361 12801 20395 12835
rect 22937 12801 22971 12835
rect 24225 12801 24259 12835
rect 27353 12801 27387 12835
rect 27537 12801 27571 12835
rect 3525 12733 3559 12767
rect 3801 12733 3835 12767
rect 4077 12733 4111 12767
rect 4169 12733 4203 12767
rect 4721 12733 4755 12767
rect 4813 12733 4847 12767
rect 8861 12733 8895 12767
rect 9321 12733 9355 12767
rect 9469 12733 9503 12767
rect 9597 12733 9631 12767
rect 9827 12733 9861 12767
rect 10517 12733 10551 12767
rect 10701 12733 10735 12767
rect 10793 12733 10827 12767
rect 11069 12733 11103 12767
rect 14013 12733 14047 12767
rect 14197 12733 14231 12767
rect 14289 12733 14323 12767
rect 15761 12733 15795 12767
rect 18337 12733 18371 12767
rect 18521 12733 18555 12767
rect 18705 12733 18739 12767
rect 18889 12733 18923 12767
rect 18981 12733 19015 12767
rect 19107 12733 19141 12767
rect 20453 12733 20487 12767
rect 20545 12733 20579 12767
rect 20729 12733 20763 12767
rect 20821 12733 20855 12767
rect 21097 12733 21131 12767
rect 21189 12733 21223 12767
rect 21557 12733 21591 12767
rect 21741 12733 21775 12767
rect 22293 12733 22327 12767
rect 24685 12733 24719 12767
rect 25329 12733 25363 12767
rect 25605 12733 25639 12767
rect 26709 12733 26743 12767
rect 27261 12733 27295 12767
rect 27997 12733 28031 12767
rect 29929 12733 29963 12767
rect 30021 12733 30055 12767
rect 1317 12665 1351 12699
rect 3985 12665 4019 12699
rect 7021 12665 7055 12699
rect 9689 12665 9723 12699
rect 10241 12665 10275 12699
rect 10425 12665 10459 12699
rect 11253 12665 11287 12699
rect 11621 12665 11655 12699
rect 15117 12665 15151 12699
rect 15485 12665 15519 12699
rect 16037 12665 16071 12699
rect 19441 12665 19475 12699
rect 22661 12665 22695 12699
rect 23121 12665 23155 12699
rect 23949 12665 23983 12699
rect 24777 12665 24811 12699
rect 26341 12665 26375 12699
rect 26893 12665 26927 12699
rect 27721 12665 27755 12699
rect 4353 12597 4387 12631
rect 5181 12597 5215 12631
rect 6745 12597 6779 12631
rect 7573 12597 7607 12631
rect 8401 12597 8435 12631
rect 8769 12597 8803 12631
rect 15301 12597 15335 12631
rect 15393 12597 15427 12631
rect 17601 12597 17635 12631
rect 19625 12597 19659 12631
rect 19809 12597 19843 12631
rect 22109 12597 22143 12631
rect 23331 12597 23365 12631
rect 24961 12597 24995 12631
rect 25421 12597 25455 12631
rect 27905 12597 27939 12631
rect 1501 12393 1535 12427
rect 4813 12393 4847 12427
rect 6653 12393 6687 12427
rect 9229 12393 9263 12427
rect 11897 12393 11931 12427
rect 14289 12393 14323 12427
rect 16405 12393 16439 12427
rect 16773 12393 16807 12427
rect 18337 12393 18371 12427
rect 19073 12393 19107 12427
rect 22109 12393 22143 12427
rect 24409 12393 24443 12427
rect 25145 12393 25179 12427
rect 25579 12393 25613 12427
rect 2421 12325 2455 12359
rect 3985 12325 4019 12359
rect 4077 12325 4111 12359
rect 10517 12325 10551 12359
rect 15577 12325 15611 12359
rect 15793 12325 15827 12359
rect 16129 12325 16163 12359
rect 16681 12325 16715 12359
rect 18705 12325 18739 12359
rect 20545 12325 20579 12359
rect 25329 12325 25363 12359
rect 25789 12325 25823 12359
rect 1685 12257 1719 12291
rect 3801 12257 3835 12291
rect 4169 12257 4203 12291
rect 6101 12257 6135 12291
rect 6561 12257 6595 12291
rect 9413 12257 9447 12291
rect 9873 12257 9907 12291
rect 10057 12257 10091 12291
rect 10149 12257 10183 12291
rect 10242 12257 10276 12291
rect 10425 12257 10459 12291
rect 10614 12257 10648 12291
rect 11161 12257 11195 12291
rect 11345 12257 11379 12291
rect 11437 12257 11471 12291
rect 11529 12257 11563 12291
rect 11713 12257 11747 12291
rect 13645 12257 13679 12291
rect 13792 12257 13826 12291
rect 14657 12257 14691 12291
rect 15393 12257 15427 12291
rect 16273 12257 16307 12291
rect 16497 12257 16531 12291
rect 16957 12257 16991 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 17417 12257 17451 12291
rect 18061 12257 18095 12291
rect 18245 12257 18279 12291
rect 18429 12257 18463 12291
rect 18797 12257 18831 12291
rect 18889 12257 18923 12291
rect 19625 12257 19659 12291
rect 20085 12257 20119 12291
rect 20177 12257 20211 12291
rect 20361 12257 20395 12291
rect 21097 12257 21131 12291
rect 21373 12257 21407 12291
rect 21833 12257 21867 12291
rect 22293 12257 22327 12291
rect 22753 12257 22787 12291
rect 23581 12257 23615 12291
rect 23765 12257 23799 12291
rect 23857 12257 23891 12291
rect 24501 12257 24535 12291
rect 24593 12257 24627 12291
rect 24869 12257 24903 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 4629 12189 4663 12223
rect 4721 12189 4755 12223
rect 6837 12189 6871 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 9965 12189 9999 12223
rect 12173 12189 12207 12223
rect 13001 12189 13035 12223
rect 14013 12189 14047 12223
rect 17785 12189 17819 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 19717 12189 19751 12223
rect 21741 12189 21775 12223
rect 22477 12189 22511 12223
rect 23397 12189 23431 12223
rect 24133 12189 24167 12223
rect 24225 12189 24259 12223
rect 24777 12189 24811 12223
rect 27537 12189 27571 12223
rect 2053 12121 2087 12155
rect 6193 12121 6227 12155
rect 14749 12121 14783 12155
rect 15945 12121 15979 12155
rect 18521 12121 18555 12155
rect 20269 12121 20303 12155
rect 21005 12121 21039 12155
rect 22017 12121 22051 12155
rect 24041 12121 24075 12155
rect 25421 12121 25455 12155
rect 4353 12053 4387 12087
rect 5181 12053 5215 12087
rect 5917 12053 5951 12087
rect 9689 12053 9723 12087
rect 10793 12053 10827 12087
rect 12817 12053 12851 12087
rect 13553 12053 13587 12087
rect 13921 12053 13955 12087
rect 15761 12053 15795 12087
rect 17601 12053 17635 12087
rect 19901 12053 19935 12087
rect 21833 12053 21867 12087
rect 22293 12053 22327 12087
rect 22845 12053 22879 12087
rect 23581 12053 23615 12087
rect 25145 12053 25179 12087
rect 25605 12053 25639 12087
rect 26985 12053 27019 12087
rect 5043 11849 5077 11883
rect 7757 11849 7791 11883
rect 9137 11849 9171 11883
rect 9505 11849 9539 11883
rect 10977 11849 11011 11883
rect 11345 11849 11379 11883
rect 12265 11849 12299 11883
rect 13369 11849 13403 11883
rect 15301 11849 15335 11883
rect 15485 11849 15519 11883
rect 17601 11849 17635 11883
rect 17877 11849 17911 11883
rect 18337 11849 18371 11883
rect 21189 11849 21223 11883
rect 21465 11849 21499 11883
rect 23949 11849 23983 11883
rect 24593 11849 24627 11883
rect 26755 11849 26789 11883
rect 3065 11781 3099 11815
rect 7481 11781 7515 11815
rect 10517 11781 10551 11815
rect 16773 11781 16807 11815
rect 20545 11781 20579 11815
rect 20913 11781 20947 11815
rect 3249 11713 3283 11747
rect 6009 11713 6043 11747
rect 8493 11713 8527 11747
rect 11069 11713 11103 11747
rect 11805 11713 11839 11747
rect 12909 11713 12943 11747
rect 13829 11713 13863 11747
rect 16497 11713 16531 11747
rect 18705 11713 18739 11747
rect 19901 11713 19935 11747
rect 24961 11713 24995 11747
rect 27169 11713 27203 11747
rect 857 11645 891 11679
rect 2881 11645 2915 11679
rect 3617 11645 3651 11679
rect 5733 11645 5767 11679
rect 7941 11645 7975 11679
rect 8033 11645 8067 11679
rect 9229 11645 9263 11679
rect 9505 11645 9539 11679
rect 9597 11645 9631 11679
rect 9689 11645 9723 11679
rect 9873 11645 9907 11679
rect 9965 11645 9999 11679
rect 10241 11645 10275 11679
rect 10425 11645 10459 11679
rect 10517 11645 10551 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 11161 11645 11195 11679
rect 11529 11645 11563 11679
rect 11713 11645 11747 11679
rect 11897 11645 11931 11679
rect 12081 11645 12115 11679
rect 12633 11645 12667 11679
rect 12817 11645 12851 11679
rect 13001 11645 13035 11679
rect 13185 11645 13219 11679
rect 13553 11645 13587 11679
rect 16313 11645 16347 11679
rect 16589 11645 16623 11679
rect 17049 11645 17083 11679
rect 17325 11645 17359 11679
rect 17785 11645 17819 11679
rect 17969 11645 18003 11679
rect 18521 11645 18555 11679
rect 18981 11645 19015 11679
rect 19073 11645 19107 11679
rect 19993 11645 20027 11679
rect 20361 11645 20395 11679
rect 20729 11645 20763 11679
rect 20821 11645 20855 11679
rect 20993 11645 21027 11679
rect 21373 11645 21407 11679
rect 21833 11645 21867 11679
rect 22293 11645 22327 11679
rect 22661 11645 22695 11679
rect 23213 11645 23247 11679
rect 24501 11645 24535 11679
rect 25329 11645 25363 11679
rect 26893 11645 26927 11679
rect 1133 11577 1167 11611
rect 8677 11577 8711 11611
rect 8769 11577 8803 11611
rect 10333 11577 10367 11611
rect 15761 11577 15795 11611
rect 16037 11577 16071 11611
rect 19441 11577 19475 11611
rect 24225 11577 24259 11611
rect 2605 11509 2639 11543
rect 8217 11509 8251 11543
rect 9321 11509 9355 11543
rect 10149 11509 10183 11543
rect 10701 11509 10735 11543
rect 15669 11509 15703 11543
rect 15853 11509 15887 11543
rect 16129 11509 16163 11543
rect 17233 11509 17267 11543
rect 17417 11509 17451 11543
rect 20177 11509 20211 11543
rect 20269 11509 20303 11543
rect 28641 11509 28675 11543
rect 1225 11305 1259 11339
rect 3249 11305 3283 11339
rect 9505 11305 9539 11339
rect 13737 11305 13771 11339
rect 13921 11305 13955 11339
rect 19717 11305 19751 11339
rect 20361 11305 20395 11339
rect 29745 11305 29779 11339
rect 3617 11237 3651 11271
rect 5089 11237 5123 11271
rect 5181 11237 5215 11271
rect 8861 11237 8895 11271
rect 9321 11237 9355 11271
rect 10333 11237 10367 11271
rect 10977 11237 11011 11271
rect 11253 11237 11287 11271
rect 11345 11237 11379 11271
rect 12265 11237 12299 11271
rect 14089 11237 14123 11271
rect 14289 11237 14323 11271
rect 17325 11237 17359 11271
rect 19901 11237 19935 11271
rect 26617 11237 26651 11271
rect 8631 11203 8665 11237
rect 1409 11169 1443 11203
rect 2053 11169 2087 11203
rect 2145 11169 2179 11203
rect 2513 11169 2547 11203
rect 4813 11169 4847 11203
rect 4906 11169 4940 11203
rect 5278 11169 5312 11203
rect 5825 11169 5859 11203
rect 7665 11169 7699 11203
rect 7813 11169 7847 11203
rect 7941 11169 7975 11203
rect 8033 11169 8067 11203
rect 8130 11169 8164 11203
rect 9781 11169 9815 11203
rect 10057 11169 10091 11203
rect 10150 11169 10184 11203
rect 10425 11169 10459 11203
rect 10522 11169 10556 11203
rect 11161 11169 11195 11203
rect 11529 11169 11563 11203
rect 11713 11169 11747 11203
rect 14657 11169 14691 11203
rect 14749 11169 14783 11203
rect 15577 11169 15611 11203
rect 16313 11169 16347 11203
rect 16497 11169 16531 11203
rect 16681 11169 16715 11203
rect 16865 11169 16899 11203
rect 16957 11169 16991 11203
rect 17141 11169 17175 11203
rect 17785 11169 17819 11203
rect 17877 11169 17911 11203
rect 17969 11169 18003 11203
rect 18521 11169 18555 11203
rect 18613 11169 18647 11203
rect 18981 11169 19015 11203
rect 20085 11169 20119 11203
rect 20637 11169 20671 11203
rect 21097 11169 21131 11203
rect 21465 11169 21499 11203
rect 21557 11169 21591 11203
rect 26801 11169 26835 11203
rect 27077 11169 27111 11203
rect 27445 11169 27479 11203
rect 28457 11169 28491 11203
rect 28917 11169 28951 11203
rect 29929 11169 29963 11203
rect 30021 11169 30055 11203
rect 2329 11101 2363 11135
rect 3065 11101 3099 11135
rect 3709 11101 3743 11135
rect 3893 11101 3927 11135
rect 9965 11101 9999 11135
rect 11989 11101 12023 11135
rect 14473 11101 14507 11135
rect 15485 11101 15519 11135
rect 16589 11101 16623 11135
rect 17693 11101 17727 11135
rect 18429 11101 18463 11135
rect 18705 11101 18739 11135
rect 19625 11101 19659 11135
rect 20821 11101 20855 11135
rect 23121 11101 23155 11135
rect 23397 11101 23431 11135
rect 25421 11101 25455 11135
rect 27629 11101 27663 11135
rect 28181 11101 28215 11135
rect 1685 11033 1719 11067
rect 5457 11033 5491 11067
rect 8493 11033 8527 11067
rect 8953 11033 8987 11067
rect 9597 11033 9631 11067
rect 10701 11033 10735 11067
rect 15117 11033 15151 11067
rect 15209 11033 15243 11067
rect 16129 11033 16163 11067
rect 18245 11033 18279 11067
rect 20913 11033 20947 11067
rect 6082 10965 6116 10999
rect 7573 10965 7607 10999
rect 8309 10965 8343 10999
rect 8677 10965 8711 10999
rect 9321 10965 9355 10999
rect 11897 10965 11931 10999
rect 14105 10965 14139 10999
rect 18153 10965 18187 10999
rect 20729 10965 20763 10999
rect 21373 10965 21407 10999
rect 25157 10965 25191 10999
rect 29561 10965 29595 10999
rect 30205 10965 30239 10999
rect 2651 10761 2685 10795
rect 5549 10761 5583 10795
rect 6929 10761 6963 10795
rect 13185 10761 13219 10795
rect 15025 10761 15059 10795
rect 16497 10761 16531 10795
rect 17785 10761 17819 10795
rect 18521 10761 18555 10795
rect 24225 10761 24259 10795
rect 24593 10761 24627 10795
rect 9413 10693 9447 10727
rect 17233 10693 17267 10727
rect 26525 10693 26559 10727
rect 857 10625 891 10659
rect 3801 10625 3835 10659
rect 6285 10625 6319 10659
rect 10333 10625 10367 10659
rect 10609 10625 10643 10659
rect 12357 10625 12391 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 15853 10625 15887 10659
rect 18153 10625 18187 10659
rect 20453 10625 20487 10659
rect 20729 10625 20763 10659
rect 23673 10625 23707 10659
rect 26341 10625 26375 10659
rect 1225 10557 1259 10591
rect 2973 10557 3007 10591
rect 4445 10557 4479 10591
rect 4538 10557 4572 10591
rect 4813 10557 4847 10591
rect 4910 10557 4944 10591
rect 5365 10557 5399 10591
rect 6009 10557 6043 10591
rect 8401 10557 8435 10591
rect 8494 10557 8528 10591
rect 8769 10557 8803 10591
rect 8907 10557 8941 10591
rect 10149 10557 10183 10591
rect 16129 10557 16163 10591
rect 17417 10557 17451 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 18337 10557 18371 10591
rect 18521 10557 18555 10591
rect 18705 10557 18739 10591
rect 21557 10557 21591 10591
rect 21649 10557 21683 10591
rect 28273 10557 28307 10591
rect 29377 10557 29411 10591
rect 29837 10557 29871 10591
rect 3617 10489 3651 10523
rect 4721 10489 4755 10523
rect 6101 10489 6135 10523
rect 8217 10489 8251 10523
rect 8677 10489 8711 10523
rect 9597 10489 9631 10523
rect 10885 10489 10919 10523
rect 13553 10489 13587 10523
rect 16681 10489 16715 10523
rect 23397 10489 23431 10523
rect 23949 10489 23983 10523
rect 26065 10489 26099 10523
rect 27997 10489 28031 10523
rect 29009 10489 29043 10523
rect 2789 10421 2823 10455
rect 3249 10421 3283 10455
rect 3709 10421 3743 10455
rect 5089 10421 5123 10455
rect 5641 10421 5675 10455
rect 9045 10421 9079 10455
rect 9781 10421 9815 10455
rect 10241 10421 10275 10455
rect 12817 10421 12851 10455
rect 16037 10421 16071 10455
rect 16773 10421 16807 10455
rect 20913 10421 20947 10455
rect 29653 10421 29687 10455
rect 1041 10217 1075 10251
rect 1317 10217 1351 10251
rect 1777 10217 1811 10251
rect 3985 10217 4019 10251
rect 5273 10217 5307 10251
rect 8309 10217 8343 10251
rect 10241 10217 10275 10251
rect 10977 10217 11011 10251
rect 11621 10217 11655 10251
rect 14565 10217 14599 10251
rect 14933 10217 14967 10251
rect 15025 10217 15059 10251
rect 15393 10217 15427 10251
rect 16865 10217 16899 10251
rect 17325 10217 17359 10251
rect 18889 10217 18923 10251
rect 24225 10217 24259 10251
rect 25237 10217 25271 10251
rect 25605 10217 25639 10251
rect 25697 10217 25731 10251
rect 26157 10217 26191 10251
rect 26801 10217 26835 10251
rect 27169 10217 27203 10251
rect 27445 10217 27479 10251
rect 2421 10149 2455 10183
rect 8217 10149 8251 10183
rect 9781 10149 9815 10183
rect 12173 10149 12207 10183
rect 13093 10149 13127 10183
rect 15485 10149 15519 10183
rect 15853 10149 15887 10183
rect 19073 10149 19107 10183
rect 19901 10149 19935 10183
rect 21281 10149 21315 10183
rect 23029 10149 23063 10183
rect 1225 10081 1259 10115
rect 1685 10081 1719 10115
rect 2145 10081 2179 10115
rect 4721 10081 4755 10115
rect 4905 10081 4939 10115
rect 4997 10081 5031 10115
rect 5089 10081 5123 10115
rect 6193 10081 6227 10115
rect 10057 10081 10091 10115
rect 10425 10081 10459 10115
rect 11253 10081 11287 10115
rect 11437 10081 11471 10115
rect 11805 10081 11839 10115
rect 12081 10081 12115 10115
rect 16497 10081 16531 10115
rect 17417 10081 17451 10115
rect 17509 10081 17543 10115
rect 17969 10081 18003 10115
rect 18061 10081 18095 10115
rect 18245 10081 18279 10115
rect 18429 10081 18463 10115
rect 18705 10081 18739 10115
rect 20269 10081 20303 10115
rect 20729 10081 20763 10115
rect 23305 10081 23339 10115
rect 23765 10081 23799 10115
rect 24409 10081 24443 10115
rect 24501 10081 24535 10115
rect 24593 10081 24627 10115
rect 24685 10081 24719 10115
rect 25881 10081 25915 10115
rect 25973 10081 26007 10115
rect 27261 10081 27295 10115
rect 29377 10081 29411 10115
rect 1961 10013 1995 10047
rect 3893 10013 3927 10047
rect 4537 10013 4571 10047
rect 6377 10013 6411 10047
rect 10517 10013 10551 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 12173 10013 12207 10047
rect 12817 10013 12851 10047
rect 14749 10013 14783 10047
rect 16221 10013 16255 10047
rect 16405 10013 16439 10047
rect 17785 10013 17819 10047
rect 19625 10013 19659 10047
rect 20545 10013 20579 10047
rect 20637 10013 20671 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 24961 10013 24995 10047
rect 25145 10013 25179 10047
rect 26525 10013 26559 10047
rect 26709 10013 26743 10047
rect 27629 10013 27663 10047
rect 29101 10013 29135 10047
rect 6009 9945 6043 9979
rect 17141 9945 17175 9979
rect 17693 9945 17727 9979
rect 24133 9945 24167 9979
rect 6929 9877 6963 9911
rect 12633 9877 12667 9911
rect 18337 9877 18371 9911
rect 21097 9877 21131 9911
rect 17325 9673 17359 9707
rect 18245 9673 18279 9707
rect 21189 9673 21223 9707
rect 21373 9673 21407 9707
rect 21741 9673 21775 9707
rect 6561 9605 6595 9639
rect 8401 9605 8435 9639
rect 10517 9605 10551 9639
rect 15577 9605 15611 9639
rect 16681 9605 16715 9639
rect 16773 9605 16807 9639
rect 17233 9605 17267 9639
rect 25973 9605 26007 9639
rect 857 9537 891 9571
rect 2605 9537 2639 9571
rect 3709 9537 3743 9571
rect 3893 9537 3927 9571
rect 6009 9537 6043 9571
rect 9045 9537 9079 9571
rect 9781 9537 9815 9571
rect 11989 9537 12023 9571
rect 12265 9537 12299 9571
rect 13185 9537 13219 9571
rect 13645 9537 13679 9571
rect 15945 9537 15979 9571
rect 16865 9537 16899 9571
rect 24409 9537 24443 9571
rect 27077 9537 27111 9571
rect 28089 9537 28123 9571
rect 2881 9469 2915 9503
rect 3617 9469 3651 9503
rect 4537 9469 4571 9503
rect 4685 9469 4719 9503
rect 4905 9469 4939 9503
rect 5043 9469 5077 9503
rect 6101 9469 6135 9503
rect 6837 9469 6871 9503
rect 6985 9469 7019 9503
rect 7113 9469 7147 9503
rect 7205 9469 7239 9503
rect 7343 9469 7377 9503
rect 7573 9469 7607 9503
rect 7666 9469 7700 9503
rect 8038 9469 8072 9503
rect 8769 9469 8803 9503
rect 9229 9469 9263 9503
rect 10057 9469 10091 9503
rect 12357 9469 12391 9503
rect 17417 9469 17451 9503
rect 17693 9469 17727 9503
rect 18061 9469 18095 9503
rect 18889 9469 18923 9503
rect 19073 9469 19107 9503
rect 19165 9469 19199 9503
rect 19441 9469 19475 9503
rect 21281 9469 21315 9503
rect 21925 9469 21959 9503
rect 24225 9469 24259 9503
rect 24685 9469 24719 9503
rect 25697 9469 25731 9503
rect 26157 9469 26191 9503
rect 27905 9469 27939 9503
rect 1133 9401 1167 9435
rect 4813 9401 4847 9435
rect 6193 9401 6227 9435
rect 7849 9401 7883 9435
rect 7941 9401 7975 9435
rect 8861 9401 8895 9435
rect 9413 9401 9447 9435
rect 9597 9401 9631 9435
rect 13921 9401 13955 9435
rect 16129 9401 16163 9435
rect 16313 9401 16347 9435
rect 19717 9401 19751 9435
rect 24961 9401 24995 9435
rect 25237 9401 25271 9435
rect 25421 9401 25455 9435
rect 25789 9401 25823 9435
rect 2697 9333 2731 9367
rect 3249 9333 3283 9367
rect 5181 9333 5215 9367
rect 7481 9333 7515 9367
rect 8217 9333 8251 9367
rect 9965 9333 9999 9367
rect 10425 9333 10459 9367
rect 12541 9333 12575 9367
rect 12633 9333 12667 9367
rect 13001 9333 13035 9367
rect 13093 9333 13127 9367
rect 15393 9333 15427 9367
rect 16037 9333 16071 9367
rect 17601 9333 17635 9367
rect 17877 9333 17911 9367
rect 18705 9333 18739 9367
rect 23213 9333 23247 9367
rect 23857 9333 23891 9367
rect 24317 9333 24351 9367
rect 25605 9333 25639 9367
rect 26433 9333 26467 9367
rect 26801 9333 26835 9367
rect 26893 9333 26927 9367
rect 27445 9333 27479 9367
rect 27813 9333 27847 9367
rect 1593 9129 1627 9163
rect 4721 9129 4755 9163
rect 5825 9129 5859 9163
rect 9238 9129 9272 9163
rect 9597 9129 9631 9163
rect 10517 9129 10551 9163
rect 11069 9129 11103 9163
rect 11253 9129 11287 9163
rect 12357 9129 12391 9163
rect 12725 9129 12759 9163
rect 19901 9129 19935 9163
rect 19993 9129 20027 9163
rect 20545 9129 20579 9163
rect 21281 9129 21315 9163
rect 21649 9129 21683 9163
rect 21741 9129 21775 9163
rect 24593 9129 24627 9163
rect 25605 9129 25639 9163
rect 30113 9129 30147 9163
rect 6193 9061 6227 9095
rect 7757 9061 7791 9095
rect 8401 9061 8435 9095
rect 8769 9061 8803 9095
rect 10701 9061 10735 9095
rect 11437 9061 11471 9095
rect 15761 9061 15795 9095
rect 18061 9061 18095 9095
rect 21005 9061 21039 9095
rect 23121 9061 23155 9095
rect 25513 9061 25547 9095
rect 1685 8993 1719 9027
rect 2145 8993 2179 9027
rect 4905 8993 4939 9027
rect 4997 8993 5031 9027
rect 5089 8993 5123 9027
rect 5273 8993 5307 9027
rect 5549 8993 5583 9027
rect 6837 8993 6871 9027
rect 6985 8993 7019 9027
rect 7113 8993 7147 9027
rect 7205 8993 7239 9027
rect 7302 8993 7336 9027
rect 7665 8993 7699 9027
rect 8861 8993 8895 9027
rect 10149 8993 10183 9027
rect 11713 8993 11747 9027
rect 12081 8993 12115 9027
rect 12817 8993 12851 9027
rect 13185 8993 13219 9027
rect 16221 8993 16255 9027
rect 18337 8993 18371 9027
rect 18521 8993 18555 9027
rect 19533 8993 19567 9027
rect 20177 8993 20211 9027
rect 20361 8993 20395 9027
rect 22293 8993 22327 9027
rect 22477 8993 22511 9027
rect 22845 8993 22879 9027
rect 25053 8993 25087 9027
rect 26065 8993 26099 9027
rect 1501 8925 1535 8959
rect 2421 8925 2455 8959
rect 3893 8925 3927 8959
rect 4537 8925 4571 8959
rect 6285 8925 6319 8959
rect 6377 8925 6411 8959
rect 9873 8925 9907 8959
rect 12909 8925 12943 8959
rect 13461 8925 13495 8959
rect 14933 8925 14967 8959
rect 15669 8925 15703 8959
rect 15853 8925 15887 8959
rect 16589 8925 16623 8959
rect 18797 8925 18831 8959
rect 19349 8925 19383 8959
rect 19441 8925 19475 8959
rect 20729 8925 20763 8959
rect 21833 8925 21867 8959
rect 25789 8925 25823 8959
rect 27997 8925 28031 8959
rect 28273 8925 28307 8959
rect 28365 8925 28399 8959
rect 28641 8925 28675 8959
rect 8125 8857 8159 8891
rect 9413 8857 9447 8891
rect 22753 8857 22787 8891
rect 25145 8857 25179 8891
rect 26249 8857 26283 8891
rect 2053 8789 2087 8823
rect 3985 8789 4019 8823
rect 5365 8789 5399 8823
rect 7481 8789 7515 8823
rect 9229 8789 9263 8823
rect 9781 8789 9815 8823
rect 10333 8789 10367 8823
rect 10517 8789 10551 8823
rect 11253 8789 11287 8823
rect 15301 8789 15335 8823
rect 16405 8789 16439 8823
rect 24869 8789 24903 8823
rect 26525 8789 26559 8823
rect 2697 8585 2731 8619
rect 5076 8585 5110 8619
rect 6653 8585 6687 8619
rect 7757 8585 7791 8619
rect 7941 8585 7975 8619
rect 8677 8585 8711 8619
rect 9321 8585 9355 8619
rect 9873 8585 9907 8619
rect 13185 8585 13219 8619
rect 13369 8585 13403 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 16497 8585 16531 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 19165 8585 19199 8619
rect 20269 8585 20303 8619
rect 22477 8585 22511 8619
rect 22845 8585 22879 8619
rect 23673 8585 23707 8619
rect 23949 8585 23983 8619
rect 24317 8585 24351 8619
rect 24672 8585 24706 8619
rect 26157 8585 26191 8619
rect 26433 8585 26467 8619
rect 27813 8585 27847 8619
rect 3249 8517 3283 8551
rect 6561 8517 6595 8551
rect 8493 8517 8527 8551
rect 10885 8517 10919 8551
rect 16129 8517 16163 8551
rect 18705 8517 18739 8551
rect 27445 8517 27479 8551
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 4813 8449 4847 8483
rect 7297 8449 7331 8483
rect 9689 8449 9723 8483
rect 11069 8449 11103 8483
rect 13001 8449 13035 8483
rect 14105 8449 14139 8483
rect 16405 8449 16439 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 18337 8449 18371 8483
rect 19717 8449 19751 8483
rect 19809 8449 19843 8483
rect 20729 8449 20763 8483
rect 23121 8449 23155 8483
rect 23213 8449 23247 8483
rect 24409 8449 24443 8483
rect 26985 8449 27019 8483
rect 857 8381 891 8415
rect 2881 8381 2915 8415
rect 3617 8381 3651 8415
rect 4077 8381 4111 8415
rect 4353 8381 4387 8415
rect 4445 8381 4479 8415
rect 7389 8381 7423 8415
rect 9045 8381 9079 8415
rect 9137 8381 9171 8415
rect 9965 8381 9999 8415
rect 10701 8381 10735 8415
rect 10977 8381 11011 8415
rect 13185 8381 13219 8415
rect 14381 8381 14415 8415
rect 14933 8381 14967 8415
rect 15669 8381 15703 8415
rect 15761 8381 15795 8415
rect 16497 8381 16531 8415
rect 17049 8381 17083 8415
rect 18889 8381 18923 8415
rect 22661 8381 22695 8415
rect 23862 8381 23896 8415
rect 27629 8381 27663 8415
rect 28089 8381 28123 8415
rect 1133 8313 1167 8347
rect 4261 8313 4295 8347
rect 7803 8313 7837 8347
rect 10241 8313 10275 8347
rect 11345 8313 11379 8347
rect 12909 8313 12943 8347
rect 15485 8313 15519 8347
rect 18153 8313 18187 8347
rect 18245 8313 18279 8347
rect 19901 8313 19935 8347
rect 21005 8313 21039 8347
rect 26893 8313 26927 8347
rect 26985 8313 27019 8347
rect 2605 8245 2639 8279
rect 4629 8245 4663 8279
rect 8668 8245 8702 8279
rect 9413 8245 9447 8279
rect 12817 8245 12851 8279
rect 13553 8245 13587 8279
rect 13921 8245 13955 8279
rect 14013 8245 14047 8279
rect 15209 8245 15243 8279
rect 23305 8245 23339 8279
rect 27905 8245 27939 8279
rect 4813 8041 4847 8075
rect 10701 8041 10735 8075
rect 11161 8041 11195 8075
rect 12449 8041 12483 8075
rect 25421 8041 25455 8075
rect 2237 7973 2271 8007
rect 8585 7973 8619 8007
rect 9873 7973 9907 8007
rect 9965 7973 9999 8007
rect 12541 7973 12575 8007
rect 15669 7973 15703 8007
rect 16405 7973 16439 8007
rect 19699 7973 19733 8007
rect 20177 7973 20211 8007
rect 20269 7973 20303 8007
rect 20453 7973 20487 8007
rect 20637 7973 20671 8007
rect 21465 7973 21499 8007
rect 22845 7973 22879 8007
rect 24869 7973 24903 8007
rect 1041 7905 1075 7939
rect 1317 7905 1351 7939
rect 1409 7905 1443 7939
rect 1593 7905 1627 7939
rect 1685 7905 1719 7939
rect 4905 7905 4939 7939
rect 5273 7905 5307 7939
rect 5365 7905 5399 7939
rect 6101 7905 6135 7939
rect 6193 7905 6227 7939
rect 6469 7905 6503 7939
rect 6745 7905 6779 7939
rect 6837 7905 6871 7939
rect 7021 7905 7055 7939
rect 7113 7905 7147 7939
rect 7941 7905 7975 7939
rect 8401 7905 8435 7939
rect 8493 7905 8527 7939
rect 8769 7905 8803 7939
rect 9137 7905 9171 7939
rect 9229 7905 9263 7939
rect 9689 7905 9723 7939
rect 10057 7905 10091 7939
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 11621 7905 11655 7939
rect 13645 7905 13679 7939
rect 13829 7905 13863 7939
rect 18245 7905 18279 7939
rect 18337 7905 18371 7939
rect 18521 7905 18555 7939
rect 19349 7905 19383 7939
rect 19993 7905 20027 7939
rect 21833 7905 21867 7939
rect 22385 7905 22419 7939
rect 23029 7905 23063 7939
rect 25145 7905 25179 7939
rect 25237 7905 25271 7939
rect 25421 7905 25455 7939
rect 25881 7905 25915 7939
rect 26525 7905 26559 7939
rect 28733 7905 28767 7939
rect 1961 7837 1995 7871
rect 3709 7837 3743 7871
rect 4353 7837 4387 7871
rect 5641 7837 5675 7871
rect 5917 7837 5951 7871
rect 6377 7837 6411 7871
rect 9505 7837 9539 7871
rect 11713 7837 11747 7871
rect 11897 7837 11931 7871
rect 12633 7837 12667 7871
rect 13461 7837 13495 7871
rect 16129 7837 16163 7871
rect 17877 7837 17911 7871
rect 18981 7837 19015 7871
rect 21649 7837 21683 7871
rect 22569 7837 22603 7871
rect 23397 7837 23431 7871
rect 25605 7837 25639 7871
rect 25789 7837 25823 7871
rect 26801 7837 26835 7871
rect 28273 7837 28307 7871
rect 1225 7769 1259 7803
rect 10241 7769 10275 7803
rect 12081 7769 12115 7803
rect 12909 7769 12943 7803
rect 14381 7769 14415 7803
rect 28457 7769 28491 7803
rect 1869 7701 1903 7735
rect 3801 7701 3835 7735
rect 5089 7701 5123 7735
rect 5549 7701 5583 7735
rect 6561 7701 6595 7735
rect 7389 7701 7423 7735
rect 8217 7701 8251 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 10333 7701 10367 7735
rect 11253 7701 11287 7735
rect 13737 7701 13771 7735
rect 20821 7701 20855 7735
rect 23213 7701 23247 7735
rect 26249 7701 26283 7735
rect 3249 7497 3283 7531
rect 5733 7497 5767 7531
rect 6377 7497 6411 7531
rect 6561 7497 6595 7531
rect 7021 7497 7055 7531
rect 9689 7497 9723 7531
rect 10425 7497 10459 7531
rect 11161 7497 11195 7531
rect 11529 7497 11563 7531
rect 20453 7497 20487 7531
rect 26065 7497 26099 7531
rect 2697 7429 2731 7463
rect 8493 7429 8527 7463
rect 9505 7429 9539 7463
rect 13553 7429 13587 7463
rect 15577 7429 15611 7463
rect 15761 7429 15795 7463
rect 17233 7429 17267 7463
rect 23121 7429 23155 7463
rect 25237 7429 25271 7463
rect 2605 7361 2639 7395
rect 3709 7361 3743 7395
rect 3801 7361 3835 7395
rect 7113 7361 7147 7395
rect 10149 7361 10183 7395
rect 10885 7361 10919 7395
rect 13277 7361 13311 7395
rect 13829 7361 13863 7395
rect 16129 7361 16163 7395
rect 16313 7361 16347 7395
rect 16681 7361 16715 7395
rect 18245 7361 18279 7395
rect 18705 7361 18739 7395
rect 21189 7361 21223 7395
rect 22661 7361 22695 7395
rect 25513 7361 25547 7395
rect 26801 7361 26835 7395
rect 857 7293 891 7327
rect 2881 7293 2915 7327
rect 4629 7293 4663 7327
rect 4997 7293 5031 7327
rect 5181 7293 5215 7327
rect 5549 7293 5583 7327
rect 5825 7293 5859 7327
rect 6101 7293 6135 7327
rect 6193 7293 6227 7327
rect 6745 7293 6779 7327
rect 6837 7293 6871 7327
rect 7711 7293 7745 7327
rect 7941 7293 7975 7327
rect 8069 7293 8103 7327
rect 8217 7293 8251 7327
rect 8493 7293 8527 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 9009 7293 9043 7327
rect 9326 7293 9360 7327
rect 9873 7293 9907 7327
rect 9965 7293 9999 7327
rect 10241 7293 10275 7327
rect 10609 7293 10643 7327
rect 10701 7293 10735 7327
rect 10977 7293 11011 7327
rect 11069 7293 11103 7327
rect 11161 7293 11195 7327
rect 13737 7293 13771 7327
rect 17785 7293 17819 7327
rect 18153 7293 18187 7327
rect 18337 7293 18371 7327
rect 18429 7293 18463 7327
rect 21097 7293 21131 7327
rect 21465 7293 21499 7327
rect 21925 7293 21959 7327
rect 22201 7293 22235 7327
rect 22385 7293 22419 7327
rect 22569 7293 22603 7327
rect 23489 7293 23523 7327
rect 23673 7293 23707 7327
rect 23949 7293 23983 7327
rect 24041 7293 24075 7327
rect 24152 7293 24186 7327
rect 24317 7293 24351 7327
rect 24593 7293 24627 7327
rect 24777 7293 24811 7327
rect 24869 7293 24903 7327
rect 24961 7293 24995 7327
rect 26341 7293 26375 7327
rect 26433 7293 26467 7327
rect 1133 7225 1167 7259
rect 5365 7225 5399 7259
rect 5453 7225 5487 7259
rect 6009 7225 6043 7259
rect 7297 7225 7331 7259
rect 7849 7225 7883 7259
rect 9137 7225 9171 7259
rect 9229 7225 9263 7259
rect 13001 7225 13035 7259
rect 14105 7225 14139 7259
rect 16221 7225 16255 7259
rect 17969 7225 18003 7259
rect 18981 7225 19015 7259
rect 22661 7225 22695 7259
rect 24501 7225 24535 7259
rect 26617 7225 26651 7259
rect 27077 7225 27111 7259
rect 28825 7225 28859 7259
rect 3617 7157 3651 7191
rect 4077 7157 4111 7191
rect 4813 7157 4847 7191
rect 7389 7157 7423 7191
rect 7573 7157 7607 7191
rect 11437 7157 11471 7191
rect 16773 7157 16807 7191
rect 16865 7157 16899 7191
rect 17601 7157 17635 7191
rect 22293 7157 22327 7191
rect 23581 7157 23615 7191
rect 25605 7157 25639 7191
rect 25697 7157 25731 7191
rect 26525 7157 26559 7191
rect 4629 6953 4663 6987
rect 11621 6953 11655 6987
rect 11713 6953 11747 6987
rect 12081 6953 12115 6987
rect 14749 6953 14783 6987
rect 16497 6953 16531 6987
rect 20821 6953 20855 6987
rect 25881 6953 25915 6987
rect 26617 6953 26651 6987
rect 28733 6953 28767 6987
rect 2053 6885 2087 6919
rect 8033 6885 8067 6919
rect 15393 6885 15427 6919
rect 18429 6885 18463 6919
rect 22569 6885 22603 6919
rect 22661 6885 22695 6919
rect 1041 6817 1075 6851
rect 1225 6817 1259 6851
rect 1317 6817 1351 6851
rect 1501 6817 1535 6851
rect 1593 6817 1627 6851
rect 2145 6817 2179 6851
rect 2881 6817 2915 6851
rect 3433 6817 3467 6851
rect 3617 6817 3651 6851
rect 3709 6817 3743 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 4353 6817 4387 6851
rect 4445 6817 4479 6851
rect 4721 6817 4755 6851
rect 5089 6817 5123 6851
rect 5273 6817 5307 6851
rect 5365 6817 5399 6851
rect 6193 6817 6227 6851
rect 7757 6817 7791 6851
rect 9965 6817 9999 6851
rect 10057 6817 10091 6851
rect 10609 6817 10643 6851
rect 10977 6817 11011 6851
rect 11161 6817 11195 6851
rect 12173 6817 12207 6851
rect 12541 6817 12575 6851
rect 15301 6817 15335 6851
rect 17417 6817 17451 6851
rect 17601 6817 17635 6851
rect 17969 6817 18003 6851
rect 18061 6817 18095 6851
rect 18797 6817 18831 6851
rect 19901 6817 19935 6851
rect 20085 6817 20119 6851
rect 20177 6817 20211 6851
rect 20361 6817 20395 6851
rect 21465 6817 21499 6851
rect 21833 6817 21867 6851
rect 22201 6817 22235 6851
rect 23581 6817 23615 6851
rect 24133 6817 24167 6851
rect 24225 6817 24259 6851
rect 24685 6817 24719 6851
rect 25053 6817 25087 6851
rect 26433 6817 26467 6851
rect 26709 6817 26743 6851
rect 26893 6817 26927 6851
rect 28917 6817 28951 6851
rect 29193 6817 29227 6851
rect 2329 6749 2363 6783
rect 2973 6749 3007 6783
rect 3065 6749 3099 6783
rect 5641 6749 5675 6783
rect 6837 6749 6871 6783
rect 7113 6749 7147 6783
rect 9505 6749 9539 6783
rect 10333 6749 10367 6783
rect 11069 6749 11103 6783
rect 11529 6749 11563 6783
rect 12817 6749 12851 6783
rect 14473 6749 14507 6783
rect 14657 6749 14691 6783
rect 15393 6749 15427 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 19073 6749 19107 6783
rect 19717 6749 19751 6783
rect 22661 6749 22695 6783
rect 24593 6749 24627 6783
rect 25605 6749 25639 6783
rect 25789 6749 25823 6783
rect 27169 6749 27203 6783
rect 1685 6681 1719 6715
rect 3985 6681 4019 6715
rect 4905 6681 4939 6715
rect 10793 6681 10827 6715
rect 15117 6681 15151 6715
rect 18981 6681 19015 6715
rect 20545 6681 20579 6715
rect 21465 6681 21499 6715
rect 23121 6681 23155 6715
rect 29009 6681 29043 6715
rect 2513 6613 2547 6647
rect 5549 6613 5583 6647
rect 6101 6613 6135 6647
rect 6285 6613 6319 6647
rect 7665 6613 7699 6647
rect 9781 6613 9815 6647
rect 10241 6613 10275 6647
rect 12357 6613 12391 6647
rect 14289 6613 14323 6647
rect 15853 6613 15887 6647
rect 16865 6613 16899 6647
rect 17785 6613 17819 6647
rect 18613 6613 18647 6647
rect 19349 6613 19383 6647
rect 26249 6613 26283 6647
rect 26433 6613 26467 6647
rect 28641 6613 28675 6647
rect 2651 6409 2685 6443
rect 4721 6409 4755 6443
rect 7665 6409 7699 6443
rect 8217 6409 8251 6443
rect 10609 6409 10643 6443
rect 14013 6409 14047 6443
rect 14749 6409 14783 6443
rect 16589 6409 16623 6443
rect 16773 6409 16807 6443
rect 17877 6409 17911 6443
rect 23397 6409 23431 6443
rect 3249 6341 3283 6375
rect 8401 6341 8435 6375
rect 11437 6341 11471 6375
rect 13921 6341 13955 6375
rect 15853 6341 15887 6375
rect 857 6273 891 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 5917 6273 5951 6307
rect 9045 6273 9079 6307
rect 9781 6273 9815 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11575 6273 11609 6307
rect 13369 6273 13403 6307
rect 13719 6273 13753 6307
rect 14657 6273 14691 6307
rect 15301 6273 15335 6307
rect 20085 6273 20119 6307
rect 22845 6273 22879 6307
rect 22937 6273 22971 6307
rect 24593 6273 24627 6307
rect 1225 6205 1259 6239
rect 2973 6205 3007 6239
rect 4169 6205 4203 6239
rect 4261 6205 4295 6239
rect 4445 6205 4479 6239
rect 4537 6205 4571 6239
rect 4813 6205 4847 6239
rect 5733 6205 5767 6239
rect 7757 6205 7791 6239
rect 7849 6205 7883 6239
rect 8033 6205 8067 6239
rect 9965 6205 9999 6239
rect 10058 6205 10092 6239
rect 10430 6205 10464 6239
rect 13001 6205 13035 6239
rect 13553 6205 13587 6239
rect 13829 6205 13863 6239
rect 14105 6205 14139 6239
rect 14381 6205 14415 6239
rect 16313 6205 16347 6239
rect 17601 6205 17635 6239
rect 17785 6205 17819 6239
rect 18061 6205 18095 6239
rect 18153 6205 18187 6239
rect 18429 6205 18463 6239
rect 19809 6205 19843 6239
rect 19993 6205 20027 6239
rect 20177 6205 20211 6239
rect 20361 6205 20395 6239
rect 21005 6205 21039 6239
rect 21189 6205 21223 6239
rect 21281 6205 21315 6239
rect 21373 6205 21407 6239
rect 21833 6205 21867 6239
rect 22017 6205 22051 6239
rect 24036 6205 24070 6239
rect 24408 6205 24442 6239
rect 24501 6205 24535 6239
rect 24869 6205 24903 6239
rect 24961 6205 24995 6239
rect 25053 6205 25087 6239
rect 25237 6205 25271 6239
rect 25513 6205 25547 6239
rect 25605 6205 25639 6239
rect 25697 6205 25731 6239
rect 25789 6205 25823 6239
rect 26157 6205 26191 6239
rect 26433 6205 26467 6239
rect 26709 6205 26743 6239
rect 27169 6205 27203 6239
rect 27445 6205 27479 6239
rect 28089 6205 28123 6239
rect 28641 6205 28675 6239
rect 28825 6205 28859 6239
rect 29377 6205 29411 6239
rect 3617 6137 3651 6171
rect 6193 6137 6227 6171
rect 10241 6137 10275 6171
rect 10333 6137 10367 6171
rect 11069 6137 11103 6171
rect 15393 6137 15427 6171
rect 15577 6137 15611 6171
rect 17417 6137 17451 6171
rect 18245 6137 18279 6171
rect 20269 6137 20303 6171
rect 22937 6137 22971 6171
rect 24133 6137 24167 6171
rect 24225 6137 24259 6171
rect 25973 6137 26007 6171
rect 27997 6137 28031 6171
rect 28365 6137 28399 6171
rect 2789 6069 2823 6103
rect 4997 6069 5031 6103
rect 5181 6069 5215 6103
rect 8769 6069 8803 6103
rect 8861 6069 8895 6103
rect 9229 6069 9263 6103
rect 14933 6069 14967 6103
rect 19625 6069 19659 6103
rect 20821 6069 20855 6103
rect 22661 6069 22695 6103
rect 23857 6069 23891 6103
rect 25329 6069 25363 6103
rect 26341 6069 26375 6103
rect 28733 6069 28767 6103
rect 29101 6069 29135 6103
rect 1501 5865 1535 5899
rect 4031 5865 4065 5899
rect 5365 5865 5399 5899
rect 6193 5865 6227 5899
rect 6285 5865 6319 5899
rect 6653 5865 6687 5899
rect 7113 5865 7147 5899
rect 7757 5865 7791 5899
rect 9229 5865 9263 5899
rect 9321 5865 9355 5899
rect 12817 5865 12851 5899
rect 14013 5865 14047 5899
rect 18153 5865 18187 5899
rect 19625 5865 19659 5899
rect 20177 5865 20211 5899
rect 22937 5865 22971 5899
rect 25881 5865 25915 5899
rect 28549 5865 28583 5899
rect 29009 5865 29043 5899
rect 1133 5797 1167 5831
rect 1869 5797 1903 5831
rect 8677 5797 8711 5831
rect 11253 5797 11287 5831
rect 14289 5797 14323 5831
rect 17877 5797 17911 5831
rect 18337 5797 18371 5831
rect 20453 5797 20487 5831
rect 20545 5797 20579 5831
rect 23857 5797 23891 5831
rect 25329 5797 25363 5831
rect 949 5729 983 5763
rect 1225 5729 1259 5763
rect 1317 5729 1351 5763
rect 1777 5729 1811 5763
rect 1961 5729 1995 5763
rect 2145 5729 2179 5763
rect 2237 5729 2271 5763
rect 4721 5729 4755 5763
rect 5273 5729 5307 5763
rect 7021 5729 7055 5763
rect 7849 5729 7883 5763
rect 9781 5729 9815 5763
rect 10333 5729 10367 5763
rect 10425 5729 10459 5763
rect 10977 5729 11011 5763
rect 14197 5729 14231 5763
rect 14564 5729 14598 5763
rect 14657 5729 14691 5763
rect 14749 5729 14783 5763
rect 14933 5729 14967 5763
rect 15025 5729 15059 5763
rect 15485 5729 15519 5763
rect 16957 5729 16991 5763
rect 17601 5729 17635 5763
rect 17785 5729 17819 5763
rect 17969 5729 18003 5763
rect 18429 5729 18463 5763
rect 19566 5729 19600 5763
rect 20085 5729 20119 5763
rect 20315 5729 20349 5763
rect 20728 5729 20762 5763
rect 20821 5729 20855 5763
rect 21373 5729 21407 5763
rect 21557 5729 21591 5763
rect 21649 5729 21683 5763
rect 22201 5729 22235 5763
rect 22385 5729 22419 5763
rect 23397 5729 23431 5763
rect 24041 5729 24075 5763
rect 24225 5729 24259 5763
rect 24409 5729 24443 5763
rect 24869 5729 24903 5763
rect 25053 5729 25087 5763
rect 25146 5729 25180 5763
rect 25421 5729 25455 5763
rect 25559 5729 25593 5763
rect 25789 5729 25823 5763
rect 26065 5729 26099 5763
rect 26617 5729 26651 5763
rect 26801 5729 26835 5763
rect 27169 5729 27203 5763
rect 27997 5729 28031 5763
rect 29469 5729 29503 5763
rect 29653 5729 29687 5763
rect 2605 5661 2639 5695
rect 5549 5661 5583 5695
rect 6377 5661 6411 5695
rect 7297 5661 7331 5695
rect 7573 5661 7607 5695
rect 9413 5661 9447 5695
rect 10149 5661 10183 5695
rect 13369 5661 13403 5695
rect 13829 5661 13863 5695
rect 16129 5661 16163 5695
rect 16681 5661 16715 5695
rect 23305 5661 23339 5695
rect 24317 5661 24351 5695
rect 24593 5661 24627 5695
rect 26893 5661 26927 5695
rect 27537 5661 27571 5695
rect 1593 5593 1627 5627
rect 5825 5593 5859 5627
rect 8401 5593 8435 5627
rect 9965 5593 9999 5627
rect 19993 5593 20027 5627
rect 21925 5593 21959 5627
rect 22569 5593 22603 5627
rect 25697 5593 25731 5627
rect 28181 5593 28215 5627
rect 28733 5593 28767 5627
rect 29377 5593 29411 5627
rect 4169 5525 4203 5559
rect 4905 5525 4939 5559
rect 8217 5525 8251 5559
rect 8861 5525 8895 5559
rect 10793 5525 10827 5559
rect 12725 5525 12759 5559
rect 13829 5525 13863 5559
rect 15669 5525 15703 5559
rect 19441 5525 19475 5559
rect 22201 5525 22235 5559
rect 22937 5525 22971 5559
rect 23121 5525 23155 5559
rect 23765 5525 23799 5559
rect 24501 5525 24535 5559
rect 24731 5525 24765 5559
rect 26249 5525 26283 5559
rect 26433 5525 26467 5559
rect 28549 5525 28583 5559
rect 28825 5525 28859 5559
rect 29009 5525 29043 5559
rect 29561 5525 29595 5559
rect 6193 5321 6227 5355
rect 10333 5321 10367 5355
rect 10701 5321 10735 5355
rect 11878 5321 11912 5355
rect 13967 5321 14001 5355
rect 16313 5321 16347 5355
rect 17693 5321 17727 5355
rect 19625 5321 19659 5355
rect 21005 5321 21039 5355
rect 22753 5321 22787 5355
rect 23581 5321 23615 5355
rect 25329 5321 25363 5355
rect 27261 5321 27295 5355
rect 6469 5253 6503 5287
rect 13369 5253 13403 5287
rect 14197 5253 14231 5287
rect 15853 5253 15887 5287
rect 19257 5253 19291 5287
rect 23857 5253 23891 5287
rect 24777 5253 24811 5287
rect 25513 5253 25547 5287
rect 857 5185 891 5219
rect 3893 5185 3927 5219
rect 4445 5185 4479 5219
rect 11437 5185 11471 5219
rect 11621 5185 11655 5219
rect 13645 5185 13679 5219
rect 14473 5185 14507 5219
rect 16957 5185 16991 5219
rect 17325 5185 17359 5219
rect 18061 5185 18095 5219
rect 18337 5185 18371 5219
rect 20821 5185 20855 5219
rect 21925 5185 21959 5219
rect 24869 5185 24903 5219
rect 25605 5185 25639 5219
rect 27997 5185 28031 5219
rect 3065 5117 3099 5151
rect 3709 5117 3743 5151
rect 8217 5117 8251 5151
rect 8585 5117 8619 5151
rect 10517 5117 10551 5151
rect 11161 5117 11195 5151
rect 13737 5117 13771 5151
rect 13829 5117 13863 5151
rect 14105 5117 14139 5151
rect 14289 5117 14323 5151
rect 14643 5117 14677 5151
rect 16037 5117 16071 5151
rect 16129 5117 16163 5151
rect 16865 5117 16899 5151
rect 17785 5117 17819 5151
rect 18153 5117 18187 5151
rect 18245 5117 18279 5151
rect 19533 5117 19567 5151
rect 19809 5117 19843 5151
rect 21097 5117 21131 5151
rect 21833 5117 21867 5151
rect 22201 5117 22235 5151
rect 22385 5117 22419 5151
rect 22661 5117 22695 5151
rect 23029 5117 23063 5151
rect 23121 5117 23155 5151
rect 24041 5117 24075 5151
rect 24133 5117 24167 5151
rect 25421 5117 25455 5151
rect 25697 5117 25731 5151
rect 26433 5117 26467 5151
rect 26617 5117 26651 5151
rect 26801 5117 26835 5151
rect 26893 5117 26927 5151
rect 27813 5117 27847 5151
rect 28273 5117 28307 5151
rect 28457 5117 28491 5151
rect 29469 5117 29503 5151
rect 1133 5049 1167 5083
rect 4721 5049 4755 5083
rect 7941 5049 7975 5083
rect 8861 5049 8895 5083
rect 15485 5049 15519 5083
rect 16313 5049 16347 5083
rect 21189 5049 21223 5083
rect 23305 5049 23339 5083
rect 23489 5049 23523 5083
rect 23857 5049 23891 5083
rect 24409 5049 24443 5083
rect 25881 5049 25915 5083
rect 25973 5049 26007 5083
rect 27261 5049 27295 5083
rect 27445 5049 27479 5083
rect 28089 5049 28123 5083
rect 29193 5049 29227 5083
rect 29377 5049 29411 5083
rect 2605 4981 2639 5015
rect 2881 4981 2915 5015
rect 3249 4981 3283 5015
rect 3617 4981 3651 5015
rect 10793 4981 10827 5015
rect 11253 4981 11287 5015
rect 14933 4981 14967 5015
rect 15945 4981 15979 5015
rect 17233 4981 17267 5015
rect 17877 4981 17911 5015
rect 20545 4981 20579 5015
rect 22477 4981 22511 5015
rect 24961 4981 24995 5015
rect 27077 4981 27111 5015
rect 27629 4981 27663 5015
rect 29009 4981 29043 5015
rect 29653 4981 29687 5015
rect 1133 4777 1167 4811
rect 2053 4777 2087 4811
rect 4261 4777 4295 4811
rect 4905 4777 4939 4811
rect 5273 4777 5307 4811
rect 8125 4777 8159 4811
rect 10701 4777 10735 4811
rect 14565 4777 14599 4811
rect 15025 4777 15059 4811
rect 15761 4777 15795 4811
rect 17601 4777 17635 4811
rect 18153 4777 18187 4811
rect 24225 4777 24259 4811
rect 2789 4709 2823 4743
rect 6193 4709 6227 4743
rect 13921 4709 13955 4743
rect 17049 4709 17083 4743
rect 18245 4709 18279 4743
rect 20637 4709 20671 4743
rect 21741 4709 21775 4743
rect 26433 4709 26467 4743
rect 26649 4709 26683 4743
rect 27721 4709 27755 4743
rect 27905 4709 27939 4743
rect 949 4641 983 4675
rect 1409 4641 1443 4675
rect 2513 4641 2547 4675
rect 4629 4641 4663 4675
rect 5365 4641 5399 4675
rect 10149 4641 10183 4675
rect 10425 4641 10459 4675
rect 10517 4641 10551 4675
rect 10977 4641 11011 4675
rect 11253 4641 11287 4675
rect 13277 4641 13311 4675
rect 14473 4641 14507 4675
rect 14657 4641 14691 4675
rect 14749 4641 14783 4675
rect 14933 4641 14967 4675
rect 15209 4641 15243 4675
rect 15393 4641 15427 4675
rect 15485 4641 15519 4675
rect 15577 4641 15611 4675
rect 16129 4641 16163 4675
rect 16313 4641 16347 4675
rect 16865 4641 16899 4675
rect 17141 4641 17175 4675
rect 17785 4641 17819 4675
rect 18521 4641 18555 4675
rect 19257 4641 19291 4675
rect 19441 4641 19475 4675
rect 19533 4641 19567 4675
rect 19901 4641 19935 4675
rect 20448 4641 20482 4675
rect 20545 4641 20579 4675
rect 20820 4641 20854 4675
rect 20913 4641 20947 4675
rect 21649 4641 21683 4675
rect 22109 4641 22143 4675
rect 22477 4641 22511 4675
rect 22661 4641 22695 4675
rect 22937 4641 22971 4675
rect 23121 4641 23155 4675
rect 23213 4641 23247 4675
rect 23305 4641 23339 4675
rect 23673 4641 23707 4675
rect 23949 4641 23983 4675
rect 24041 4641 24075 4675
rect 24961 4641 24995 4675
rect 25605 4641 25639 4675
rect 25697 4641 25731 4675
rect 25881 4641 25915 4675
rect 25973 4641 26007 4675
rect 27077 4641 27111 4675
rect 27537 4641 27571 4675
rect 2145 4573 2179 4607
rect 2329 4573 2363 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 9873 4573 9907 4607
rect 11529 4573 11563 4607
rect 13921 4573 13955 4607
rect 14013 4573 14047 4607
rect 14841 4573 14875 4607
rect 16221 4573 16255 4607
rect 17877 4573 17911 4607
rect 18245 4573 18279 4607
rect 19625 4573 19659 4607
rect 19993 4573 20027 4607
rect 22017 4573 22051 4607
rect 23581 4573 23615 4607
rect 25053 4573 25087 4607
rect 27169 4573 27203 4607
rect 1685 4505 1719 4539
rect 10241 4505 10275 4539
rect 11161 4505 11195 4539
rect 13001 4505 13035 4539
rect 13093 4505 13127 4539
rect 13461 4505 13495 4539
rect 20269 4505 20303 4539
rect 26801 4505 26835 4539
rect 27445 4505 27479 4539
rect 1225 4437 1259 4471
rect 4813 4437 4847 4471
rect 6101 4437 6135 4471
rect 8401 4437 8435 4471
rect 16681 4437 16715 4471
rect 17233 4437 17267 4471
rect 17785 4437 17819 4471
rect 18429 4437 18463 4471
rect 19349 4437 19383 4471
rect 20177 4437 20211 4471
rect 23765 4437 23799 4471
rect 24685 4437 24719 4471
rect 25421 4437 25455 4471
rect 26617 4437 26651 4471
rect 1041 4233 1075 4267
rect 4794 4233 4828 4267
rect 6285 4233 6319 4267
rect 8217 4233 8251 4267
rect 9781 4233 9815 4267
rect 10885 4233 10919 4267
rect 14749 4233 14783 4267
rect 15117 4233 15151 4267
rect 15669 4233 15703 4267
rect 18981 4233 19015 4267
rect 24133 4233 24167 4267
rect 25881 4233 25915 4267
rect 26249 4233 26283 4267
rect 9413 4165 9447 4199
rect 15485 4165 15519 4199
rect 17785 4165 17819 4199
rect 17877 4165 17911 4199
rect 23489 4165 23523 4199
rect 26341 4165 26375 4199
rect 27629 4165 27663 4199
rect 27997 4165 28031 4199
rect 1133 4097 1167 4131
rect 2881 4097 2915 4131
rect 3801 4097 3835 4131
rect 7665 4097 7699 4131
rect 8769 4097 8803 4131
rect 8953 4097 8987 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 11529 4097 11563 4131
rect 13645 4097 13679 4131
rect 16221 4097 16255 4131
rect 16497 4097 16531 4131
rect 21925 4097 21959 4131
rect 22017 4097 22051 4131
rect 22385 4097 22419 4131
rect 22753 4097 22787 4131
rect 24133 4097 24167 4131
rect 24961 4097 24995 4131
rect 28089 4097 28123 4131
rect 857 4029 891 4063
rect 4445 4029 4479 4063
rect 4537 4029 4571 4063
rect 6469 4029 6503 4063
rect 7481 4029 7515 4063
rect 8033 4029 8067 4063
rect 8401 4029 8435 4063
rect 11253 4029 11287 4063
rect 11345 4029 11379 4063
rect 14105 4029 14139 4063
rect 14289 4029 14323 4063
rect 14381 4029 14415 4063
rect 15025 4029 15059 4063
rect 15117 4029 15151 4063
rect 15393 4029 15427 4063
rect 15577 4029 15611 4063
rect 16405 4029 16439 4063
rect 16957 4029 16991 4063
rect 17141 4029 17175 4063
rect 17785 4029 17819 4063
rect 19165 4029 19199 4063
rect 19257 4029 19291 4063
rect 19441 4029 19475 4063
rect 19533 4029 19567 4063
rect 20085 4029 20119 4063
rect 20177 4029 20211 4063
rect 20361 4029 20395 4063
rect 20453 4029 20487 4063
rect 20821 4029 20855 4063
rect 20914 4029 20948 4063
rect 21189 4029 21223 4063
rect 21286 4029 21320 4063
rect 21741 4029 21775 4063
rect 22569 4029 22603 4063
rect 23029 4029 23063 4063
rect 23213 4029 23247 4063
rect 23489 4029 23523 4063
rect 23673 4029 23707 4063
rect 24409 4029 24443 4063
rect 25053 4029 25087 4063
rect 25513 4029 25547 4063
rect 25697 4029 25731 4063
rect 25789 4029 25823 4063
rect 26065 4029 26099 4063
rect 26520 4029 26554 4063
rect 26617 4029 26651 4063
rect 26892 4029 26926 4063
rect 26985 4029 27019 4063
rect 27077 4029 27111 4063
rect 27169 4029 27203 4063
rect 27353 4029 27387 4063
rect 27445 4029 27479 4063
rect 27905 4029 27939 4063
rect 1409 3961 1443 3995
rect 7021 3961 7055 3995
rect 7573 3961 7607 3995
rect 9045 3961 9079 3995
rect 9781 3961 9815 3995
rect 9965 3961 9999 3995
rect 15209 3961 15243 3995
rect 16865 3961 16899 3995
rect 18061 3961 18095 3995
rect 21097 3961 21131 3995
rect 25605 3961 25639 3995
rect 26709 3961 26743 3995
rect 27721 3961 27755 3995
rect 28181 3961 28215 3995
rect 3249 3893 3283 3927
rect 3617 3893 3651 3927
rect 3709 3893 3743 3927
rect 4261 3893 4295 3927
rect 7113 3893 7147 3927
rect 8585 3893 8619 3927
rect 9597 3893 9631 3927
rect 10057 3893 10091 3927
rect 10425 3893 10459 3927
rect 17049 3893 17083 3927
rect 19901 3893 19935 3927
rect 21465 3893 21499 3927
rect 21557 3893 21591 3927
rect 23857 3893 23891 3927
rect 24777 3893 24811 3927
rect 25421 3893 25455 3927
rect 9965 3689 9999 3723
rect 11253 3689 11287 3723
rect 13093 3689 13127 3723
rect 14933 3689 14967 3723
rect 16221 3689 16255 3723
rect 17969 3689 18003 3723
rect 18153 3689 18187 3723
rect 20913 3689 20947 3723
rect 24041 3689 24075 3723
rect 26249 3689 26283 3723
rect 4169 3621 4203 3655
rect 6561 3621 6595 3655
rect 8401 3621 8435 3655
rect 11621 3621 11655 3655
rect 13829 3621 13863 3655
rect 21649 3621 21683 3655
rect 24409 3621 24443 3655
rect 1685 3553 1719 3587
rect 2053 3553 2087 3587
rect 3893 3553 3927 3587
rect 6009 3553 6043 3587
rect 10517 3553 10551 3587
rect 11069 3553 11103 3587
rect 11345 3553 11379 3587
rect 14289 3553 14323 3587
rect 14473 3553 14507 3587
rect 15301 3553 15335 3587
rect 16589 3553 16623 3587
rect 17325 3553 17359 3587
rect 17509 3553 17543 3587
rect 17601 3553 17635 3587
rect 17785 3553 17819 3587
rect 18061 3553 18095 3587
rect 18245 3553 18279 3587
rect 18521 3553 18555 3587
rect 18705 3553 18739 3587
rect 19073 3553 19107 3587
rect 19809 3553 19843 3587
rect 20821 3553 20855 3587
rect 21005 3553 21039 3587
rect 21281 3553 21315 3587
rect 21429 3553 21463 3587
rect 21557 3553 21591 3587
rect 21746 3553 21780 3587
rect 22201 3553 22235 3587
rect 22293 3553 22327 3587
rect 23489 3553 23523 3587
rect 23949 3553 23983 3587
rect 24225 3553 24259 3587
rect 24685 3553 24719 3587
rect 24777 3553 24811 3587
rect 26065 3553 26099 3587
rect 26249 3553 26283 3587
rect 27445 3553 27479 3587
rect 27813 3553 27847 3587
rect 2329 3485 2363 3519
rect 3801 3485 3835 3519
rect 5641 3485 5675 3519
rect 6285 3485 6319 3519
rect 8125 3485 8159 3519
rect 9873 3485 9907 3519
rect 14565 3485 14599 3519
rect 15209 3485 15243 3519
rect 16681 3485 16715 3519
rect 17141 3485 17175 3519
rect 20729 3485 20763 3519
rect 23305 3485 23339 3519
rect 23397 3485 23431 3519
rect 23581 3485 23615 3519
rect 24317 3485 24351 3519
rect 26709 3485 26743 3519
rect 27537 3485 27571 3519
rect 27905 3485 27939 3519
rect 1501 3417 1535 3451
rect 18337 3417 18371 3451
rect 21925 3417 21959 3451
rect 22017 3417 22051 3451
rect 6193 3349 6227 3383
rect 8033 3349 8067 3383
rect 23121 3349 23155 3383
rect 24225 3349 24259 3383
rect 24961 3349 24995 3383
rect 1869 3145 1903 3179
rect 2789 3145 2823 3179
rect 3801 3145 3835 3179
rect 5825 3145 5859 3179
rect 6745 3145 6779 3179
rect 8033 3145 8067 3179
rect 8493 3145 8527 3179
rect 11713 3145 11747 3179
rect 14933 3145 14967 3179
rect 15301 3145 15335 3179
rect 15485 3145 15519 3179
rect 16681 3145 16715 3179
rect 17509 3145 17543 3179
rect 18889 3145 18923 3179
rect 19809 3145 19843 3179
rect 20453 3145 20487 3179
rect 23305 3145 23339 3179
rect 24041 3145 24075 3179
rect 25697 3145 25731 3179
rect 26801 3145 26835 3179
rect 27169 3145 27203 3179
rect 8769 3077 8803 3111
rect 19993 3077 20027 3111
rect 25053 3077 25087 3111
rect 2513 3009 2547 3043
rect 4353 3009 4387 3043
rect 6469 3009 6503 3043
rect 7665 3009 7699 3043
rect 9321 3009 9355 3043
rect 9873 3009 9907 3043
rect 10149 3009 10183 3043
rect 12265 3009 12299 3043
rect 13553 3009 13587 3043
rect 14289 3009 14323 3043
rect 15945 3009 15979 3043
rect 19901 3009 19935 3043
rect 21005 3009 21039 3043
rect 23121 3009 23155 3043
rect 27077 3009 27111 3043
rect 2329 2941 2363 2975
rect 2973 2941 3007 2975
rect 6929 2941 6963 2975
rect 7389 2941 7423 2975
rect 8217 2941 8251 2975
rect 8677 2941 8711 2975
rect 9137 2941 9171 2975
rect 12173 2941 12207 2975
rect 14013 2941 14047 2975
rect 14197 2941 14231 2975
rect 15393 2941 15427 2975
rect 15669 2941 15703 2975
rect 15853 2941 15887 2975
rect 16865 2941 16899 2975
rect 17141 2941 17175 2975
rect 17233 2941 17267 2975
rect 17785 2941 17819 2975
rect 17969 2941 18003 2975
rect 18153 2941 18187 2975
rect 19438 2941 19472 2975
rect 19993 2941 20027 2975
rect 20177 2941 20211 2975
rect 20913 2941 20947 2975
rect 21649 2941 21683 2975
rect 21833 2941 21867 2975
rect 22661 2941 22695 2975
rect 22845 2941 22879 2975
rect 22937 2941 22971 2975
rect 23213 2941 23247 2975
rect 23489 2941 23523 2975
rect 23857 2941 23891 2975
rect 24041 2941 24075 2975
rect 24133 2941 24167 2975
rect 24317 2941 24351 2975
rect 24409 2941 24443 2975
rect 24557 2941 24591 2975
rect 24777 2941 24811 2975
rect 24915 2941 24949 2975
rect 25145 2941 25179 2975
rect 25237 2941 25271 2975
rect 25421 2941 25455 2975
rect 25513 2941 25547 2975
rect 26617 2941 26651 2975
rect 26893 2941 26927 2975
rect 26985 2941 27019 2975
rect 2237 2873 2271 2907
rect 12081 2873 12115 2907
rect 18705 2873 18739 2907
rect 20821 2873 20855 2907
rect 22201 2873 22235 2907
rect 22385 2873 22419 2907
rect 23673 2873 23707 2907
rect 24685 2873 24719 2907
rect 7021 2805 7055 2839
rect 7481 2805 7515 2839
rect 9229 2805 9263 2839
rect 11621 2805 11655 2839
rect 17049 2805 17083 2839
rect 17693 2805 17727 2839
rect 18905 2805 18939 2839
rect 19073 2805 19107 2839
rect 19257 2805 19291 2839
rect 19441 2805 19475 2839
rect 21465 2805 21499 2839
rect 22017 2805 22051 2839
rect 24133 2805 24167 2839
rect 26433 2805 26467 2839
rect 27353 2805 27387 2839
rect 7757 2601 7791 2635
rect 9597 2601 9631 2635
rect 15577 2601 15611 2635
rect 17325 2601 17359 2635
rect 18245 2601 18279 2635
rect 18521 2601 18555 2635
rect 21373 2601 21407 2635
rect 22661 2601 22695 2635
rect 23305 2601 23339 2635
rect 26157 2601 26191 2635
rect 27077 2601 27111 2635
rect 13553 2533 13587 2567
rect 15761 2533 15795 2567
rect 18797 2533 18831 2567
rect 21557 2533 21591 2567
rect 23489 2533 23523 2567
rect 25605 2533 25639 2567
rect 27537 2533 27571 2567
rect 8401 2465 8435 2499
rect 10149 2465 10183 2499
rect 14013 2465 14047 2499
rect 14197 2465 14231 2499
rect 14289 2465 14323 2499
rect 15209 2465 15243 2499
rect 15393 2465 15427 2499
rect 15669 2465 15703 2499
rect 15853 2455 15887 2489
rect 16681 2465 16715 2499
rect 16957 2465 16991 2499
rect 17601 2465 17635 2499
rect 18429 2465 18463 2499
rect 18613 2465 18647 2499
rect 19073 2465 19107 2499
rect 19165 2465 19199 2499
rect 19349 2465 19383 2499
rect 19441 2465 19475 2499
rect 19809 2465 19843 2499
rect 20821 2465 20855 2499
rect 21005 2465 21039 2499
rect 21097 2465 21131 2499
rect 21281 2465 21315 2499
rect 21741 2465 21775 2499
rect 22017 2465 22051 2499
rect 22201 2465 22235 2499
rect 22385 2465 22419 2499
rect 23397 2465 23431 2499
rect 23581 2465 23615 2499
rect 23949 2465 23983 2499
rect 24133 2465 24167 2499
rect 24225 2465 24259 2499
rect 24409 2465 24443 2499
rect 24593 2465 24627 2499
rect 25513 2465 25547 2499
rect 25697 2465 25731 2499
rect 25973 2465 26007 2499
rect 26249 2465 26283 2499
rect 26433 2465 26467 2499
rect 26801 2465 26835 2499
rect 15117 2397 15151 2431
rect 15301 2397 15335 2431
rect 16221 2397 16255 2431
rect 17325 2397 17359 2431
rect 17877 2397 17911 2431
rect 18061 2397 18095 2431
rect 19717 2397 19751 2431
rect 22845 2397 22879 2431
rect 22937 2397 22971 2431
rect 25329 2397 25363 2431
rect 26985 2397 27019 2431
rect 20637 2329 20671 2363
rect 21557 2329 21591 2363
rect 25973 2329 26007 2363
rect 26525 2329 26559 2363
rect 27261 2329 27295 2363
rect 18889 2261 18923 2295
rect 21741 2261 21775 2295
rect 23765 2261 23799 2295
rect 14565 2057 14599 2091
rect 18153 2057 18187 2091
rect 18889 2057 18923 2091
rect 19349 2057 19383 2091
rect 21097 2057 21131 2091
rect 22293 2057 22327 2091
rect 24409 2057 24443 2091
rect 25145 2057 25179 2091
rect 25421 2057 25455 2091
rect 26525 2057 26559 2091
rect 26617 2057 26651 2091
rect 15117 1989 15151 2023
rect 19993 1989 20027 2023
rect 15577 1921 15611 1955
rect 17141 1921 17175 1955
rect 17417 1921 17451 1955
rect 19165 1921 19199 1955
rect 20453 1921 20487 1955
rect 20729 1921 20763 1955
rect 21925 1921 21959 1955
rect 24869 1921 24903 1955
rect 26433 1921 26467 1955
rect 14933 1853 14967 1887
rect 15485 1853 15519 1887
rect 17049 1853 17083 1887
rect 18337 1853 18371 1887
rect 19441 1853 19475 1887
rect 19539 1853 19573 1887
rect 19717 1853 19751 1887
rect 20361 1853 20395 1887
rect 20821 1853 20855 1887
rect 21281 1853 21315 1887
rect 21465 1853 21499 1887
rect 22017 1853 22051 1887
rect 24777 1853 24811 1887
rect 25053 1853 25087 1887
rect 25237 1853 25271 1887
rect 25329 1853 25363 1887
rect 26709 1853 26743 1887
rect 14749 1785 14783 1819
rect 18521 1785 18555 1819
rect 21373 1785 21407 1819
rect 19625 1717 19659 1751
rect 18981 1513 19015 1547
rect 18981 1377 19015 1411
rect 19349 1377 19383 1411
rect 19533 1377 19567 1411
rect 19717 1377 19751 1411
rect 19073 1309 19107 1343
rect 19257 1173 19291 1207
rect 19533 1173 19567 1207
<< metal1 >>
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5132 21984 10364 22012
rect 5132 21972 5138 21984
rect 10336 21956 10364 21984
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 24578 22012 24584 22024
rect 15252 21984 24584 22012
rect 15252 21972 15258 21984
rect 24578 21972 24584 21984
rect 24636 22012 24642 22024
rect 26878 22012 26884 22024
rect 24636 21984 26884 22012
rect 24636 21972 24642 21984
rect 26878 21972 26884 21984
rect 26936 22012 26942 22024
rect 30374 22012 30380 22024
rect 26936 21984 30380 22012
rect 26936 21972 26942 21984
rect 30374 21972 30380 21984
rect 30432 21972 30438 22024
rect 4062 21904 4068 21956
rect 4120 21944 4126 21956
rect 10134 21944 10140 21956
rect 4120 21916 10140 21944
rect 4120 21904 4126 21916
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 10318 21904 10324 21956
rect 10376 21904 10382 21956
rect 3510 21836 3516 21888
rect 3568 21876 3574 21888
rect 15838 21876 15844 21888
rect 3568 21848 15844 21876
rect 3568 21836 3574 21848
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 25314 21836 25320 21888
rect 25372 21876 25378 21888
rect 30834 21876 30840 21888
rect 25372 21848 30840 21876
rect 25372 21836 25378 21848
rect 30834 21836 30840 21848
rect 30892 21836 30898 21888
rect 552 21786 31648 21808
rect 552 21734 4285 21786
rect 4337 21734 4349 21786
rect 4401 21734 4413 21786
rect 4465 21734 4477 21786
rect 4529 21734 4541 21786
rect 4593 21734 12059 21786
rect 12111 21734 12123 21786
rect 12175 21734 12187 21786
rect 12239 21734 12251 21786
rect 12303 21734 12315 21786
rect 12367 21734 19833 21786
rect 19885 21734 19897 21786
rect 19949 21734 19961 21786
rect 20013 21734 20025 21786
rect 20077 21734 20089 21786
rect 20141 21734 27607 21786
rect 27659 21734 27671 21786
rect 27723 21734 27735 21786
rect 27787 21734 27799 21786
rect 27851 21734 27863 21786
rect 27915 21734 31648 21786
rect 552 21712 31648 21734
rect 6362 21632 6368 21684
rect 6420 21632 6426 21684
rect 7006 21632 7012 21684
rect 7064 21632 7070 21684
rect 8128 21644 8708 21672
rect 4982 21564 4988 21616
rect 5040 21604 5046 21616
rect 6380 21604 6408 21632
rect 8128 21604 8156 21644
rect 5040 21576 5672 21604
rect 6380 21576 8156 21604
rect 8205 21607 8263 21613
rect 5040 21564 5046 21576
rect 1302 21496 1308 21548
rect 1360 21496 1366 21548
rect 3605 21539 3663 21545
rect 3605 21505 3617 21539
rect 3651 21536 3663 21539
rect 5534 21536 5540 21548
rect 3651 21508 5540 21536
rect 3651 21505 3663 21508
rect 3605 21499 3663 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5644 21545 5672 21576
rect 8205 21573 8217 21607
rect 8251 21573 8263 21607
rect 8205 21567 8263 21573
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 6270 21496 6276 21548
rect 6328 21536 6334 21548
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 6328 21508 6377 21536
rect 6328 21496 6334 21508
rect 6365 21505 6377 21508
rect 6411 21536 6423 21539
rect 7561 21539 7619 21545
rect 7561 21536 7573 21539
rect 6411 21508 7573 21536
rect 6411 21505 6423 21508
rect 6365 21499 6423 21505
rect 7561 21505 7573 21508
rect 7607 21505 7619 21539
rect 7561 21499 7619 21505
rect 2682 21428 2688 21480
rect 2740 21428 2746 21480
rect 3053 21471 3111 21477
rect 3053 21437 3065 21471
rect 3099 21437 3111 21471
rect 3053 21431 3111 21437
rect 2222 21360 2228 21412
rect 2280 21360 2286 21412
rect 3068 21400 3096 21431
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7024 21440 7849 21468
rect 7024 21412 7052 21440
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 8220 21468 8248 21567
rect 8680 21536 8708 21644
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 8904 21644 10241 21672
rect 8904 21632 8910 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 12526 21632 12532 21684
rect 12584 21632 12590 21684
rect 13814 21632 13820 21684
rect 13872 21632 13878 21684
rect 14093 21675 14151 21681
rect 14093 21641 14105 21675
rect 14139 21672 14151 21675
rect 14369 21675 14427 21681
rect 14369 21672 14381 21675
rect 14139 21644 14381 21672
rect 14139 21641 14151 21644
rect 14093 21635 14151 21641
rect 14369 21641 14381 21644
rect 14415 21641 14427 21675
rect 14369 21635 14427 21641
rect 16574 21632 16580 21684
rect 16632 21632 16638 21684
rect 20438 21672 20444 21684
rect 16960 21644 20444 21672
rect 8757 21607 8815 21613
rect 8757 21573 8769 21607
rect 8803 21604 8815 21607
rect 12342 21604 12348 21616
rect 8803 21576 9904 21604
rect 8803 21573 8815 21576
rect 8757 21567 8815 21573
rect 9030 21536 9036 21548
rect 8680 21508 9036 21536
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 9766 21536 9772 21548
rect 9539 21508 9772 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8220 21440 9137 21468
rect 7837 21431 7895 21437
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9416 21468 9444 21499
rect 9766 21496 9772 21508
rect 9824 21496 9830 21548
rect 9876 21536 9904 21576
rect 11072 21576 12348 21604
rect 11072 21536 11100 21576
rect 12342 21564 12348 21576
rect 12400 21564 12406 21616
rect 13541 21607 13599 21613
rect 13541 21573 13553 21607
rect 13587 21604 13599 21607
rect 13630 21604 13636 21616
rect 13587 21576 13636 21604
rect 13587 21573 13599 21576
rect 13541 21567 13599 21573
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 13832 21604 13860 21632
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 13832 21576 14841 21604
rect 14829 21573 14841 21576
rect 14875 21573 14887 21607
rect 16960 21604 16988 21644
rect 20438 21632 20444 21644
rect 20496 21672 20502 21684
rect 20625 21675 20683 21681
rect 20496 21644 20576 21672
rect 20496 21632 20502 21644
rect 14829 21567 14887 21573
rect 16546 21576 16988 21604
rect 17037 21607 17095 21613
rect 9876 21508 11100 21536
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 13170 21536 13176 21548
rect 11195 21508 13176 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 13280 21508 13860 21536
rect 9674 21468 9680 21480
rect 9416 21440 9680 21468
rect 9125 21431 9183 21437
rect 9674 21428 9680 21440
rect 9732 21428 9738 21480
rect 9876 21440 10272 21468
rect 3602 21400 3608 21412
rect 3068 21372 3608 21400
rect 3602 21360 3608 21372
rect 3660 21360 3666 21412
rect 3878 21360 3884 21412
rect 3936 21360 3942 21412
rect 6914 21400 6920 21412
rect 5106 21372 6920 21400
rect 6914 21360 6920 21372
rect 6972 21360 6978 21412
rect 7006 21360 7012 21412
rect 7064 21360 7070 21412
rect 7282 21360 7288 21412
rect 7340 21360 7346 21412
rect 7374 21360 7380 21412
rect 7432 21400 7438 21412
rect 8481 21403 8539 21409
rect 8481 21400 8493 21403
rect 7432 21372 8493 21400
rect 7432 21360 7438 21372
rect 8481 21369 8493 21372
rect 8527 21369 8539 21403
rect 9876 21400 9904 21440
rect 8481 21363 8539 21369
rect 8864 21372 9904 21400
rect 10137 21403 10195 21409
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 3329 21335 3387 21341
rect 3329 21332 3341 21335
rect 3016 21304 3341 21332
rect 3016 21292 3022 21304
rect 3329 21301 3341 21304
rect 3375 21332 3387 21335
rect 3786 21332 3792 21344
rect 3375 21304 3792 21332
rect 3375 21301 3387 21304
rect 3329 21295 3387 21301
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 4672 21304 5825 21332
rect 4672 21292 4678 21304
rect 5813 21301 5825 21304
rect 5859 21301 5871 21335
rect 5813 21295 5871 21301
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 6273 21335 6331 21341
rect 6273 21301 6285 21335
rect 6319 21332 6331 21335
rect 6362 21332 6368 21344
rect 6319 21304 6368 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6825 21335 6883 21341
rect 6825 21301 6837 21335
rect 6871 21332 6883 21335
rect 7190 21332 7196 21344
rect 6871 21304 7196 21332
rect 6871 21301 6883 21304
rect 6825 21295 6883 21301
rect 7190 21292 7196 21304
rect 7248 21292 7254 21344
rect 7745 21335 7803 21341
rect 7745 21301 7757 21335
rect 7791 21332 7803 21335
rect 8864 21332 8892 21372
rect 10137 21369 10149 21403
rect 10183 21369 10195 21403
rect 10244 21400 10272 21440
rect 10502 21428 10508 21480
rect 10560 21468 10566 21480
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 10560 21440 12449 21468
rect 10560 21428 10566 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 12897 21471 12955 21477
rect 12897 21437 12909 21471
rect 12943 21468 12955 21471
rect 13280 21468 13308 21508
rect 12943 21440 13308 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 13725 21471 13783 21477
rect 13725 21470 13737 21471
rect 13648 21468 13737 21470
rect 13596 21442 13737 21468
rect 13596 21440 13676 21442
rect 13596 21428 13602 21440
rect 13725 21437 13737 21442
rect 13771 21437 13783 21471
rect 13832 21468 13860 21508
rect 13906 21496 13912 21548
rect 13964 21536 13970 21548
rect 16546 21536 16574 21576
rect 17037 21573 17049 21607
rect 17083 21573 17095 21607
rect 17037 21567 17095 21573
rect 18969 21607 19027 21613
rect 18969 21573 18981 21607
rect 19015 21604 19027 21607
rect 20254 21604 20260 21616
rect 19015 21576 20260 21604
rect 19015 21573 19027 21576
rect 18969 21567 19027 21573
rect 13964 21508 16574 21536
rect 17052 21536 17080 21567
rect 20254 21564 20260 21576
rect 20312 21564 20318 21616
rect 20548 21604 20576 21644
rect 20625 21641 20637 21675
rect 20671 21672 20683 21675
rect 20714 21672 20720 21684
rect 20671 21644 20720 21672
rect 20671 21641 20683 21644
rect 20625 21635 20683 21641
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 26697 21675 26755 21681
rect 26697 21672 26709 21675
rect 22060 21644 26709 21672
rect 22060 21632 22066 21644
rect 26697 21641 26709 21644
rect 26743 21641 26755 21675
rect 26697 21635 26755 21641
rect 28442 21632 28448 21684
rect 28500 21672 28506 21684
rect 29825 21675 29883 21681
rect 29825 21672 29837 21675
rect 28500 21644 29837 21672
rect 28500 21632 28506 21644
rect 29825 21641 29837 21644
rect 29871 21641 29883 21675
rect 29825 21635 29883 21641
rect 21450 21604 21456 21616
rect 20548 21576 21456 21604
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 21545 21607 21603 21613
rect 21545 21573 21557 21607
rect 21591 21604 21603 21607
rect 24489 21607 24547 21613
rect 24489 21604 24501 21607
rect 21591 21576 24501 21604
rect 21591 21573 21603 21576
rect 21545 21567 21603 21573
rect 24489 21573 24501 21576
rect 24535 21573 24547 21607
rect 24489 21567 24547 21573
rect 25501 21607 25559 21613
rect 25501 21573 25513 21607
rect 25547 21604 25559 21607
rect 26421 21607 26479 21613
rect 26421 21604 26433 21607
rect 25547 21576 26433 21604
rect 25547 21573 25559 21576
rect 25501 21567 25559 21573
rect 26421 21573 26433 21576
rect 26467 21573 26479 21607
rect 26421 21567 26479 21573
rect 26881 21607 26939 21613
rect 26881 21573 26893 21607
rect 26927 21604 26939 21607
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 26927 21576 27537 21604
rect 26927 21573 26939 21576
rect 26881 21567 26939 21573
rect 27525 21573 27537 21576
rect 27571 21573 27583 21607
rect 29549 21607 29607 21613
rect 29549 21604 29561 21607
rect 27525 21567 27583 21573
rect 27632 21576 29561 21604
rect 25866 21536 25872 21548
rect 17052 21508 24072 21536
rect 13964 21496 13970 21508
rect 14645 21471 14703 21477
rect 14645 21468 14657 21471
rect 13832 21440 14657 21468
rect 13725 21431 13783 21437
rect 14645 21437 14657 21440
rect 14691 21437 14703 21471
rect 14645 21431 14703 21437
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 16485 21471 16543 21477
rect 16485 21468 16497 21471
rect 15344 21440 16497 21468
rect 15344 21428 15350 21440
rect 16485 21437 16497 21440
rect 16531 21437 16543 21471
rect 16485 21431 16543 21437
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21468 16911 21471
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 16899 21440 18705 21468
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21437 18935 21471
rect 18877 21431 18935 21437
rect 11238 21400 11244 21412
rect 10244 21372 11244 21400
rect 10137 21363 10195 21369
rect 7791 21304 8892 21332
rect 7791 21301 7803 21304
rect 7745 21295 7803 21301
rect 8938 21292 8944 21344
rect 8996 21292 9002 21344
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 9585 21335 9643 21341
rect 9585 21332 9597 21335
rect 9180 21304 9597 21332
rect 9180 21292 9186 21304
rect 9585 21301 9597 21304
rect 9631 21301 9643 21335
rect 9585 21295 9643 21301
rect 9953 21335 10011 21341
rect 9953 21301 9965 21335
rect 9999 21332 10011 21335
rect 10152 21332 10180 21363
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 11330 21360 11336 21412
rect 11388 21400 11394 21412
rect 11425 21403 11483 21409
rect 11425 21400 11437 21403
rect 11388 21372 11437 21400
rect 11388 21360 11394 21372
rect 11425 21369 11437 21372
rect 11471 21369 11483 21403
rect 11425 21363 11483 21369
rect 11698 21360 11704 21412
rect 11756 21400 11762 21412
rect 11885 21403 11943 21409
rect 11885 21400 11897 21403
rect 11756 21372 11897 21400
rect 11756 21360 11762 21372
rect 11885 21369 11897 21372
rect 11931 21369 11943 21403
rect 11885 21363 11943 21369
rect 12342 21360 12348 21412
rect 12400 21360 12406 21412
rect 12986 21360 12992 21412
rect 13044 21400 13050 21412
rect 13081 21403 13139 21409
rect 13081 21400 13093 21403
rect 13044 21372 13093 21400
rect 13044 21360 13050 21372
rect 13081 21369 13093 21372
rect 13127 21369 13139 21403
rect 13081 21363 13139 21369
rect 13262 21360 13268 21412
rect 13320 21360 13326 21412
rect 14200 21372 14504 21400
rect 9999 21304 10180 21332
rect 12161 21335 12219 21341
rect 9999 21301 10011 21304
rect 9953 21295 10011 21301
rect 12161 21301 12173 21335
rect 12207 21332 12219 21335
rect 12250 21332 12256 21344
rect 12207 21304 12256 21332
rect 12207 21301 12219 21304
rect 12161 21295 12219 21301
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12360 21332 12388 21360
rect 14200 21344 14228 21372
rect 13354 21332 13360 21344
rect 12360 21304 13360 21332
rect 13354 21292 13360 21304
rect 13412 21332 13418 21344
rect 13817 21335 13875 21341
rect 13817 21332 13829 21335
rect 13412 21304 13829 21332
rect 13412 21292 13418 21304
rect 13817 21301 13829 21304
rect 13863 21301 13875 21335
rect 13817 21295 13875 21301
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 14182 21292 14188 21344
rect 14240 21292 14246 21344
rect 14366 21341 14372 21344
rect 14353 21335 14372 21341
rect 14353 21301 14365 21335
rect 14353 21295 14372 21301
rect 14366 21292 14372 21295
rect 14424 21292 14430 21344
rect 14476 21332 14504 21372
rect 14550 21360 14556 21412
rect 14608 21400 14614 21412
rect 15102 21400 15108 21412
rect 14608 21372 15108 21400
rect 14608 21360 14614 21372
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 16666 21332 16672 21344
rect 14476 21304 16672 21332
rect 16666 21292 16672 21304
rect 16724 21292 16730 21344
rect 18892 21332 18920 21431
rect 19058 21428 19064 21480
rect 19116 21428 19122 21480
rect 19150 21428 19156 21480
rect 19208 21428 19214 21480
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21437 19395 21471
rect 19337 21431 19395 21437
rect 19352 21400 19380 21431
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 20441 21471 20499 21477
rect 20441 21468 20453 21471
rect 19576 21440 20453 21468
rect 19576 21428 19582 21440
rect 20441 21437 20453 21440
rect 20487 21437 20499 21471
rect 20441 21431 20499 21437
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 20625 21471 20683 21477
rect 20625 21468 20637 21471
rect 20588 21440 20637 21468
rect 20588 21428 20594 21440
rect 20625 21437 20637 21440
rect 20671 21437 20683 21471
rect 20625 21431 20683 21437
rect 21450 21428 21456 21480
rect 21508 21468 21514 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 21508 21440 21833 21468
rect 21508 21428 21514 21440
rect 21821 21437 21833 21440
rect 21867 21468 21879 21471
rect 23934 21468 23940 21480
rect 21867 21440 23940 21468
rect 21867 21437 21879 21440
rect 21821 21431 21879 21437
rect 23934 21428 23940 21440
rect 23992 21428 23998 21480
rect 24044 21477 24072 21508
rect 24228 21508 25872 21536
rect 24029 21471 24087 21477
rect 24029 21437 24041 21471
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 20990 21400 20996 21412
rect 19352 21372 20996 21400
rect 20990 21360 20996 21372
rect 21048 21360 21054 21412
rect 24228 21400 24256 21508
rect 25866 21496 25872 21508
rect 25924 21496 25930 21548
rect 24670 21428 24676 21480
rect 24728 21428 24734 21480
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 24912 21440 25789 21468
rect 24912 21428 24918 21440
rect 25777 21437 25789 21440
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 26602 21428 26608 21480
rect 26660 21428 26666 21480
rect 27430 21428 27436 21480
rect 27488 21428 27494 21480
rect 27522 21428 27528 21480
rect 27580 21468 27586 21480
rect 27632 21468 27660 21576
rect 29549 21573 29561 21576
rect 29595 21573 29607 21607
rect 29549 21567 29607 21573
rect 28810 21496 28816 21548
rect 28868 21536 28874 21548
rect 29273 21539 29331 21545
rect 29273 21536 29285 21539
rect 28868 21508 29285 21536
rect 28868 21496 28874 21508
rect 29273 21505 29285 21508
rect 29319 21505 29331 21539
rect 29273 21499 29331 21505
rect 27580 21440 27660 21468
rect 27580 21428 27586 21440
rect 27706 21428 27712 21480
rect 27764 21428 27770 21480
rect 28074 21428 28080 21480
rect 28132 21428 28138 21480
rect 28994 21428 29000 21480
rect 29052 21428 29058 21480
rect 29178 21477 29184 21480
rect 29135 21471 29184 21477
rect 29135 21437 29147 21471
rect 29181 21437 29184 21471
rect 29135 21431 29184 21437
rect 29178 21428 29184 21431
rect 29236 21428 29242 21480
rect 29457 21471 29515 21477
rect 29457 21437 29469 21471
rect 29503 21437 29515 21471
rect 29457 21431 29515 21437
rect 23952 21372 24256 21400
rect 24397 21403 24455 21409
rect 19610 21332 19616 21344
rect 18892 21304 19616 21332
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 23952 21341 23980 21372
rect 24397 21369 24409 21403
rect 24443 21400 24455 21403
rect 24443 21372 25360 21400
rect 24443 21369 24455 21372
rect 24397 21363 24455 21369
rect 21361 21335 21419 21341
rect 21361 21332 21373 21335
rect 20680 21304 21373 21332
rect 20680 21292 20686 21304
rect 21361 21301 21373 21304
rect 21407 21301 21419 21335
rect 21361 21295 21419 21301
rect 23937 21335 23995 21341
rect 23937 21301 23949 21335
rect 23983 21301 23995 21335
rect 23937 21295 23995 21301
rect 24118 21292 24124 21344
rect 24176 21292 24182 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24854 21332 24860 21344
rect 24268 21304 24860 21332
rect 24268 21292 24274 21304
rect 24854 21292 24860 21304
rect 24912 21292 24918 21344
rect 25332 21341 25360 21372
rect 26326 21360 26332 21412
rect 26384 21400 26390 21412
rect 27157 21403 27215 21409
rect 27157 21400 27169 21403
rect 26384 21372 27169 21400
rect 26384 21360 26390 21372
rect 27157 21369 27169 21372
rect 27203 21400 27215 21403
rect 29472 21400 29500 21431
rect 29730 21428 29736 21480
rect 29788 21428 29794 21480
rect 30006 21428 30012 21480
rect 30064 21428 30070 21480
rect 30282 21428 30288 21480
rect 30340 21468 30346 21480
rect 30469 21471 30527 21477
rect 30469 21468 30481 21471
rect 30340 21440 30481 21468
rect 30340 21428 30346 21440
rect 30469 21437 30481 21440
rect 30515 21437 30527 21471
rect 30469 21431 30527 21437
rect 29638 21400 29644 21412
rect 27203 21372 29644 21400
rect 27203 21369 27215 21372
rect 27157 21363 27215 21369
rect 29638 21360 29644 21372
rect 29696 21360 29702 21412
rect 25317 21335 25375 21341
rect 25317 21301 25329 21335
rect 25363 21301 25375 21335
rect 25317 21295 25375 21301
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 27246 21292 27252 21344
rect 27304 21292 27310 21344
rect 28261 21335 28319 21341
rect 28261 21301 28273 21335
rect 28307 21332 28319 21335
rect 28994 21332 29000 21344
rect 28307 21304 29000 21332
rect 28307 21301 28319 21304
rect 28261 21295 28319 21301
rect 28994 21292 29000 21304
rect 29052 21292 29058 21344
rect 29362 21292 29368 21344
rect 29420 21292 29426 21344
rect 30282 21292 30288 21344
rect 30340 21292 30346 21344
rect 552 21242 31808 21264
rect 552 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 15946 21242
rect 15998 21190 16010 21242
rect 16062 21190 16074 21242
rect 16126 21190 16138 21242
rect 16190 21190 16202 21242
rect 16254 21190 23720 21242
rect 23772 21190 23784 21242
rect 23836 21190 23848 21242
rect 23900 21190 23912 21242
rect 23964 21190 23976 21242
rect 24028 21190 31494 21242
rect 31546 21190 31558 21242
rect 31610 21190 31622 21242
rect 31674 21190 31686 21242
rect 31738 21190 31750 21242
rect 31802 21190 31808 21242
rect 552 21168 31808 21190
rect 2130 21088 2136 21140
rect 2188 21128 2194 21140
rect 3513 21131 3571 21137
rect 2188 21100 2452 21128
rect 2188 21088 2194 21100
rect 2424 21060 2452 21100
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 3878 21128 3884 21140
rect 3559 21100 3884 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 3970 21088 3976 21140
rect 4028 21088 4034 21140
rect 4062 21088 4068 21140
rect 4120 21088 4126 21140
rect 4617 21131 4675 21137
rect 4617 21097 4629 21131
rect 4663 21097 4675 21131
rect 4617 21091 4675 21097
rect 2869 21063 2927 21069
rect 2869 21060 2881 21063
rect 2424 21032 2881 21060
rect 2869 21029 2881 21032
rect 2915 21029 2927 21063
rect 4632 21060 4660 21091
rect 4982 21088 4988 21140
rect 5040 21088 5046 21140
rect 5074 21088 5080 21140
rect 5132 21088 5138 21140
rect 6454 21088 6460 21140
rect 6512 21088 6518 21140
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 6825 21131 6883 21137
rect 6825 21128 6837 21131
rect 6696 21100 6837 21128
rect 6696 21088 6702 21100
rect 6825 21097 6837 21100
rect 6871 21097 6883 21131
rect 8938 21128 8944 21140
rect 6825 21091 6883 21097
rect 8772 21100 8944 21128
rect 2869 21023 2927 21029
rect 3344 21032 4660 21060
rect 2222 20952 2228 21004
rect 2280 20952 2286 21004
rect 3344 21001 3372 21032
rect 4706 21020 4712 21072
rect 4764 21060 4770 21072
rect 7006 21060 7012 21072
rect 4764 21032 7012 21060
rect 4764 21020 4770 21032
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 8772 21069 8800 21100
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 9030 21088 9036 21140
rect 9088 21088 9094 21140
rect 9398 21088 9404 21140
rect 9456 21128 9462 21140
rect 10045 21131 10103 21137
rect 10045 21128 10057 21131
rect 9456 21100 10057 21128
rect 9456 21088 9462 21100
rect 10045 21097 10057 21100
rect 10091 21097 10103 21131
rect 13078 21128 13084 21140
rect 10045 21091 10103 21097
rect 11072 21100 13084 21128
rect 8757 21063 8815 21069
rect 8757 21029 8769 21063
rect 8803 21029 8815 21063
rect 9048 21060 9076 21088
rect 9585 21063 9643 21069
rect 9585 21060 9597 21063
rect 9048 21032 9597 21060
rect 8757 21023 8815 21029
rect 9585 21029 9597 21032
rect 9631 21029 9643 21063
rect 9585 21023 9643 21029
rect 9677 21063 9735 21069
rect 9677 21029 9689 21063
rect 9723 21060 9735 21063
rect 11072 21060 11100 21100
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13722 21128 13728 21140
rect 13780 21137 13786 21140
rect 13780 21131 13799 21137
rect 13228 21100 13728 21128
rect 13228 21088 13234 21100
rect 13722 21088 13728 21100
rect 13787 21097 13799 21131
rect 13780 21091 13799 21097
rect 13909 21131 13967 21137
rect 13909 21097 13921 21131
rect 13955 21128 13967 21131
rect 14366 21128 14372 21140
rect 13955 21100 14372 21128
rect 13955 21097 13967 21100
rect 13909 21091 13967 21097
rect 13780 21088 13786 21091
rect 14366 21088 14372 21100
rect 14424 21088 14430 21140
rect 15746 21088 15752 21140
rect 15804 21088 15810 21140
rect 15856 21100 18000 21128
rect 9723 21032 11100 21060
rect 11164 21032 11468 21060
rect 9723 21029 9735 21032
rect 9677 21023 9735 21029
rect 3053 20995 3111 21001
rect 3053 20961 3065 20995
rect 3099 20961 3111 20995
rect 3053 20955 3111 20961
rect 3329 20995 3387 21001
rect 3329 20961 3341 20995
rect 3375 20961 3387 20995
rect 3329 20955 3387 20961
rect 3804 20964 5212 20992
rect 845 20927 903 20933
rect 845 20893 857 20927
rect 891 20924 903 20927
rect 1121 20927 1179 20933
rect 891 20896 980 20924
rect 891 20893 903 20896
rect 845 20887 903 20893
rect 952 20800 980 20896
rect 1121 20893 1133 20927
rect 1167 20924 1179 20927
rect 1210 20924 1216 20936
rect 1167 20896 1216 20924
rect 1167 20893 1179 20896
rect 1121 20887 1179 20893
rect 1210 20884 1216 20896
rect 1268 20884 1274 20936
rect 3068 20924 3096 20955
rect 3804 20936 3832 20964
rect 3068 20896 3648 20924
rect 3620 20865 3648 20896
rect 3786 20884 3792 20936
rect 3844 20884 3850 20936
rect 4172 20933 4200 20964
rect 5184 20933 5212 20964
rect 5442 20952 5448 21004
rect 5500 20952 5506 21004
rect 5810 20952 5816 21004
rect 5868 20952 5874 21004
rect 6365 20995 6423 21001
rect 6365 20961 6377 20995
rect 6411 20961 6423 20995
rect 6365 20955 6423 20961
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 6181 20927 6239 20933
rect 6181 20924 6193 20927
rect 5215 20896 6193 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 6181 20893 6193 20896
rect 6227 20924 6239 20927
rect 6270 20924 6276 20936
rect 6227 20896 6276 20924
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6270 20884 6276 20896
rect 6328 20884 6334 20936
rect 3605 20859 3663 20865
rect 3605 20825 3617 20859
rect 3651 20825 3663 20859
rect 3605 20819 3663 20825
rect 934 20748 940 20800
rect 992 20748 998 20800
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 5626 20748 5632 20800
rect 5684 20748 5690 20800
rect 5997 20791 6055 20797
rect 5997 20757 6009 20791
rect 6043 20788 6055 20791
rect 6086 20788 6092 20800
rect 6043 20760 6092 20788
rect 6043 20757 6055 20760
rect 5997 20751 6055 20757
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6380 20788 6408 20955
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 6972 20964 7682 20992
rect 6972 20952 6978 20964
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 10376 20964 10425 20992
rect 10376 20952 10382 20964
rect 10413 20961 10425 20964
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 10594 20992 10600 21004
rect 10551 20964 10600 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 11164 20992 11192 21032
rect 10836 20964 11192 20992
rect 10836 20952 10842 20964
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11333 20995 11391 21001
rect 11333 20992 11345 20995
rect 11296 20964 11345 20992
rect 11296 20952 11302 20964
rect 11333 20961 11345 20964
rect 11379 20961 11391 20995
rect 11440 20992 11468 21032
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 13541 21063 13599 21069
rect 13541 21060 13553 21063
rect 12308 21032 13553 21060
rect 12308 21020 12314 21032
rect 13541 21029 13553 21032
rect 13587 21060 13599 21063
rect 14734 21060 14740 21072
rect 13587 21032 14740 21060
rect 13587 21029 13599 21032
rect 13541 21023 13599 21029
rect 14734 21020 14740 21032
rect 14792 21020 14798 21072
rect 15856 21060 15884 21100
rect 17972 21072 18000 21100
rect 18506 21088 18512 21140
rect 18564 21088 18570 21140
rect 19058 21088 19064 21140
rect 19116 21088 19122 21140
rect 19242 21137 19248 21140
rect 19229 21131 19248 21137
rect 19229 21097 19241 21131
rect 19229 21091 19248 21097
rect 19242 21088 19248 21091
rect 19300 21088 19306 21140
rect 20530 21128 20536 21140
rect 19352 21100 20536 21128
rect 15626 21032 15884 21060
rect 15626 21004 15654 21032
rect 16022 21020 16028 21072
rect 16080 21060 16086 21072
rect 16393 21063 16451 21069
rect 16393 21060 16405 21063
rect 16080 21032 16405 21060
rect 16080 21020 16086 21032
rect 16393 21029 16405 21032
rect 16439 21060 16451 21063
rect 16439 21032 16620 21060
rect 16439 21029 16451 21032
rect 16393 21023 16451 21029
rect 12342 20992 12348 21004
rect 11440 20964 12348 20992
rect 11333 20955 11391 20961
rect 12342 20952 12348 20964
rect 12400 20992 12406 21004
rect 12437 20995 12495 21001
rect 12437 20992 12449 20995
rect 12400 20964 12449 20992
rect 12400 20952 12406 20964
rect 12437 20961 12449 20964
rect 12483 20961 12495 20995
rect 12437 20955 12495 20961
rect 12529 20995 12587 21001
rect 12529 20961 12541 20995
rect 12575 20992 12587 20995
rect 12802 20992 12808 21004
rect 12575 20964 12808 20992
rect 12575 20961 12587 20964
rect 12529 20955 12587 20961
rect 12802 20952 12808 20964
rect 12860 20952 12866 21004
rect 13262 20952 13268 21004
rect 13320 20952 13326 21004
rect 13906 20952 13912 21004
rect 13964 20952 13970 21004
rect 14090 20952 14096 21004
rect 14148 20992 14154 21004
rect 14185 20995 14243 21001
rect 14185 20992 14197 20995
rect 14148 20964 14197 20992
rect 14148 20952 14154 20964
rect 14185 20961 14197 20964
rect 14231 20961 14243 20995
rect 14185 20955 14243 20961
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 14700 20964 15117 20992
rect 14700 20952 14706 20964
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 15194 20952 15200 21004
rect 15252 20992 15258 21004
rect 15252 20964 15297 20992
rect 15252 20952 15258 20964
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 15626 21001 15660 21004
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20961 15531 20995
rect 15473 20955 15531 20961
rect 15611 20995 15660 21001
rect 15611 20961 15623 20995
rect 15657 20961 15660 20995
rect 15611 20955 15660 20961
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7340 20896 8984 20924
rect 7340 20884 7346 20896
rect 8956 20856 8984 20896
rect 9030 20884 9036 20936
rect 9088 20884 9094 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9732 20896 9873 20924
rect 9732 20884 9738 20896
rect 9861 20893 9873 20896
rect 9907 20924 9919 20927
rect 9950 20924 9956 20936
rect 9907 20896 9956 20924
rect 9907 20893 9919 20896
rect 9861 20887 9919 20893
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10689 20927 10747 20933
rect 10689 20924 10701 20927
rect 10008 20896 10701 20924
rect 10008 20884 10014 20896
rect 10689 20893 10701 20896
rect 10735 20924 10747 20927
rect 10735 20896 11008 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 8956 20828 9229 20856
rect 9217 20825 9229 20828
rect 9263 20825 9275 20859
rect 9217 20819 9275 20825
rect 9766 20816 9772 20868
rect 9824 20856 9830 20868
rect 10870 20856 10876 20868
rect 9824 20828 10876 20856
rect 9824 20816 9830 20828
rect 10870 20816 10876 20828
rect 10928 20816 10934 20868
rect 10980 20856 11008 20896
rect 11422 20884 11428 20936
rect 11480 20884 11486 20936
rect 11514 20884 11520 20936
rect 11572 20924 11578 20936
rect 12621 20927 12679 20933
rect 12621 20924 12633 20927
rect 11572 20896 12633 20924
rect 11572 20884 11578 20896
rect 12621 20893 12633 20896
rect 12667 20893 12679 20927
rect 12621 20887 12679 20893
rect 13078 20884 13084 20936
rect 13136 20924 13142 20936
rect 13814 20924 13820 20936
rect 13136 20896 13820 20924
rect 13136 20884 13142 20896
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 13924 20924 13952 20952
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 13924 20896 14473 20924
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 15488 20924 15516 20955
rect 15654 20952 15660 20955
rect 15712 20952 15718 21004
rect 15838 20952 15844 21004
rect 15896 20992 15902 21004
rect 16117 20995 16175 21001
rect 16117 20992 16129 20995
rect 15896 20964 16129 20992
rect 15896 20952 15902 20964
rect 16117 20961 16129 20964
rect 16163 20961 16175 20995
rect 16117 20955 16175 20961
rect 16298 20952 16304 21004
rect 16356 20952 16362 21004
rect 16482 20952 16488 21004
rect 16540 20952 16546 21004
rect 16592 20992 16620 21032
rect 16666 21020 16672 21072
rect 16724 21020 16730 21072
rect 17954 21020 17960 21072
rect 18012 21060 18018 21072
rect 19352 21060 19380 21100
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 21545 21131 21603 21137
rect 21545 21097 21557 21131
rect 21591 21128 21603 21131
rect 21591 21100 22324 21128
rect 21591 21097 21603 21100
rect 21545 21091 21603 21097
rect 18012 21032 19380 21060
rect 18012 21020 18018 21032
rect 19426 21020 19432 21072
rect 19484 21060 19490 21072
rect 19484 21032 20852 21060
rect 19484 21020 19490 21032
rect 18230 20992 18236 21004
rect 16592 20964 18236 20992
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 18322 20952 18328 21004
rect 18380 20952 18386 21004
rect 18723 20995 18781 21001
rect 18723 20992 18735 20995
rect 18708 20961 18735 20992
rect 18769 20961 18781 20995
rect 18708 20955 18781 20961
rect 20165 20995 20223 21001
rect 20165 20961 20177 20995
rect 20211 20961 20223 20995
rect 20165 20955 20223 20961
rect 16390 20924 16396 20936
rect 15488 20896 16396 20924
rect 11532 20856 11560 20884
rect 10980 20828 11560 20856
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 15488 20856 15516 20896
rect 16390 20884 16396 20896
rect 16448 20924 16454 20936
rect 18340 20924 18368 20952
rect 16448 20896 18368 20924
rect 16448 20884 16454 20896
rect 12032 20828 15516 20856
rect 12032 20816 12038 20828
rect 10778 20788 10784 20800
rect 6380 20760 10784 20788
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 10962 20748 10968 20800
rect 11020 20748 11026 20800
rect 11606 20748 11612 20800
rect 11664 20788 11670 20800
rect 12069 20791 12127 20797
rect 12069 20788 12081 20791
rect 11664 20760 12081 20788
rect 11664 20748 11670 20760
rect 12069 20757 12081 20760
rect 12115 20757 12127 20791
rect 12069 20751 12127 20757
rect 12388 20748 12394 20800
rect 12446 20788 12452 20800
rect 12989 20791 13047 20797
rect 12989 20788 13001 20791
rect 12446 20760 13001 20788
rect 12446 20748 12452 20760
rect 12989 20757 13001 20760
rect 13035 20757 13047 20791
rect 12989 20751 13047 20757
rect 13722 20748 13728 20800
rect 13780 20748 13786 20800
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 18708 20788 18736 20955
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 18969 20927 19027 20933
rect 18969 20893 18981 20927
rect 19015 20924 19027 20927
rect 19058 20924 19064 20936
rect 19015 20896 19064 20924
rect 19015 20893 19027 20896
rect 18969 20887 19027 20893
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 20180 20856 20208 20955
rect 20254 20952 20260 21004
rect 20312 20952 20318 21004
rect 20349 20995 20407 21001
rect 20349 20961 20361 20995
rect 20395 20982 20407 20995
rect 20714 20992 20720 21004
rect 20640 20982 20720 20992
rect 20395 20964 20720 20982
rect 20395 20961 20668 20964
rect 20349 20955 20668 20961
rect 20364 20954 20668 20955
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 20824 20992 20852 21032
rect 21450 21020 21456 21072
rect 21508 21060 21514 21072
rect 22296 21060 22324 21100
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 22428 21100 24075 21128
rect 22428 21088 22434 21100
rect 22462 21060 22468 21072
rect 21508 21032 21956 21060
rect 22296 21032 22468 21060
rect 21508 21020 21514 21032
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 20824 20964 21649 20992
rect 21637 20961 21649 20964
rect 21683 20992 21695 20995
rect 21818 20992 21824 21004
rect 21683 20964 21824 20992
rect 21683 20961 21695 20964
rect 21637 20955 21695 20961
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 21928 20992 21956 21032
rect 22462 21020 22468 21032
rect 22520 21020 22526 21072
rect 23842 21060 23848 21072
rect 22572 21032 23848 21060
rect 22572 21001 22600 21032
rect 23842 21020 23848 21032
rect 23900 21020 23906 21072
rect 24047 21060 24075 21100
rect 24118 21088 24124 21140
rect 24176 21128 24182 21140
rect 24305 21131 24363 21137
rect 24305 21128 24317 21131
rect 24176 21100 24317 21128
rect 24176 21088 24182 21100
rect 24305 21097 24317 21100
rect 24351 21097 24363 21131
rect 24305 21091 24363 21097
rect 25148 21100 26832 21128
rect 25148 21060 25176 21100
rect 24047 21032 25176 21060
rect 25240 21032 26740 21060
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 21928 20964 22569 20992
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20961 22799 20995
rect 22741 20955 22799 20961
rect 20732 20924 20760 20952
rect 22370 20924 22376 20936
rect 20732 20896 22376 20924
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22756 20924 22784 20955
rect 22830 20952 22836 21004
rect 22888 20952 22894 21004
rect 22922 20952 22928 21004
rect 22980 20952 22986 21004
rect 23290 20952 23296 21004
rect 23348 20952 23354 21004
rect 23382 20952 23388 21004
rect 23440 20992 23446 21004
rect 23477 20995 23535 21001
rect 23477 20992 23489 20995
rect 23440 20964 23489 20992
rect 23440 20952 23446 20964
rect 23477 20961 23489 20964
rect 23523 20961 23535 20995
rect 23477 20955 23535 20961
rect 23566 20952 23572 21004
rect 23624 20952 23630 21004
rect 24486 20952 24492 21004
rect 24544 20952 24550 21004
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 24627 20964 24961 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24949 20961 24961 20964
rect 24995 20961 25007 20995
rect 24949 20955 25007 20961
rect 25130 20952 25136 21004
rect 25188 20952 25194 21004
rect 23658 20924 23664 20936
rect 22756 20896 23664 20924
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 23768 20896 24685 20924
rect 21821 20859 21879 20865
rect 21821 20856 21833 20859
rect 19392 20828 21833 20856
rect 19392 20816 19398 20828
rect 21821 20825 21833 20828
rect 21867 20825 21879 20859
rect 21821 20819 21879 20825
rect 21910 20816 21916 20868
rect 21968 20856 21974 20868
rect 23768 20865 23796 20896
rect 24673 20893 24685 20896
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 25240 20924 25268 21032
rect 26712 21004 26740 21032
rect 25314 20952 25320 21004
rect 25372 20952 25378 21004
rect 25406 20952 25412 21004
rect 25464 20952 25470 21004
rect 25498 20952 25504 21004
rect 25556 20952 25562 21004
rect 25682 20952 25688 21004
rect 25740 20952 25746 21004
rect 25774 20952 25780 21004
rect 25832 20952 25838 21004
rect 26513 20995 26571 21001
rect 26513 20961 26525 20995
rect 26559 20961 26571 20995
rect 26513 20955 26571 20961
rect 24811 20896 25268 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 23753 20859 23811 20865
rect 21968 20828 23704 20856
rect 21968 20816 21974 20828
rect 17368 20760 18736 20788
rect 17368 20748 17374 20760
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 19245 20791 19303 20797
rect 19245 20788 19257 20791
rect 18840 20760 19257 20788
rect 18840 20748 18846 20760
rect 19245 20757 19257 20760
rect 19291 20757 19303 20791
rect 19245 20751 19303 20757
rect 21266 20748 21272 20800
rect 21324 20748 21330 20800
rect 23201 20791 23259 20797
rect 23201 20757 23213 20791
rect 23247 20788 23259 20791
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 23247 20760 23305 20788
rect 23247 20757 23259 20760
rect 23201 20751 23259 20757
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23676 20788 23704 20828
rect 23753 20825 23765 20859
rect 23799 20825 23811 20859
rect 23753 20819 23811 20825
rect 23842 20816 23848 20868
rect 23900 20856 23906 20868
rect 25332 20856 25360 20952
rect 23900 20828 25360 20856
rect 25424 20856 25452 20952
rect 26528 20924 26556 20955
rect 26694 20952 26700 21004
rect 26752 20952 26758 21004
rect 26804 20992 26832 21100
rect 26878 21088 26884 21140
rect 26936 21128 26942 21140
rect 28077 21131 28135 21137
rect 26936 21100 27660 21128
rect 26936 21088 26942 21100
rect 27062 21020 27068 21072
rect 27120 21060 27126 21072
rect 27338 21060 27344 21072
rect 27120 21032 27344 21060
rect 27120 21020 27126 21032
rect 27338 21020 27344 21032
rect 27396 21020 27402 21072
rect 27632 21069 27660 21100
rect 28077 21097 28089 21131
rect 28123 21097 28135 21131
rect 28077 21091 28135 21097
rect 27617 21063 27675 21069
rect 27617 21029 27629 21063
rect 27663 21029 27675 21063
rect 27617 21023 27675 21029
rect 27709 21063 27767 21069
rect 27709 21029 27721 21063
rect 27755 21060 27767 21063
rect 28092 21060 28120 21091
rect 29178 21088 29184 21140
rect 29236 21128 29242 21140
rect 30101 21131 30159 21137
rect 30101 21128 30113 21131
rect 29236 21100 30113 21128
rect 29236 21088 29242 21100
rect 30101 21097 30113 21100
rect 30147 21097 30159 21131
rect 30101 21091 30159 21097
rect 30834 21088 30840 21140
rect 30892 21088 30898 21140
rect 29086 21060 29092 21072
rect 27755 21032 28120 21060
rect 28368 21032 29092 21060
rect 27755 21029 27767 21032
rect 27709 21023 27767 21029
rect 27479 20995 27537 21001
rect 27479 20992 27491 20995
rect 26804 20964 27491 20992
rect 27479 20961 27491 20964
rect 27525 20992 27537 20995
rect 27798 20992 27804 21004
rect 27525 20964 27804 20992
rect 27525 20961 27537 20964
rect 27479 20955 27537 20961
rect 27798 20952 27804 20964
rect 27856 20952 27862 21004
rect 27890 20952 27896 21004
rect 27948 20952 27954 21004
rect 27985 20995 28043 21001
rect 27985 20961 27997 20995
rect 28031 20992 28043 20995
rect 28368 20992 28396 21032
rect 29086 21020 29092 21032
rect 29144 21020 29150 21072
rect 28031 20964 28396 20992
rect 28445 20995 28503 21001
rect 28031 20961 28043 20964
rect 27985 20955 28043 20961
rect 28445 20961 28457 20995
rect 28491 20961 28503 20995
rect 28445 20955 28503 20961
rect 25608 20896 26556 20924
rect 26605 20927 26663 20933
rect 25608 20868 25636 20896
rect 26605 20893 26617 20927
rect 26651 20924 26663 20927
rect 28000 20924 28028 20955
rect 26651 20896 28028 20924
rect 26651 20893 26663 20896
rect 26605 20887 26663 20893
rect 28350 20884 28356 20936
rect 28408 20884 28414 20936
rect 28460 20924 28488 20955
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 30285 20995 30343 21001
rect 30285 20992 30297 20995
rect 28592 20964 30297 20992
rect 28592 20952 28598 20964
rect 30285 20961 30297 20964
rect 30331 20961 30343 20995
rect 30285 20955 30343 20961
rect 30745 20995 30803 21001
rect 30745 20961 30757 20995
rect 30791 20992 30803 20995
rect 30926 20992 30932 21004
rect 30791 20964 30932 20992
rect 30791 20961 30803 20964
rect 30745 20955 30803 20961
rect 30926 20952 30932 20964
rect 30984 20952 30990 21004
rect 30558 20924 30564 20936
rect 28460 20896 30564 20924
rect 25501 20859 25559 20865
rect 25501 20856 25513 20859
rect 25424 20828 25513 20856
rect 23900 20816 23906 20828
rect 25501 20825 25513 20828
rect 25547 20825 25559 20859
rect 25501 20819 25559 20825
rect 25590 20816 25596 20868
rect 25648 20816 25654 20868
rect 28460 20856 28488 20896
rect 30558 20884 30564 20896
rect 30616 20884 30622 20936
rect 27264 20828 28488 20856
rect 27264 20788 27292 20828
rect 23676 20760 27292 20788
rect 23293 20751 23351 20757
rect 27338 20748 27344 20800
rect 27396 20748 27402 20800
rect 27798 20748 27804 20800
rect 27856 20788 27862 20800
rect 28074 20788 28080 20800
rect 27856 20760 28080 20788
rect 27856 20748 27862 20760
rect 28074 20748 28080 20760
rect 28132 20788 28138 20800
rect 28261 20791 28319 20797
rect 28261 20788 28273 20791
rect 28132 20760 28273 20788
rect 28132 20748 28138 20760
rect 28261 20757 28273 20760
rect 28307 20757 28319 20791
rect 28261 20751 28319 20757
rect 30466 20748 30472 20800
rect 30524 20748 30530 20800
rect 552 20698 31648 20720
rect 552 20646 4285 20698
rect 4337 20646 4349 20698
rect 4401 20646 4413 20698
rect 4465 20646 4477 20698
rect 4529 20646 4541 20698
rect 4593 20646 12059 20698
rect 12111 20646 12123 20698
rect 12175 20646 12187 20698
rect 12239 20646 12251 20698
rect 12303 20646 12315 20698
rect 12367 20646 19833 20698
rect 19885 20646 19897 20698
rect 19949 20646 19961 20698
rect 20013 20646 20025 20698
rect 20077 20646 20089 20698
rect 20141 20646 27607 20698
rect 27659 20646 27671 20698
rect 27723 20646 27735 20698
rect 27787 20646 27799 20698
rect 27851 20646 27863 20698
rect 27915 20646 31648 20698
rect 552 20624 31648 20646
rect 2682 20544 2688 20596
rect 2740 20584 2746 20596
rect 2869 20587 2927 20593
rect 2869 20584 2881 20587
rect 2740 20556 2881 20584
rect 2740 20544 2746 20556
rect 2869 20553 2881 20556
rect 2915 20553 2927 20587
rect 4614 20584 4620 20596
rect 2869 20547 2927 20553
rect 3068 20556 4620 20584
rect 1688 20488 3004 20516
rect 937 20383 995 20389
rect 937 20349 949 20383
rect 983 20380 995 20383
rect 983 20352 1256 20380
rect 983 20349 995 20352
rect 937 20343 995 20349
rect 1118 20204 1124 20256
rect 1176 20204 1182 20256
rect 1228 20253 1256 20352
rect 1578 20340 1584 20392
rect 1636 20340 1642 20392
rect 1688 20389 1716 20488
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20417 1915 20451
rect 1857 20411 1915 20417
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20349 1731 20383
rect 1872 20380 1900 20411
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2556 20420 2605 20448
rect 2556 20408 2562 20420
rect 2593 20417 2605 20420
rect 2639 20417 2651 20451
rect 2593 20411 2651 20417
rect 2866 20380 2872 20392
rect 1872 20352 2872 20380
rect 1673 20343 1731 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 2409 20315 2467 20321
rect 2409 20281 2421 20315
rect 2455 20312 2467 20315
rect 2774 20312 2780 20324
rect 2455 20284 2780 20312
rect 2455 20281 2467 20284
rect 2409 20275 2467 20281
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 1213 20247 1271 20253
rect 1213 20213 1225 20247
rect 1259 20213 1271 20247
rect 1213 20207 1271 20213
rect 2038 20204 2044 20256
rect 2096 20204 2102 20256
rect 2501 20247 2559 20253
rect 2501 20213 2513 20247
rect 2547 20244 2559 20247
rect 2590 20244 2596 20256
rect 2547 20216 2596 20244
rect 2547 20213 2559 20216
rect 2501 20207 2559 20213
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 2976 20244 3004 20488
rect 3068 20389 3096 20556
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 5276 20556 7972 20584
rect 4522 20476 4528 20528
rect 4580 20516 4586 20528
rect 5276 20516 5304 20556
rect 4580 20488 5304 20516
rect 4580 20476 4586 20488
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3602 20448 3608 20460
rect 3283 20420 3608 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 5261 20451 5319 20457
rect 5261 20448 5273 20451
rect 4212 20420 5273 20448
rect 4212 20408 4218 20420
rect 5261 20417 5273 20420
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 7190 20408 7196 20460
rect 7248 20448 7254 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 7248 20420 7297 20448
rect 7248 20408 7254 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 7944 20448 7972 20556
rect 8662 20544 8668 20596
rect 8720 20544 8726 20596
rect 10502 20544 10508 20596
rect 10560 20544 10566 20596
rect 11057 20587 11115 20593
rect 11057 20553 11069 20587
rect 11103 20584 11115 20587
rect 11790 20584 11796 20596
rect 11103 20556 11796 20584
rect 11103 20553 11115 20556
rect 11057 20547 11115 20553
rect 11790 20544 11796 20556
rect 11848 20544 11854 20596
rect 13998 20584 14004 20596
rect 11900 20556 14004 20584
rect 8018 20476 8024 20528
rect 8076 20516 8082 20528
rect 8941 20519 8999 20525
rect 8941 20516 8953 20519
rect 8076 20488 8953 20516
rect 8076 20476 8082 20488
rect 8941 20485 8953 20488
rect 8987 20485 8999 20519
rect 11900 20516 11928 20556
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 15286 20584 15292 20596
rect 14139 20556 15292 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20584 15623 20587
rect 16022 20584 16028 20596
rect 15611 20556 16028 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 16298 20544 16304 20596
rect 16356 20544 16362 20596
rect 17865 20587 17923 20593
rect 17865 20553 17877 20587
rect 17911 20584 17923 20587
rect 17954 20584 17960 20596
rect 17911 20556 17960 20584
rect 17911 20553 17923 20556
rect 17865 20547 17923 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 18288 20556 20668 20584
rect 18288 20544 18294 20556
rect 8941 20479 8999 20485
rect 10888 20488 11928 20516
rect 9585 20451 9643 20457
rect 7944 20420 9536 20448
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20380 7619 20383
rect 8757 20383 8815 20389
rect 7607 20352 8064 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 3234 20272 3240 20324
rect 3292 20312 3298 20324
rect 3513 20315 3571 20321
rect 3513 20312 3525 20315
rect 3292 20284 3525 20312
rect 3292 20272 3298 20284
rect 3513 20281 3525 20284
rect 3559 20281 3571 20315
rect 4982 20312 4988 20324
rect 4738 20284 4988 20312
rect 3513 20275 3571 20281
rect 4982 20272 4988 20284
rect 5040 20272 5046 20324
rect 5537 20315 5595 20321
rect 5537 20281 5549 20315
rect 5583 20281 5595 20315
rect 6854 20284 6960 20312
rect 5537 20275 5595 20281
rect 4154 20244 4160 20256
rect 2976 20216 4160 20244
rect 4154 20204 4160 20216
rect 4212 20244 4218 20256
rect 4522 20244 4528 20256
rect 4212 20216 4528 20244
rect 4212 20204 4218 20216
rect 4522 20204 4528 20216
rect 4580 20204 4586 20256
rect 5552 20244 5580 20275
rect 6932 20256 6960 20284
rect 6454 20244 6460 20256
rect 5552 20216 6460 20244
rect 6454 20204 6460 20216
rect 6512 20204 6518 20256
rect 6914 20204 6920 20256
rect 6972 20204 6978 20256
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 8036 20244 8064 20352
rect 8757 20349 8769 20383
rect 8803 20380 8815 20383
rect 9398 20380 9404 20392
rect 8803 20352 9404 20380
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 8113 20315 8171 20321
rect 8113 20281 8125 20315
rect 8159 20312 8171 20315
rect 8846 20312 8852 20324
rect 8159 20284 8852 20312
rect 8159 20281 8171 20284
rect 8113 20275 8171 20281
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 9030 20272 9036 20324
rect 9088 20272 9094 20324
rect 9309 20315 9367 20321
rect 9309 20281 9321 20315
rect 9355 20312 9367 20315
rect 9508 20312 9536 20420
rect 9585 20417 9597 20451
rect 9631 20448 9643 20451
rect 9950 20448 9956 20460
rect 9631 20420 9956 20448
rect 9631 20417 9643 20420
rect 9585 20411 9643 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10778 20448 10784 20460
rect 10091 20420 10784 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 10888 20380 10916 20488
rect 13814 20476 13820 20528
rect 13872 20516 13878 20528
rect 16574 20516 16580 20528
rect 13872 20488 16580 20516
rect 13872 20476 13878 20488
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 16853 20519 16911 20525
rect 16853 20485 16865 20519
rect 16899 20516 16911 20519
rect 17681 20519 17739 20525
rect 16899 20488 17264 20516
rect 16899 20485 16911 20488
rect 16853 20479 16911 20485
rect 11379 20451 11437 20457
rect 11379 20417 11391 20451
rect 11425 20448 11437 20451
rect 12986 20448 12992 20460
rect 11425 20420 12992 20448
rect 11425 20417 11437 20420
rect 11379 20411 11437 20417
rect 12986 20408 12992 20420
rect 13044 20448 13050 20460
rect 15746 20448 15752 20460
rect 13044 20420 13584 20448
rect 13044 20408 13050 20420
rect 9355 20284 9536 20312
rect 9968 20352 10916 20380
rect 11149 20383 11207 20389
rect 9355 20281 9367 20284
rect 9309 20275 9367 20281
rect 8570 20244 8576 20256
rect 7892 20216 8576 20244
rect 7892 20204 7898 20216
rect 8570 20204 8576 20216
rect 8628 20244 8634 20256
rect 9048 20244 9076 20272
rect 8628 20216 9076 20244
rect 9401 20247 9459 20253
rect 8628 20204 8634 20216
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 9968 20244 9996 20352
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11606 20380 11612 20392
rect 11195 20352 11612 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11606 20340 11612 20352
rect 11664 20340 11670 20392
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20380 12863 20383
rect 12894 20380 12900 20392
rect 12851 20352 12900 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 13170 20340 13176 20392
rect 13228 20340 13234 20392
rect 13556 20389 13584 20420
rect 14476 20420 15752 20448
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 14182 20340 14188 20392
rect 14240 20380 14246 20392
rect 14277 20383 14335 20389
rect 14277 20380 14289 20383
rect 14240 20352 14289 20380
rect 14240 20340 14246 20352
rect 14277 20349 14289 20352
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 14366 20340 14372 20392
rect 14424 20340 14430 20392
rect 12250 20272 12256 20324
rect 12308 20272 12314 20324
rect 13633 20315 13691 20321
rect 13633 20281 13645 20315
rect 13679 20312 13691 20315
rect 14476 20312 14504 20420
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 14734 20340 14740 20392
rect 14792 20340 14798 20392
rect 14826 20340 14832 20392
rect 14884 20340 14890 20392
rect 15010 20340 15016 20392
rect 15068 20340 15074 20392
rect 15102 20340 15108 20392
rect 15160 20380 15166 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15160 20352 15485 20380
rect 15160 20340 15166 20352
rect 15473 20349 15485 20352
rect 15519 20380 15531 20383
rect 15562 20380 15568 20392
rect 15519 20352 15568 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 15654 20340 15660 20392
rect 15712 20340 15718 20392
rect 15930 20340 15936 20392
rect 15988 20340 15994 20392
rect 16393 20383 16451 20389
rect 16393 20349 16405 20383
rect 16439 20380 16451 20383
rect 16482 20380 16488 20392
rect 16439 20352 16488 20380
rect 16439 20349 16451 20352
rect 16393 20343 16451 20349
rect 16482 20340 16488 20352
rect 16540 20340 16546 20392
rect 16592 20389 16620 20476
rect 17236 20457 17264 20488
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 18414 20516 18420 20528
rect 17681 20479 17739 20485
rect 17926 20488 18420 20516
rect 17221 20451 17279 20457
rect 16776 20420 17080 20448
rect 16776 20389 16804 20420
rect 17052 20392 17080 20420
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 17696 20448 17724 20479
rect 17543 20420 17724 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 16577 20383 16635 20389
rect 16577 20349 16589 20383
rect 16623 20349 16635 20383
rect 16577 20343 16635 20349
rect 16761 20383 16819 20389
rect 16761 20349 16773 20383
rect 16807 20349 16819 20383
rect 16761 20343 16819 20349
rect 16942 20340 16948 20392
rect 17000 20340 17006 20392
rect 17034 20340 17040 20392
rect 17092 20340 17098 20392
rect 17310 20340 17316 20392
rect 17368 20340 17374 20392
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20380 17463 20383
rect 17586 20380 17592 20392
rect 17451 20352 17592 20380
rect 17451 20349 17463 20352
rect 17405 20343 17463 20349
rect 17586 20340 17592 20352
rect 17644 20380 17650 20392
rect 17926 20380 17954 20488
rect 18414 20476 18420 20488
rect 18472 20476 18478 20528
rect 18598 20476 18604 20528
rect 18656 20516 18662 20528
rect 19794 20516 19800 20528
rect 18656 20488 19800 20516
rect 18656 20476 18662 20488
rect 19794 20476 19800 20488
rect 19852 20476 19858 20528
rect 20254 20476 20260 20528
rect 20312 20476 20318 20528
rect 20349 20519 20407 20525
rect 20349 20485 20361 20519
rect 20395 20516 20407 20519
rect 20640 20516 20668 20556
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 21910 20584 21916 20596
rect 20772 20556 21916 20584
rect 20772 20544 20778 20556
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22554 20544 22560 20596
rect 22612 20544 22618 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 23290 20584 23296 20596
rect 22695 20556 23296 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23566 20584 23572 20596
rect 23492 20556 23572 20584
rect 22572 20516 22600 20544
rect 23492 20516 23520 20556
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 24670 20544 24676 20596
rect 24728 20544 24734 20596
rect 24765 20587 24823 20593
rect 24765 20553 24777 20587
rect 24811 20584 24823 20587
rect 25130 20584 25136 20596
rect 24811 20556 25136 20584
rect 24811 20553 24823 20556
rect 24765 20547 24823 20553
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 26206 20556 29040 20584
rect 25498 20516 25504 20528
rect 20395 20488 20576 20516
rect 20640 20488 21680 20516
rect 22572 20488 23520 20516
rect 23584 20488 25504 20516
rect 20395 20485 20407 20488
rect 20349 20479 20407 20485
rect 18506 20408 18512 20460
rect 18564 20448 18570 20460
rect 19150 20448 19156 20460
rect 18564 20420 19156 20448
rect 18564 20408 18570 20420
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 20272 20448 20300 20476
rect 20180 20420 20300 20448
rect 20548 20448 20576 20488
rect 20548 20420 21312 20448
rect 19702 20380 19708 20392
rect 17644 20352 17954 20380
rect 18064 20352 19708 20380
rect 17644 20340 17650 20352
rect 15378 20312 15384 20324
rect 13679 20284 14504 20312
rect 14568 20284 15384 20312
rect 13679 20281 13691 20284
rect 13633 20275 13691 20281
rect 9447 20216 9996 20244
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 10134 20204 10140 20256
rect 10192 20204 10198 20256
rect 10594 20204 10600 20256
rect 10652 20244 10658 20256
rect 11606 20244 11612 20256
rect 10652 20216 11612 20244
rect 10652 20204 10658 20216
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 14568 20253 14596 20284
rect 15378 20272 15384 20284
rect 15436 20272 15442 20324
rect 17862 20321 17868 20324
rect 17849 20315 17868 20321
rect 16040 20284 17540 20312
rect 14553 20247 14611 20253
rect 14553 20213 14565 20247
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14691 20216 14841 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 14829 20207 14887 20213
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 16040 20253 16068 20284
rect 17512 20256 17540 20284
rect 17849 20281 17861 20315
rect 17849 20275 17868 20281
rect 17862 20272 17868 20275
rect 17920 20272 17926 20324
rect 18064 20321 18092 20352
rect 19702 20340 19708 20352
rect 19760 20340 19766 20392
rect 20180 20389 20208 20420
rect 21284 20392 21312 20420
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 20254 20340 20260 20392
rect 20312 20340 20318 20392
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20349 20499 20383
rect 20441 20343 20499 20349
rect 18049 20315 18107 20321
rect 18049 20281 18061 20315
rect 18095 20281 18107 20315
rect 20456 20312 20484 20343
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 20772 20352 21189 20380
rect 20772 20340 20778 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 21266 20340 21272 20392
rect 21324 20340 21330 20392
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21407 20352 21496 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 18049 20275 18107 20281
rect 18156 20284 20484 20312
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 14976 20216 16037 20244
rect 14976 20204 14982 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 16117 20247 16175 20253
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16485 20247 16543 20253
rect 16485 20244 16497 20247
rect 16163 20216 16497 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16485 20213 16497 20216
rect 16531 20244 16543 20247
rect 16574 20244 16580 20256
rect 16531 20216 16580 20244
rect 16531 20213 16543 20216
rect 16485 20207 16543 20213
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17037 20247 17095 20253
rect 17037 20244 17049 20247
rect 17000 20216 17049 20244
rect 17000 20204 17006 20216
rect 17037 20213 17049 20216
rect 17083 20213 17095 20247
rect 17037 20207 17095 20213
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 18156 20244 18184 20284
rect 20898 20272 20904 20324
rect 20956 20272 20962 20324
rect 21468 20256 21496 20352
rect 21542 20340 21548 20392
rect 21600 20340 21606 20392
rect 21652 20380 21680 20488
rect 23584 20460 23612 20488
rect 25498 20476 25504 20488
rect 25556 20516 25562 20528
rect 26206 20516 26234 20556
rect 25556 20488 26234 20516
rect 25556 20476 25562 20488
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 22244 20420 22569 20448
rect 22244 20408 22250 20420
rect 22557 20417 22569 20420
rect 22603 20417 22615 20451
rect 22557 20411 22615 20417
rect 23566 20408 23572 20460
rect 23624 20408 23630 20460
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 23716 20420 24440 20448
rect 23716 20408 23722 20420
rect 22465 20383 22523 20389
rect 21652 20352 22232 20380
rect 22204 20321 22232 20352
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 24302 20380 24308 20392
rect 22511 20352 24308 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 24302 20340 24308 20352
rect 24360 20340 24366 20392
rect 22189 20315 22247 20321
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 23382 20312 23388 20324
rect 22235 20284 23388 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 23750 20272 23756 20324
rect 23808 20272 23814 20324
rect 17552 20216 18184 20244
rect 17552 20204 17558 20216
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 19334 20244 19340 20256
rect 18380 20216 19340 20244
rect 18380 20204 18386 20216
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 20530 20244 20536 20256
rect 20312 20216 20536 20244
rect 20312 20204 20318 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 21450 20204 21456 20256
rect 21508 20204 21514 20256
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 22462 20244 22468 20256
rect 22327 20216 22468 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 22462 20204 22468 20216
rect 22520 20244 22526 20256
rect 22646 20244 22652 20256
rect 22520 20216 22652 20244
rect 22520 20204 22526 20216
rect 22646 20204 22652 20216
rect 22704 20244 22710 20256
rect 23768 20244 23796 20272
rect 22704 20216 23796 20244
rect 24412 20244 24440 20420
rect 24578 20408 24584 20460
rect 24636 20408 24642 20460
rect 24857 20451 24915 20457
rect 24857 20417 24869 20451
rect 24903 20448 24915 20451
rect 25590 20448 25596 20460
rect 24903 20420 25596 20448
rect 24903 20417 24915 20420
rect 24857 20411 24915 20417
rect 24596 20380 24624 20408
rect 24964 20392 24992 20420
rect 25590 20408 25596 20420
rect 25648 20408 25654 20460
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20448 27675 20451
rect 28442 20448 28448 20460
rect 27663 20420 28448 20448
rect 27663 20417 27675 20420
rect 27617 20411 27675 20417
rect 28442 20408 28448 20420
rect 28500 20408 28506 20460
rect 29012 20448 29040 20556
rect 29086 20544 29092 20596
rect 29144 20584 29150 20596
rect 29365 20587 29423 20593
rect 29365 20584 29377 20587
rect 29144 20556 29377 20584
rect 29144 20544 29150 20556
rect 29365 20553 29377 20556
rect 29411 20553 29423 20587
rect 29365 20547 29423 20553
rect 29454 20544 29460 20596
rect 29512 20544 29518 20596
rect 30466 20544 30472 20596
rect 30524 20584 30530 20596
rect 31113 20587 31171 20593
rect 31113 20584 31125 20587
rect 30524 20556 31125 20584
rect 30524 20544 30530 20556
rect 31113 20553 31125 20556
rect 31159 20553 31171 20587
rect 31113 20547 31171 20553
rect 30558 20476 30564 20528
rect 30616 20476 30622 20528
rect 29012 20420 29132 20448
rect 24596 20367 24625 20380
rect 24582 20361 24640 20367
rect 24582 20327 24594 20361
rect 24628 20327 24640 20361
rect 24946 20340 24952 20392
rect 25004 20340 25010 20392
rect 27062 20340 27068 20392
rect 27120 20380 27126 20392
rect 27155 20383 27213 20389
rect 27155 20380 27167 20383
rect 27120 20352 27167 20380
rect 27120 20340 27126 20352
rect 27155 20349 27167 20352
rect 27201 20349 27213 20383
rect 27155 20343 27213 20349
rect 27479 20383 27537 20389
rect 27479 20349 27491 20383
rect 27525 20349 27537 20383
rect 27479 20343 27537 20349
rect 24582 20321 24640 20327
rect 24854 20272 24860 20324
rect 24912 20312 24918 20324
rect 27494 20312 27522 20343
rect 28626 20340 28632 20392
rect 28684 20380 28690 20392
rect 29104 20380 29132 20420
rect 30190 20408 30196 20460
rect 30248 20448 30254 20460
rect 30834 20448 30840 20460
rect 30248 20420 30840 20448
rect 30248 20408 30254 20420
rect 30834 20408 30840 20420
rect 30892 20448 30898 20460
rect 30892 20420 31248 20448
rect 30892 20408 30898 20420
rect 29457 20383 29515 20389
rect 28684 20354 28764 20380
rect 28997 20357 29055 20363
rect 28997 20354 29009 20357
rect 28684 20352 29009 20354
rect 28684 20340 28690 20352
rect 28736 20326 29009 20352
rect 28997 20323 29009 20326
rect 29043 20323 29055 20357
rect 29104 20352 29408 20380
rect 28997 20317 29055 20323
rect 24912 20284 27522 20312
rect 24912 20272 24918 20284
rect 29178 20272 29184 20324
rect 29236 20321 29242 20324
rect 29236 20315 29265 20321
rect 29253 20281 29265 20315
rect 29380 20312 29408 20352
rect 29457 20349 29469 20383
rect 29503 20380 29515 20383
rect 29914 20380 29920 20392
rect 29503 20352 29920 20380
rect 29503 20349 29515 20352
rect 29457 20343 29515 20349
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 30561 20383 30619 20389
rect 30561 20380 30573 20383
rect 30300 20352 30573 20380
rect 30300 20324 30328 20352
rect 30561 20349 30573 20352
rect 30607 20349 30619 20383
rect 30561 20343 30619 20349
rect 30742 20340 30748 20392
rect 30800 20340 30806 20392
rect 31018 20340 31024 20392
rect 31076 20340 31082 20392
rect 31220 20389 31248 20420
rect 31205 20383 31263 20389
rect 31205 20349 31217 20383
rect 31251 20349 31263 20383
rect 31205 20343 31263 20349
rect 29546 20312 29552 20324
rect 29380 20284 29552 20312
rect 29236 20275 29265 20281
rect 29236 20272 29242 20275
rect 29546 20272 29552 20284
rect 29604 20312 29610 20324
rect 29733 20315 29791 20321
rect 29733 20312 29745 20315
rect 29604 20284 29745 20312
rect 29604 20272 29610 20284
rect 29733 20281 29745 20284
rect 29779 20281 29791 20315
rect 29733 20275 29791 20281
rect 30282 20272 30288 20324
rect 30340 20272 30346 20324
rect 25314 20244 25320 20256
rect 24412 20216 25320 20244
rect 22704 20204 22710 20216
rect 25314 20204 25320 20216
rect 25372 20204 25378 20256
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 26786 20244 26792 20256
rect 25740 20216 26792 20244
rect 25740 20204 25746 20216
rect 26786 20204 26792 20216
rect 26844 20204 26850 20256
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 28350 20204 28356 20256
rect 28408 20244 28414 20256
rect 29089 20247 29147 20253
rect 29089 20244 29101 20247
rect 28408 20216 29101 20244
rect 28408 20204 28414 20216
rect 29089 20213 29101 20216
rect 29135 20244 29147 20247
rect 29825 20247 29883 20253
rect 29825 20244 29837 20247
rect 29135 20216 29837 20244
rect 29135 20213 29147 20216
rect 29089 20207 29147 20213
rect 29825 20213 29837 20216
rect 29871 20244 29883 20247
rect 30098 20244 30104 20256
rect 29871 20216 30104 20244
rect 29871 20213 29883 20216
rect 29825 20207 29883 20213
rect 30098 20204 30104 20216
rect 30156 20204 30162 20256
rect 552 20154 31808 20176
rect 552 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 15946 20154
rect 15998 20102 16010 20154
rect 16062 20102 16074 20154
rect 16126 20102 16138 20154
rect 16190 20102 16202 20154
rect 16254 20102 23720 20154
rect 23772 20102 23784 20154
rect 23836 20102 23848 20154
rect 23900 20102 23912 20154
rect 23964 20102 23976 20154
rect 24028 20102 31494 20154
rect 31546 20102 31558 20154
rect 31610 20102 31622 20154
rect 31674 20102 31686 20154
rect 31738 20102 31750 20154
rect 31802 20102 31808 20154
rect 552 20080 31808 20102
rect 1118 20000 1124 20052
rect 1176 20000 1182 20052
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4028 20012 7512 20040
rect 4028 20000 4034 20012
rect 1136 19972 1164 20000
rect 1213 19975 1271 19981
rect 1213 19972 1225 19975
rect 1136 19944 1225 19972
rect 1213 19941 1225 19944
rect 1259 19941 1271 19975
rect 1213 19935 1271 19941
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19972 3019 19975
rect 3326 19972 3332 19984
rect 3007 19944 3332 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 3326 19932 3332 19944
rect 3384 19932 3390 19984
rect 4982 19932 4988 19984
rect 5040 19972 5046 19984
rect 5092 19972 5120 20012
rect 7484 19984 7512 20012
rect 9030 20000 9036 20052
rect 9088 20040 9094 20052
rect 9088 20012 9674 20040
rect 9088 20000 9094 20012
rect 5040 19944 5120 19972
rect 5040 19932 5046 19944
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 6181 19975 6239 19981
rect 6181 19972 6193 19975
rect 5684 19944 6193 19972
rect 5684 19932 5690 19944
rect 6181 19941 6193 19944
rect 6227 19941 6239 19975
rect 6181 19935 6239 19941
rect 6914 19932 6920 19984
rect 6972 19932 6978 19984
rect 7466 19932 7472 19984
rect 7524 19932 7530 19984
rect 2222 19864 2228 19916
rect 2280 19904 2286 19916
rect 2682 19904 2688 19916
rect 2280 19876 2688 19904
rect 2280 19864 2286 19876
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 3660 19876 4108 19904
rect 3660 19864 3666 19876
rect 937 19839 995 19845
rect 937 19805 949 19839
rect 983 19805 995 19839
rect 937 19799 995 19805
rect 952 19712 980 19799
rect 3050 19796 3056 19848
rect 3108 19836 3114 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3108 19808 3985 19836
rect 3108 19796 3114 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 4080 19836 4108 19876
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5905 19907 5963 19913
rect 5905 19904 5917 19907
rect 5592 19876 5917 19904
rect 5592 19864 5598 19876
rect 5905 19873 5917 19876
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 8021 19907 8079 19913
rect 8021 19904 8033 19907
rect 7892 19876 8033 19904
rect 7892 19864 7898 19876
rect 8021 19873 8033 19876
rect 8067 19873 8079 19907
rect 8021 19867 8079 19873
rect 6178 19836 6184 19848
rect 4080 19808 6184 19836
rect 3973 19799 4031 19805
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 6638 19796 6644 19848
rect 6696 19836 6702 19848
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 6696 19808 7941 19836
rect 6696 19796 6702 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8938 19836 8944 19848
rect 8343 19808 8944 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 3602 19768 3608 19780
rect 2424 19740 3608 19768
rect 934 19660 940 19712
rect 992 19700 998 19712
rect 2424 19700 2452 19740
rect 3602 19728 3608 19740
rect 3660 19728 3666 19780
rect 9416 19768 9444 19890
rect 9646 19836 9674 20012
rect 10410 20000 10416 20052
rect 10468 20000 10474 20052
rect 12250 20040 12256 20052
rect 10520 20012 12256 20040
rect 10042 19864 10048 19916
rect 10100 19904 10106 19916
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 10100 19876 10241 19904
rect 10100 19864 10106 19876
rect 10229 19873 10241 19876
rect 10275 19904 10287 19907
rect 10520 19904 10548 20012
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 13170 20040 13176 20052
rect 12575 20012 13176 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 17678 20040 17684 20052
rect 16540 20012 17684 20040
rect 16540 20000 16546 20012
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 17957 20043 18015 20049
rect 17957 20009 17969 20043
rect 18003 20040 18015 20043
rect 18506 20040 18512 20052
rect 18003 20012 18512 20040
rect 18003 20009 18015 20012
rect 17957 20003 18015 20009
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 21634 20040 21640 20052
rect 18932 20012 21640 20040
rect 18932 20000 18938 20012
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 24946 20040 24952 20052
rect 23348 20012 24952 20040
rect 23348 20000 23354 20012
rect 24946 20000 24952 20012
rect 25004 20040 25010 20052
rect 25133 20043 25191 20049
rect 25133 20040 25145 20043
rect 25004 20012 25145 20040
rect 25004 20000 25010 20012
rect 25133 20009 25145 20012
rect 25179 20009 25191 20043
rect 25133 20003 25191 20009
rect 26786 20000 26792 20052
rect 26844 20040 26850 20052
rect 27065 20043 27123 20049
rect 26844 20012 27016 20040
rect 26844 20000 26850 20012
rect 10275 19876 10548 19904
rect 10612 19944 12480 19972
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 10612 19836 10640 19944
rect 10689 19907 10747 19913
rect 10689 19873 10701 19907
rect 10735 19904 10747 19907
rect 10962 19904 10968 19916
rect 10735 19876 10968 19904
rect 10735 19873 10747 19876
rect 10689 19867 10747 19873
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 11204 19876 11345 19904
rect 11204 19864 11210 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11606 19864 11612 19916
rect 11664 19904 11670 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 11664 19876 11897 19904
rect 11664 19864 11670 19876
rect 11885 19873 11897 19876
rect 11931 19904 11943 19907
rect 11974 19904 11980 19916
rect 11931 19876 11980 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12250 19864 12256 19916
rect 12308 19864 12314 19916
rect 12452 19913 12480 19944
rect 12802 19932 12808 19984
rect 12860 19972 12866 19984
rect 12986 19972 12992 19984
rect 12860 19944 12992 19972
rect 12860 19932 12866 19944
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 13078 19932 13084 19984
rect 13136 19972 13142 19984
rect 14826 19972 14832 19984
rect 13136 19944 14832 19972
rect 13136 19932 13142 19944
rect 14826 19932 14832 19944
rect 14884 19972 14890 19984
rect 17310 19972 17316 19984
rect 14884 19944 17316 19972
rect 14884 19932 14890 19944
rect 17310 19932 17316 19944
rect 17368 19972 17374 19984
rect 17368 19944 18092 19972
rect 17368 19932 17374 19944
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 17034 19904 17040 19916
rect 15620 19876 17040 19904
rect 15620 19864 15626 19876
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 17552 19876 17601 19904
rect 17552 19864 17558 19876
rect 17589 19873 17601 19876
rect 17635 19904 17647 19907
rect 17954 19904 17960 19916
rect 17635 19876 17960 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 18064 19904 18092 19944
rect 18414 19932 18420 19984
rect 18472 19972 18478 19984
rect 18472 19944 18828 19972
rect 18472 19932 18478 19944
rect 18800 19913 18828 19944
rect 19150 19932 19156 19984
rect 19208 19972 19214 19984
rect 21542 19972 21548 19984
rect 19208 19944 21548 19972
rect 19208 19932 19214 19944
rect 21542 19932 21548 19944
rect 21600 19932 21606 19984
rect 22278 19932 22284 19984
rect 22336 19972 22342 19984
rect 22925 19975 22983 19981
rect 22925 19972 22937 19975
rect 22336 19944 22937 19972
rect 22336 19932 22342 19944
rect 22925 19941 22937 19944
rect 22971 19941 22983 19975
rect 22925 19935 22983 19941
rect 23017 19975 23075 19981
rect 23017 19941 23029 19975
rect 23063 19972 23075 19975
rect 24121 19975 24179 19981
rect 24121 19972 24133 19975
rect 23063 19944 23177 19972
rect 23063 19941 23075 19944
rect 23017 19935 23075 19941
rect 18265 19907 18323 19913
rect 18265 19904 18277 19907
rect 18064 19876 18277 19904
rect 18265 19873 18277 19876
rect 18311 19873 18323 19907
rect 18601 19907 18659 19913
rect 18601 19904 18613 19907
rect 18265 19867 18323 19873
rect 18432 19876 18613 19904
rect 9646 19808 10640 19836
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11514 19796 11520 19848
rect 11572 19796 11578 19848
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12526 19836 12532 19848
rect 11848 19808 12532 19836
rect 11848 19796 11854 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 16482 19836 16488 19848
rect 12676 19808 16488 19836
rect 12676 19796 12682 19808
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 17862 19836 17868 19848
rect 17727 19808 17868 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18138 19836 18144 19848
rect 18095 19808 18144 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 9490 19768 9496 19780
rect 9416 19740 9496 19768
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 9769 19771 9827 19777
rect 9769 19737 9781 19771
rect 9815 19768 9827 19771
rect 9815 19740 10180 19768
rect 9815 19737 9827 19740
rect 9769 19731 9827 19737
rect 992 19672 2452 19700
rect 992 19660 998 19672
rect 2682 19660 2688 19712
rect 2740 19700 2746 19712
rect 3970 19700 3976 19712
rect 2740 19672 3976 19700
rect 2740 19660 2746 19672
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 5350 19660 5356 19712
rect 5408 19709 5414 19712
rect 5408 19703 5457 19709
rect 5408 19669 5411 19703
rect 5445 19669 5457 19703
rect 5408 19663 5457 19669
rect 5408 19660 5414 19663
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 6972 19672 10057 19700
rect 6972 19660 6978 19672
rect 10045 19669 10057 19672
rect 10091 19669 10103 19703
rect 10152 19700 10180 19740
rect 10226 19728 10232 19780
rect 10284 19768 10290 19780
rect 14550 19768 14556 19780
rect 10284 19740 14556 19768
rect 10284 19728 10290 19740
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 18432 19768 18460 19876
rect 18601 19873 18613 19876
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19873 18843 19907
rect 18785 19867 18843 19873
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18616 19836 18644 19867
rect 18874 19864 18880 19916
rect 18932 19864 18938 19916
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19904 19027 19907
rect 19334 19904 19340 19916
rect 19015 19876 19340 19904
rect 19015 19873 19027 19876
rect 18969 19867 19027 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19426 19864 19432 19916
rect 19484 19864 19490 19916
rect 19518 19864 19524 19916
rect 19576 19904 19582 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19576 19876 19625 19904
rect 19576 19864 19582 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 19935 19876 20024 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 19444 19836 19472 19864
rect 18616 19808 19472 19836
rect 19628 19836 19656 19867
rect 19996 19836 20024 19876
rect 20070 19864 20076 19916
rect 20128 19864 20134 19916
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 21174 19904 21180 19916
rect 20772 19876 21180 19904
rect 20772 19864 20778 19876
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21910 19904 21916 19916
rect 21508 19876 21916 19904
rect 21508 19864 21514 19876
rect 21910 19864 21916 19876
rect 21968 19904 21974 19916
rect 21968 19876 22324 19904
rect 21968 19864 21974 19876
rect 20898 19836 20904 19848
rect 19628 19808 19932 19836
rect 19996 19808 20904 19836
rect 18509 19799 18567 19805
rect 17552 19740 18460 19768
rect 18524 19768 18552 19799
rect 19705 19771 19763 19777
rect 19705 19768 19717 19771
rect 18524 19740 19717 19768
rect 17552 19728 17558 19740
rect 19705 19737 19717 19740
rect 19751 19737 19763 19771
rect 19705 19731 19763 19737
rect 19794 19728 19800 19780
rect 19852 19728 19858 19780
rect 19904 19768 19932 19808
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 22094 19836 22100 19848
rect 21008 19808 22100 19836
rect 21008 19768 21036 19808
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 22186 19796 22192 19848
rect 22244 19796 22250 19848
rect 22296 19845 22324 19876
rect 22370 19864 22376 19916
rect 22428 19864 22434 19916
rect 23149 19904 23177 19944
rect 23308 19944 24133 19972
rect 23308 19904 23336 19944
rect 24121 19941 24133 19944
rect 24167 19941 24179 19975
rect 24121 19935 24179 19941
rect 24394 19932 24400 19984
rect 24452 19972 24458 19984
rect 24489 19975 24547 19981
rect 24489 19972 24501 19975
rect 24452 19944 24501 19972
rect 24452 19932 24458 19944
rect 24489 19941 24501 19944
rect 24535 19972 24547 19975
rect 24670 19972 24676 19984
rect 24535 19944 24676 19972
rect 24535 19941 24547 19944
rect 24489 19935 24547 19941
rect 24670 19932 24676 19944
rect 24728 19932 24734 19984
rect 26694 19972 26700 19984
rect 25148 19944 25636 19972
rect 23149 19876 23336 19904
rect 23382 19864 23388 19916
rect 23440 19864 23446 19916
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 23661 19907 23719 19913
rect 23661 19904 23673 19907
rect 23532 19876 23673 19904
rect 23532 19864 23538 19876
rect 23661 19873 23673 19876
rect 23707 19873 23719 19907
rect 23661 19867 23719 19873
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 23934 19904 23940 19916
rect 23891 19876 23940 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 23934 19864 23940 19876
rect 23992 19864 23998 19916
rect 24302 19864 24308 19916
rect 24360 19864 24366 19916
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 22281 19839 22339 19845
rect 22281 19805 22293 19839
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19836 22615 19839
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22603 19808 22661 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 22649 19799 22707 19805
rect 19904 19740 21036 19768
rect 21450 19728 21456 19780
rect 21508 19768 21514 19780
rect 22204 19768 22232 19796
rect 21508 19740 22232 19768
rect 22296 19768 22324 19799
rect 23014 19796 23020 19848
rect 23072 19796 23078 19848
rect 23134 19839 23192 19845
rect 23134 19805 23146 19839
rect 23180 19805 23192 19839
rect 24596 19836 24624 19867
rect 24762 19864 24768 19916
rect 24820 19864 24826 19916
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19902 25007 19907
rect 25148 19904 25176 19944
rect 25608 19916 25636 19944
rect 26528 19944 26700 19972
rect 26528 19916 26556 19944
rect 26694 19932 26700 19944
rect 26752 19972 26758 19984
rect 26752 19944 26924 19972
rect 26752 19932 26758 19944
rect 25056 19902 25176 19904
rect 24995 19876 25176 19902
rect 25225 19907 25283 19913
rect 24995 19874 25084 19876
rect 24995 19873 25007 19874
rect 24949 19867 25007 19873
rect 25225 19873 25237 19907
rect 25271 19873 25283 19907
rect 25225 19867 25283 19873
rect 24857 19839 24915 19845
rect 24857 19836 24869 19839
rect 24596 19808 24869 19836
rect 23134 19799 23192 19805
rect 24857 19805 24869 19808
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 23032 19768 23060 19796
rect 22296 19740 23060 19768
rect 21508 19728 21514 19740
rect 10594 19700 10600 19712
rect 10152 19672 10600 19700
rect 10045 19663 10103 19669
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 10962 19660 10968 19712
rect 11020 19660 11026 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 14182 19700 14188 19712
rect 11112 19672 14188 19700
rect 11112 19660 11118 19672
rect 14182 19660 14188 19672
rect 14240 19700 14246 19712
rect 16390 19700 16396 19712
rect 14240 19672 16396 19700
rect 14240 19660 14246 19672
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 17460 19672 17601 19700
rect 17460 19660 17466 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 17862 19660 17868 19712
rect 17920 19700 17926 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17920 19672 18153 19700
rect 17920 19660 17926 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 19245 19703 19303 19709
rect 19245 19700 19257 19703
rect 18564 19672 19257 19700
rect 18564 19660 18570 19672
rect 19245 19669 19257 19672
rect 19291 19669 19303 19703
rect 19245 19663 19303 19669
rect 19337 19703 19395 19709
rect 19337 19669 19349 19703
rect 19383 19700 19395 19703
rect 20806 19700 20812 19712
rect 19383 19672 20812 19700
rect 19383 19669 19395 19672
rect 19337 19663 19395 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 20898 19660 20904 19712
rect 20956 19700 20962 19712
rect 23149 19700 23177 19799
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 25240 19836 25268 19867
rect 25314 19864 25320 19916
rect 25372 19864 25378 19916
rect 25590 19864 25596 19916
rect 25648 19864 25654 19916
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 26421 19907 26479 19913
rect 26421 19904 26433 19907
rect 26384 19876 26433 19904
rect 26384 19864 26390 19876
rect 26421 19873 26433 19876
rect 26467 19873 26479 19907
rect 26421 19867 26479 19873
rect 26510 19864 26516 19916
rect 26568 19864 26574 19916
rect 26602 19864 26608 19916
rect 26660 19864 26666 19916
rect 26896 19913 26924 19944
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19873 26939 19907
rect 26881 19867 26939 19873
rect 25188 19808 25268 19836
rect 25188 19796 25194 19808
rect 26786 19796 26792 19848
rect 26844 19796 26850 19848
rect 26988 19836 27016 20012
rect 27065 20009 27077 20043
rect 27111 20040 27123 20043
rect 27154 20040 27160 20052
rect 27111 20012 27160 20040
rect 27111 20009 27123 20012
rect 27065 20003 27123 20009
rect 27154 20000 27160 20012
rect 27212 20000 27218 20052
rect 29178 20000 29184 20052
rect 29236 20000 29242 20052
rect 29454 20000 29460 20052
rect 29512 20000 29518 20052
rect 30742 20040 30748 20052
rect 29564 20012 30748 20040
rect 29196 19972 29224 20000
rect 27908 19944 29224 19972
rect 27430 19864 27436 19916
rect 27488 19904 27494 19916
rect 27908 19913 27936 19944
rect 27893 19907 27951 19913
rect 27893 19904 27905 19907
rect 27488 19876 27905 19904
rect 27488 19864 27494 19876
rect 27893 19873 27905 19876
rect 27939 19873 27951 19907
rect 27893 19867 27951 19873
rect 28074 19864 28080 19916
rect 28132 19864 28138 19916
rect 28169 19907 28227 19913
rect 28169 19873 28181 19907
rect 28215 19904 28227 19907
rect 29472 19904 29500 20000
rect 28215 19876 29500 19904
rect 28215 19873 28227 19876
rect 28169 19867 28227 19873
rect 29564 19836 29592 20012
rect 30742 20000 30748 20012
rect 30800 20000 30806 20052
rect 29730 19932 29736 19984
rect 29788 19972 29794 19984
rect 30653 19975 30711 19981
rect 30653 19972 30665 19975
rect 29788 19944 30665 19972
rect 29788 19932 29794 19944
rect 30653 19941 30665 19944
rect 30699 19972 30711 19975
rect 31018 19972 31024 19984
rect 30699 19944 31024 19972
rect 30699 19941 30711 19944
rect 30653 19935 30711 19941
rect 31018 19932 31024 19944
rect 31076 19932 31082 19984
rect 30377 19907 30435 19913
rect 30377 19873 30389 19907
rect 30423 19873 30435 19907
rect 30377 19867 30435 19873
rect 26988 19808 29592 19836
rect 30392 19836 30420 19867
rect 30466 19864 30472 19916
rect 30524 19864 30530 19916
rect 30742 19864 30748 19916
rect 30800 19864 30806 19916
rect 30760 19836 30788 19864
rect 30392 19808 30788 19836
rect 23293 19771 23351 19777
rect 23293 19737 23305 19771
rect 23339 19768 23351 19771
rect 26697 19771 26755 19777
rect 26697 19768 26709 19771
rect 23339 19740 26709 19768
rect 23339 19737 23351 19740
rect 23293 19731 23351 19737
rect 26697 19737 26709 19740
rect 26743 19737 26755 19771
rect 26697 19731 26755 19737
rect 27985 19771 28043 19777
rect 27985 19737 27997 19771
rect 28031 19768 28043 19771
rect 28074 19768 28080 19780
rect 28031 19740 28080 19768
rect 28031 19737 28043 19740
rect 27985 19731 28043 19737
rect 28074 19728 28080 19740
rect 28132 19768 28138 19780
rect 28534 19768 28540 19780
rect 28132 19740 28540 19768
rect 28132 19728 28138 19740
rect 28534 19728 28540 19740
rect 28592 19728 28598 19780
rect 20956 19672 23177 19700
rect 20956 19660 20962 19672
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24029 19703 24087 19709
rect 24029 19700 24041 19703
rect 23808 19672 24041 19700
rect 23808 19660 23814 19672
rect 24029 19669 24041 19672
rect 24075 19669 24087 19703
rect 24029 19663 24087 19669
rect 26050 19660 26056 19712
rect 26108 19700 26114 19712
rect 27709 19703 27767 19709
rect 27709 19700 27721 19703
rect 26108 19672 27721 19700
rect 26108 19660 26114 19672
rect 27709 19669 27721 19672
rect 27755 19669 27767 19703
rect 27709 19663 27767 19669
rect 552 19610 31648 19632
rect 552 19558 4285 19610
rect 4337 19558 4349 19610
rect 4401 19558 4413 19610
rect 4465 19558 4477 19610
rect 4529 19558 4541 19610
rect 4593 19558 12059 19610
rect 12111 19558 12123 19610
rect 12175 19558 12187 19610
rect 12239 19558 12251 19610
rect 12303 19558 12315 19610
rect 12367 19558 19833 19610
rect 19885 19558 19897 19610
rect 19949 19558 19961 19610
rect 20013 19558 20025 19610
rect 20077 19558 20089 19610
rect 20141 19558 27607 19610
rect 27659 19558 27671 19610
rect 27723 19558 27735 19610
rect 27787 19558 27799 19610
rect 27851 19558 27863 19610
rect 27915 19558 31648 19610
rect 552 19536 31648 19558
rect 934 19456 940 19508
rect 992 19456 998 19508
rect 3050 19456 3056 19508
rect 3108 19456 3114 19508
rect 3421 19499 3479 19505
rect 3421 19465 3433 19499
rect 3467 19465 3479 19499
rect 3421 19459 3479 19465
rect 6012 19468 8616 19496
rect 845 19363 903 19369
rect 845 19329 857 19363
rect 891 19360 903 19363
rect 952 19360 980 19456
rect 891 19332 980 19360
rect 3436 19360 3464 19459
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 3436 19332 4169 19360
rect 891 19329 903 19332
rect 845 19323 903 19329
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 2682 19292 2688 19304
rect 2254 19264 2688 19292
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 4172 19292 4200 19323
rect 4338 19320 4344 19372
rect 4396 19320 4402 19372
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4672 19332 4721 19360
rect 4672 19320 4678 19332
rect 4709 19329 4721 19332
rect 4755 19360 4767 19363
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 4755 19332 5549 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5537 19329 5549 19332
rect 5583 19360 5595 19363
rect 6012 19360 6040 19468
rect 6089 19431 6147 19437
rect 6089 19397 6101 19431
rect 6135 19397 6147 19431
rect 6089 19391 6147 19397
rect 5583 19332 6040 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 5350 19292 5356 19304
rect 2915 19264 3648 19292
rect 4172 19264 5356 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 1118 19184 1124 19236
rect 1176 19184 1182 19236
rect 3234 19184 3240 19236
rect 3292 19184 3298 19236
rect 3620 19224 3648 19264
rect 5350 19252 5356 19264
rect 5408 19292 5414 19304
rect 5994 19292 6000 19304
rect 5408 19264 6000 19292
rect 5408 19252 5414 19264
rect 5994 19252 6000 19264
rect 6052 19252 6058 19304
rect 6104 19292 6132 19391
rect 7926 19388 7932 19440
rect 7984 19388 7990 19440
rect 8588 19428 8616 19468
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 10042 19496 10048 19508
rect 9088 19468 10048 19496
rect 9088 19456 9094 19468
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10137 19499 10195 19505
rect 10137 19465 10149 19499
rect 10183 19496 10195 19499
rect 10226 19496 10232 19508
rect 10183 19468 10232 19496
rect 10183 19465 10195 19468
rect 10137 19459 10195 19465
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 10686 19456 10692 19508
rect 10744 19456 10750 19508
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 12802 19496 12808 19508
rect 11480 19468 12808 19496
rect 11480 19456 11486 19468
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13630 19496 13636 19508
rect 13096 19468 13636 19496
rect 9585 19431 9643 19437
rect 8588 19400 8800 19428
rect 6270 19320 6276 19372
rect 6328 19360 6334 19372
rect 8588 19369 8616 19400
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6328 19332 6837 19360
rect 6328 19320 6334 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19329 8631 19363
rect 8772 19360 8800 19400
rect 9585 19397 9597 19431
rect 9631 19428 9643 19431
rect 13096 19428 13124 19468
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19465 14335 19499
rect 14277 19459 14335 19465
rect 9631 19400 13124 19428
rect 13173 19431 13231 19437
rect 9631 19397 9643 19400
rect 9585 19391 9643 19397
rect 13173 19397 13185 19431
rect 13219 19428 13231 19431
rect 14292 19428 14320 19459
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 14553 19499 14611 19505
rect 14553 19496 14565 19499
rect 14424 19468 14565 19496
rect 14424 19456 14430 19468
rect 14553 19465 14565 19468
rect 14599 19465 14611 19499
rect 14553 19459 14611 19465
rect 14645 19499 14703 19505
rect 14645 19465 14657 19499
rect 14691 19496 14703 19499
rect 14734 19496 14740 19508
rect 14691 19468 14740 19496
rect 14691 19465 14703 19468
rect 14645 19459 14703 19465
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 15286 19456 15292 19508
rect 15344 19456 15350 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 16209 19499 16267 19505
rect 16209 19496 16221 19499
rect 15436 19468 16221 19496
rect 15436 19456 15442 19468
rect 16209 19465 16221 19468
rect 16255 19465 16267 19499
rect 16209 19459 16267 19465
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 16540 19468 17908 19496
rect 16540 19456 16546 19468
rect 14458 19428 14464 19440
rect 13219 19400 14464 19428
rect 13219 19397 13231 19400
rect 13173 19391 13231 19397
rect 9950 19360 9956 19372
rect 8772 19332 9956 19360
rect 8573 19323 8631 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 12618 19360 12624 19372
rect 11808 19332 12624 19360
rect 7374 19292 7380 19304
rect 6104 19264 7380 19292
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 8018 19252 8024 19304
rect 8076 19292 8082 19304
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 8076 19264 8125 19292
rect 8076 19252 8082 19264
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8113 19255 8171 19261
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19292 8815 19295
rect 10594 19292 10600 19304
rect 8803 19264 10600 19292
rect 8803 19261 8815 19264
rect 8757 19255 8815 19261
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 10962 19292 10968 19304
rect 10827 19264 10968 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11422 19252 11428 19304
rect 11480 19252 11486 19304
rect 11517 19295 11575 19301
rect 11517 19261 11529 19295
rect 11563 19292 11575 19295
rect 11808 19292 11836 19332
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13188 19360 13216 19391
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 17494 19428 17500 19440
rect 14752 19400 17500 19428
rect 14752 19360 14780 19400
rect 17494 19388 17500 19400
rect 17552 19388 17558 19440
rect 17880 19428 17908 19468
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18932 19468 18981 19496
rect 18932 19456 18938 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 19153 19499 19211 19505
rect 19153 19496 19165 19499
rect 19116 19468 19165 19496
rect 19116 19456 19122 19468
rect 19153 19465 19165 19468
rect 19199 19465 19211 19499
rect 19153 19459 19211 19465
rect 19337 19499 19395 19505
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 20898 19496 20904 19508
rect 19383 19468 20904 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 22278 19496 22284 19508
rect 21928 19468 22284 19496
rect 18598 19428 18604 19440
rect 17880 19400 18604 19428
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 19484 19400 19564 19428
rect 19484 19388 19490 19400
rect 12728 19332 13216 19360
rect 14292 19332 14780 19360
rect 14829 19363 14887 19369
rect 11563 19264 11836 19292
rect 11563 19261 11575 19264
rect 11517 19255 11575 19261
rect 11882 19252 11888 19304
rect 11940 19252 11946 19304
rect 12728 19301 12756 19332
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 12691 19264 12725 19292
rect 12437 19255 12495 19261
rect 12713 19261 12725 19264
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 3620 19196 3740 19224
rect 2590 19116 2596 19168
rect 2648 19116 2654 19168
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3437 19159 3495 19165
rect 3437 19156 3449 19159
rect 3384 19128 3449 19156
rect 3384 19116 3390 19128
rect 3437 19125 3449 19128
rect 3483 19125 3495 19159
rect 3437 19119 3495 19125
rect 3602 19116 3608 19168
rect 3660 19116 3666 19168
rect 3712 19165 3740 19196
rect 4908 19196 5396 19224
rect 4908 19168 4936 19196
rect 5368 19168 5396 19196
rect 5442 19184 5448 19236
rect 5500 19224 5506 19236
rect 5500 19196 6316 19224
rect 5500 19184 5506 19196
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19125 3755 19159
rect 3697 19119 3755 19125
rect 4062 19116 4068 19168
rect 4120 19116 4126 19168
rect 4798 19116 4804 19168
rect 4856 19116 4862 19168
rect 4890 19116 4896 19168
rect 4948 19116 4954 19168
rect 5258 19116 5264 19168
rect 5316 19116 5322 19168
rect 5350 19116 5356 19168
rect 5408 19116 5414 19168
rect 5626 19116 5632 19168
rect 5684 19116 5690 19168
rect 5721 19159 5779 19165
rect 5721 19125 5733 19159
rect 5767 19156 5779 19159
rect 5994 19156 6000 19168
rect 5767 19128 6000 19156
rect 5767 19125 5779 19128
rect 5721 19119 5779 19125
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 6288 19165 6316 19196
rect 6638 19184 6644 19236
rect 6696 19184 6702 19236
rect 7561 19227 7619 19233
rect 7561 19193 7573 19227
rect 7607 19224 7619 19227
rect 7926 19224 7932 19236
rect 7607 19196 7932 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 7926 19184 7932 19196
rect 7984 19224 7990 19236
rect 9030 19224 9036 19236
rect 7984 19196 9036 19224
rect 7984 19184 7990 19196
rect 9030 19184 9036 19196
rect 9088 19184 9094 19236
rect 9309 19227 9367 19233
rect 9309 19224 9321 19227
rect 9140 19196 9321 19224
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19125 6331 19159
rect 6273 19119 6331 19125
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 6733 19159 6791 19165
rect 6733 19156 6745 19159
rect 6604 19128 6745 19156
rect 6604 19116 6610 19128
rect 6733 19125 6745 19128
rect 6779 19125 6791 19159
rect 6733 19119 6791 19125
rect 7466 19116 7472 19168
rect 7524 19116 7530 19168
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 9140 19165 9168 19196
rect 9309 19193 9321 19196
rect 9355 19193 9367 19227
rect 9309 19187 9367 19193
rect 9858 19184 9864 19236
rect 9916 19184 9922 19236
rect 11606 19184 11612 19236
rect 11664 19184 11670 19236
rect 11747 19227 11805 19233
rect 11747 19193 11759 19227
rect 11793 19224 11805 19227
rect 12253 19227 12311 19233
rect 12253 19224 12265 19227
rect 11793 19196 12265 19224
rect 11793 19193 11805 19196
rect 11747 19187 11805 19193
rect 12253 19193 12265 19196
rect 12299 19193 12311 19227
rect 12253 19187 12311 19193
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19125 9183 19159
rect 9125 19119 9183 19125
rect 11238 19116 11244 19168
rect 11296 19116 11302 19168
rect 12452 19156 12480 19255
rect 12986 19252 12992 19304
rect 13044 19252 13050 19304
rect 13173 19295 13231 19301
rect 13173 19261 13185 19295
rect 13219 19292 13231 19295
rect 13630 19292 13636 19304
rect 13219 19264 13636 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13906 19252 13912 19304
rect 13964 19252 13970 19304
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 14292 19292 14320 19332
rect 14829 19329 14841 19363
rect 14875 19360 14887 19363
rect 16390 19360 16396 19372
rect 14875 19332 16396 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 18414 19360 18420 19372
rect 17184 19332 18420 19360
rect 17184 19320 17190 19332
rect 14047 19264 14320 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14366 19252 14372 19304
rect 14424 19252 14430 19304
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14700 19264 14933 19292
rect 14700 19252 14706 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15286 19292 15292 19304
rect 15151 19264 15292 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 12621 19227 12679 19233
rect 12621 19193 12633 19227
rect 12667 19224 12679 19227
rect 13722 19224 13728 19236
rect 12667 19196 13728 19224
rect 12667 19193 12679 19196
rect 12621 19187 12679 19193
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 13814 19156 13820 19168
rect 12452 19128 13820 19156
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14660 19156 14688 19252
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 15028 19224 15056 19255
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 15562 19252 15568 19304
rect 15620 19252 15626 19304
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19261 15807 19295
rect 15749 19255 15807 19261
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 14792 19196 15056 19224
rect 14792 19184 14798 19196
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 15672 19224 15700 19255
rect 15252 19196 15700 19224
rect 15764 19224 15792 19255
rect 16390 19224 16396 19236
rect 15764 19196 16396 19224
rect 15252 19184 15258 19196
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 16500 19156 16528 19255
rect 16574 19252 16580 19304
rect 16632 19252 16638 19304
rect 16669 19295 16727 19301
rect 16669 19261 16681 19295
rect 16715 19292 16727 19295
rect 16850 19292 16856 19304
rect 16715 19264 16856 19292
rect 16715 19261 16727 19264
rect 16669 19255 16727 19261
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 16942 19252 16948 19304
rect 17000 19252 17006 19304
rect 17037 19295 17095 19301
rect 17037 19261 17049 19295
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 16574 19156 16580 19168
rect 14660 19128 16580 19156
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 17052 19156 17080 19255
rect 17218 19252 17224 19304
rect 17276 19252 17282 19304
rect 17328 19301 17356 19332
rect 18414 19320 18420 19332
rect 18472 19360 18478 19372
rect 19536 19360 19564 19400
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 21928 19428 21956 19468
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 24397 19499 24455 19505
rect 24397 19496 24409 19499
rect 23440 19468 24409 19496
rect 23440 19456 23446 19468
rect 24397 19465 24409 19468
rect 24443 19465 24455 19499
rect 24397 19459 24455 19465
rect 24854 19456 24860 19508
rect 24912 19456 24918 19508
rect 26145 19499 26203 19505
rect 26145 19465 26157 19499
rect 26191 19465 26203 19499
rect 26145 19459 26203 19465
rect 19668 19400 21956 19428
rect 19668 19388 19674 19400
rect 20714 19360 20720 19372
rect 18472 19332 19472 19360
rect 19536 19332 20208 19360
rect 18472 19320 18478 19332
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19292 17463 19295
rect 17494 19292 17500 19304
rect 17451 19264 17500 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 18966 19292 18972 19304
rect 17736 19264 18972 19292
rect 17736 19252 17742 19264
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19444 19301 19472 19332
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 19116 19264 19257 19292
rect 19116 19252 19122 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19292 19487 19295
rect 19475 19264 19748 19292
rect 19475 19261 19487 19264
rect 19429 19255 19487 19261
rect 19720 19236 19748 19264
rect 17770 19224 17776 19236
rect 17512 19196 17776 19224
rect 17512 19156 17540 19196
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 18598 19184 18604 19236
rect 18656 19224 18662 19236
rect 18785 19227 18843 19233
rect 18785 19224 18797 19227
rect 18656 19196 18797 19224
rect 18656 19184 18662 19196
rect 18785 19193 18797 19196
rect 18831 19193 18843 19227
rect 18785 19187 18843 19193
rect 18892 19196 19657 19224
rect 17052 19128 17540 19156
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 17678 19156 17684 19168
rect 17635 19128 17684 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 18892 19156 18920 19196
rect 17920 19128 18920 19156
rect 18995 19159 19053 19165
rect 17920 19116 17926 19128
rect 18995 19125 19007 19159
rect 19041 19156 19053 19159
rect 19426 19156 19432 19168
rect 19041 19128 19432 19156
rect 19041 19125 19053 19128
rect 18995 19119 19053 19125
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 19629 19156 19657 19196
rect 19702 19184 19708 19236
rect 19760 19184 19766 19236
rect 20180 19168 20208 19332
rect 20272 19332 20720 19360
rect 20272 19301 20300 19332
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 20257 19295 20315 19301
rect 20257 19261 20269 19295
rect 20303 19261 20315 19295
rect 20257 19255 20315 19261
rect 20346 19252 20352 19304
rect 20404 19252 20410 19304
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 20622 19292 20628 19304
rect 20579 19264 20628 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20718 19273 20776 19279
rect 20718 19239 20730 19273
rect 20764 19239 20776 19273
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 20990 19252 20996 19304
rect 21048 19252 21054 19304
rect 21177 19295 21235 19301
rect 21177 19261 21189 19295
rect 21223 19292 21235 19295
rect 21468 19292 21496 19323
rect 21634 19320 21640 19372
rect 21692 19320 21698 19372
rect 21928 19369 21956 19400
rect 22094 19388 22100 19440
rect 22152 19428 22158 19440
rect 24762 19428 24768 19440
rect 22152 19400 24768 19428
rect 22152 19388 22158 19400
rect 24762 19388 24768 19400
rect 24820 19428 24826 19440
rect 25130 19428 25136 19440
rect 24820 19400 25136 19428
rect 24820 19388 24826 19400
rect 25130 19388 25136 19400
rect 25188 19388 25194 19440
rect 26160 19428 26188 19459
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 26697 19499 26755 19505
rect 26697 19496 26709 19499
rect 26660 19468 26709 19496
rect 26660 19456 26666 19468
rect 26697 19465 26709 19468
rect 26743 19465 26755 19499
rect 26697 19459 26755 19465
rect 29454 19456 29460 19508
rect 29512 19456 29518 19508
rect 29914 19456 29920 19508
rect 29972 19456 29978 19508
rect 30837 19499 30895 19505
rect 30837 19465 30849 19499
rect 30883 19465 30895 19499
rect 30837 19459 30895 19465
rect 27430 19428 27436 19440
rect 26160 19400 27436 19428
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19329 21971 19363
rect 21913 19323 21971 19329
rect 22186 19320 22192 19372
rect 22244 19360 22250 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 22244 19332 22293 19360
rect 22244 19320 22250 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22281 19323 22339 19329
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19360 22431 19363
rect 22646 19360 22652 19372
rect 22419 19332 22652 19360
rect 22419 19329 22431 19332
rect 22373 19323 22431 19329
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 23106 19320 23112 19372
rect 23164 19320 23170 19372
rect 23934 19320 23940 19372
rect 23992 19360 23998 19372
rect 24210 19360 24216 19372
rect 23992 19332 24216 19360
rect 23992 19320 23998 19332
rect 24210 19320 24216 19332
rect 24268 19360 24274 19372
rect 26160 19360 26188 19400
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 28997 19431 29055 19437
rect 28997 19397 29009 19431
rect 29043 19428 29055 19431
rect 29086 19428 29092 19440
rect 29043 19400 29092 19428
rect 29043 19397 29055 19400
rect 28997 19391 29055 19397
rect 29086 19388 29092 19400
rect 29144 19388 29150 19440
rect 29472 19428 29500 19456
rect 30282 19428 30288 19440
rect 29472 19400 30288 19428
rect 30282 19388 30288 19400
rect 30340 19428 30346 19440
rect 30852 19428 30880 19459
rect 30340 19400 30880 19428
rect 30340 19388 30346 19400
rect 24268 19332 26188 19360
rect 24268 19320 24274 19332
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 27396 19332 30604 19360
rect 27396 19320 27402 19332
rect 21223 19264 21496 19292
rect 21223 19261 21235 19264
rect 21177 19255 21235 19261
rect 20718 19236 20776 19239
rect 20714 19184 20720 19236
rect 20772 19184 20778 19236
rect 21085 19227 21143 19233
rect 21085 19193 21097 19227
rect 21131 19224 21143 19227
rect 21652 19224 21680 19320
rect 21726 19252 21732 19304
rect 21784 19252 21790 19304
rect 21818 19252 21824 19304
rect 21876 19292 21882 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 21876 19264 22477 19292
rect 21876 19252 21882 19264
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22186 19224 22192 19236
rect 21131 19196 21588 19224
rect 21652 19196 22192 19224
rect 21131 19193 21143 19196
rect 21085 19187 21143 19193
rect 19794 19156 19800 19168
rect 19629 19128 19800 19156
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 20162 19116 20168 19168
rect 20220 19116 20226 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 21361 19159 21419 19165
rect 21361 19156 21373 19159
rect 20404 19128 21373 19156
rect 20404 19116 20410 19128
rect 21361 19125 21373 19128
rect 21407 19125 21419 19159
rect 21560 19156 21588 19196
rect 22186 19184 22192 19196
rect 22244 19184 22250 19236
rect 22480 19224 22508 19255
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 23017 19295 23075 19301
rect 23017 19261 23029 19295
rect 23063 19292 23075 19295
rect 23198 19292 23204 19304
rect 23063 19264 23204 19292
rect 23063 19261 23075 19264
rect 23017 19255 23075 19261
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19292 23535 19295
rect 23658 19292 23664 19304
rect 23523 19264 23664 19292
rect 23523 19261 23535 19264
rect 23477 19255 23535 19261
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 23842 19252 23848 19304
rect 23900 19252 23906 19304
rect 24029 19295 24087 19301
rect 24029 19261 24041 19295
rect 24075 19261 24087 19295
rect 24029 19255 24087 19261
rect 24581 19295 24639 19301
rect 24581 19261 24593 19295
rect 24627 19261 24639 19295
rect 24581 19255 24639 19261
rect 22646 19224 22652 19236
rect 22480 19196 22652 19224
rect 22646 19184 22652 19196
rect 22704 19184 22710 19236
rect 22756 19196 22968 19224
rect 22097 19159 22155 19165
rect 22097 19156 22109 19159
rect 21560 19128 22109 19156
rect 21361 19119 21419 19125
rect 22097 19125 22109 19128
rect 22143 19125 22155 19159
rect 22097 19119 22155 19125
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 22756 19156 22784 19196
rect 22428 19128 22784 19156
rect 22428 19116 22434 19128
rect 22830 19116 22836 19168
rect 22888 19116 22894 19168
rect 22940 19156 22968 19196
rect 23106 19184 23112 19236
rect 23164 19224 23170 19236
rect 24044 19224 24072 19255
rect 23164 19196 24072 19224
rect 24596 19224 24624 19255
rect 24670 19252 24676 19304
rect 24728 19252 24734 19304
rect 24949 19295 25007 19301
rect 24949 19261 24961 19295
rect 24995 19292 25007 19295
rect 25866 19292 25872 19304
rect 24995 19264 25872 19292
rect 24995 19261 25007 19264
rect 24949 19255 25007 19261
rect 25866 19252 25872 19264
rect 25924 19252 25930 19304
rect 26050 19252 26056 19304
rect 26108 19252 26114 19304
rect 26329 19295 26387 19301
rect 26329 19261 26341 19295
rect 26375 19261 26387 19295
rect 26329 19255 26387 19261
rect 26068 19224 26096 19252
rect 24596 19196 26096 19224
rect 23164 19184 23170 19196
rect 26142 19184 26148 19236
rect 26200 19184 26206 19236
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 22940 19128 23213 19156
rect 23201 19125 23213 19128
rect 23247 19156 23259 19159
rect 23290 19156 23296 19168
rect 23247 19128 23296 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 23385 19159 23443 19165
rect 23385 19125 23397 19159
rect 23431 19156 23443 19159
rect 23845 19159 23903 19165
rect 23845 19156 23857 19159
rect 23431 19128 23857 19156
rect 23431 19125 23443 19128
rect 23385 19119 23443 19125
rect 23845 19125 23857 19128
rect 23891 19125 23903 19159
rect 23845 19119 23903 19125
rect 24118 19116 24124 19168
rect 24176 19156 24182 19168
rect 26344 19156 26372 19255
rect 26418 19252 26424 19304
rect 26476 19252 26482 19304
rect 26878 19252 26884 19304
rect 26936 19252 26942 19304
rect 27154 19252 27160 19304
rect 27212 19252 27218 19304
rect 28994 19252 29000 19304
rect 29052 19252 29058 19304
rect 29178 19252 29184 19304
rect 29236 19252 29242 19304
rect 29270 19252 29276 19304
rect 29328 19252 29334 19304
rect 29362 19252 29368 19304
rect 29420 19252 29426 19304
rect 29457 19295 29515 19301
rect 29457 19261 29469 19295
rect 29503 19261 29515 19295
rect 29457 19255 29515 19261
rect 27065 19227 27123 19233
rect 27065 19224 27077 19227
rect 26620 19196 27077 19224
rect 26620 19165 26648 19196
rect 27065 19193 27077 19196
rect 27111 19193 27123 19227
rect 29012 19224 29040 19252
rect 29472 19224 29500 19255
rect 29638 19252 29644 19304
rect 29696 19252 29702 19304
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 30101 19295 30159 19301
rect 30101 19292 30113 19295
rect 29880 19264 30113 19292
rect 29880 19252 29886 19264
rect 30101 19261 30113 19264
rect 30147 19261 30159 19295
rect 30101 19255 30159 19261
rect 30190 19252 30196 19304
rect 30248 19292 30254 19304
rect 30370 19295 30428 19301
rect 30370 19292 30382 19295
rect 30248 19264 30382 19292
rect 30248 19252 30254 19264
rect 30370 19261 30382 19264
rect 30416 19261 30428 19295
rect 30370 19255 30428 19261
rect 30478 19295 30536 19301
rect 30478 19261 30490 19295
rect 30524 19261 30536 19295
rect 30478 19255 30536 19261
rect 29012 19196 29500 19224
rect 27065 19187 27123 19193
rect 24176 19128 26372 19156
rect 26605 19159 26663 19165
rect 24176 19116 24182 19128
rect 26605 19125 26617 19159
rect 26651 19125 26663 19159
rect 26605 19119 26663 19125
rect 26694 19116 26700 19168
rect 26752 19156 26758 19168
rect 30484 19156 30512 19255
rect 30576 19224 30604 19332
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 31018 19360 31024 19372
rect 30892 19332 31024 19360
rect 30892 19320 30898 19332
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 30650 19252 30656 19304
rect 30708 19292 30714 19304
rect 30708 19264 31064 19292
rect 30708 19252 30714 19264
rect 31036 19233 31064 19264
rect 30805 19227 30863 19233
rect 30805 19224 30817 19227
rect 30576 19196 30817 19224
rect 30805 19193 30817 19196
rect 30851 19193 30863 19227
rect 30805 19187 30863 19193
rect 31021 19227 31079 19233
rect 31021 19193 31033 19227
rect 31067 19193 31079 19227
rect 31021 19187 31079 19193
rect 26752 19128 30512 19156
rect 26752 19116 26758 19128
rect 30650 19116 30656 19168
rect 30708 19116 30714 19168
rect 552 19066 31808 19088
rect 552 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 15946 19066
rect 15998 19014 16010 19066
rect 16062 19014 16074 19066
rect 16126 19014 16138 19066
rect 16190 19014 16202 19066
rect 16254 19014 23720 19066
rect 23772 19014 23784 19066
rect 23836 19014 23848 19066
rect 23900 19014 23912 19066
rect 23964 19014 23976 19066
rect 24028 19014 31494 19066
rect 31546 19014 31558 19066
rect 31610 19014 31622 19066
rect 31674 19014 31686 19066
rect 31738 19014 31750 19066
rect 31802 19014 31808 19066
rect 552 18992 31808 19014
rect 1118 18912 1124 18964
rect 1176 18952 1182 18964
rect 1213 18955 1271 18961
rect 1213 18952 1225 18955
rect 1176 18924 1225 18952
rect 1176 18912 1182 18924
rect 1213 18921 1225 18924
rect 1259 18921 1271 18955
rect 1213 18915 1271 18921
rect 1489 18955 1547 18961
rect 1489 18921 1501 18955
rect 1535 18921 1547 18955
rect 2038 18952 2044 18964
rect 1489 18915 1547 18921
rect 1596 18924 2044 18952
rect 1504 18884 1532 18915
rect 952 18856 1532 18884
rect 952 18825 980 18856
rect 937 18819 995 18825
rect 937 18785 949 18819
rect 983 18785 995 18819
rect 937 18779 995 18785
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1596 18816 1624 18924
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 2130 18912 2136 18964
rect 2188 18912 2194 18964
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 2832 18924 3157 18952
rect 2832 18912 2838 18924
rect 3145 18921 3157 18924
rect 3191 18921 3203 18955
rect 3145 18915 3203 18921
rect 3234 18912 3240 18964
rect 3292 18912 3298 18964
rect 3973 18955 4031 18961
rect 3973 18921 3985 18955
rect 4019 18952 4031 18955
rect 4062 18952 4068 18964
rect 4019 18924 4068 18952
rect 4019 18921 4031 18924
rect 3973 18915 4031 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4341 18955 4399 18961
rect 4341 18921 4353 18955
rect 4387 18952 4399 18955
rect 4706 18952 4712 18964
rect 4387 18924 4712 18952
rect 4387 18921 4399 18924
rect 4341 18915 4399 18921
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 4798 18912 4804 18964
rect 4856 18912 4862 18964
rect 5258 18912 5264 18964
rect 5316 18912 5322 18964
rect 6270 18912 6276 18964
rect 6328 18952 6334 18964
rect 8386 18952 8392 18964
rect 6328 18924 8392 18952
rect 6328 18912 6334 18924
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 8481 18955 8539 18961
rect 8481 18921 8493 18955
rect 8527 18952 8539 18955
rect 8662 18952 8668 18964
rect 8527 18924 8668 18952
rect 8527 18921 8539 18924
rect 8481 18915 8539 18921
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 9766 18952 9772 18964
rect 9048 18924 9772 18952
rect 1857 18887 1915 18893
rect 1857 18853 1869 18887
rect 1903 18884 1915 18887
rect 2148 18884 2176 18912
rect 1903 18856 2176 18884
rect 1903 18853 1915 18856
rect 1857 18847 1915 18853
rect 2590 18844 2596 18896
rect 2648 18884 2654 18896
rect 3252 18884 3280 18912
rect 2648 18856 3280 18884
rect 3605 18887 3663 18893
rect 2648 18844 2654 18856
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 3694 18884 3700 18896
rect 3651 18856 3700 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 3694 18844 3700 18856
rect 3752 18884 3758 18896
rect 5169 18887 5227 18893
rect 5169 18884 5181 18887
rect 3752 18856 5181 18884
rect 3752 18844 3758 18856
rect 5169 18853 5181 18856
rect 5215 18853 5227 18887
rect 5276 18884 5304 18912
rect 6181 18887 6239 18893
rect 6181 18884 6193 18887
rect 5276 18856 6193 18884
rect 5169 18847 5227 18853
rect 6181 18853 6193 18856
rect 6227 18853 6239 18887
rect 6181 18847 6239 18853
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 8941 18887 8999 18893
rect 8941 18884 8953 18887
rect 7892 18856 8953 18884
rect 7892 18844 7898 18856
rect 8941 18853 8953 18856
rect 8987 18853 8999 18887
rect 8941 18847 8999 18853
rect 1443 18788 1624 18816
rect 2685 18819 2743 18825
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2685 18785 2697 18819
rect 2731 18816 2743 18819
rect 3418 18816 3424 18828
rect 2731 18788 3424 18816
rect 2731 18785 2743 18788
rect 2685 18779 2743 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 3510 18776 3516 18828
rect 3568 18776 3574 18828
rect 4433 18819 4491 18825
rect 3620 18788 4292 18816
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 1121 18615 1179 18621
rect 1121 18581 1133 18615
rect 1167 18612 1179 18615
rect 1210 18612 1216 18624
rect 1167 18584 1216 18612
rect 1167 18581 1179 18584
rect 1121 18575 1179 18581
rect 1210 18572 1216 18584
rect 1268 18572 1274 18624
rect 1964 18612 1992 18711
rect 2148 18680 2176 18711
rect 2498 18708 2504 18760
rect 2556 18708 2562 18760
rect 2590 18708 2596 18760
rect 2648 18708 2654 18760
rect 2866 18680 2872 18692
rect 2148 18652 2872 18680
rect 2866 18640 2872 18652
rect 2924 18640 2930 18692
rect 3620 18680 3648 18788
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18748 3847 18751
rect 4062 18748 4068 18760
rect 3835 18720 4068 18748
rect 3835 18717 3847 18720
rect 3789 18711 3847 18717
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 2976 18652 3648 18680
rect 2976 18612 3004 18652
rect 1964 18584 3004 18612
rect 3050 18572 3056 18624
rect 3108 18572 3114 18624
rect 4080 18612 4108 18708
rect 4264 18692 4292 18788
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 5074 18816 5080 18828
rect 4479 18788 5080 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5736 18788 5825 18816
rect 5736 18760 5764 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4246 18640 4252 18692
rect 4304 18640 4310 18692
rect 4540 18612 4568 18711
rect 4706 18708 4712 18760
rect 4764 18748 4770 18760
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4764 18720 5273 18748
rect 4764 18708 4770 18720
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 5442 18708 5448 18760
rect 5500 18708 5506 18760
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 5813 18683 5871 18689
rect 5813 18680 5825 18683
rect 4856 18652 5825 18680
rect 4856 18640 4862 18652
rect 5813 18649 5825 18652
rect 5859 18649 5871 18683
rect 5813 18643 5871 18649
rect 4080 18584 4568 18612
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 6012 18612 6040 18779
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7024 18748 7052 18802
rect 8386 18776 8392 18828
rect 8444 18776 8450 18828
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 8849 18819 8907 18825
rect 8849 18816 8861 18819
rect 8720 18788 8861 18816
rect 8720 18776 8726 18788
rect 8849 18785 8861 18788
rect 8895 18816 8907 18819
rect 9048 18816 9076 18924
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 10045 18955 10103 18961
rect 10045 18952 10057 18955
rect 9916 18924 10057 18952
rect 9916 18912 9922 18924
rect 10045 18921 10057 18924
rect 10091 18921 10103 18955
rect 10045 18915 10103 18921
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 11296 18924 11560 18952
rect 11296 18912 11302 18924
rect 9585 18887 9643 18893
rect 9585 18853 9597 18887
rect 9631 18884 9643 18887
rect 10134 18884 10140 18896
rect 9631 18856 10140 18884
rect 9631 18853 9643 18856
rect 9585 18847 9643 18853
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 11532 18893 11560 18924
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 17126 18952 17132 18964
rect 12584 18924 17132 18952
rect 12584 18912 12590 18924
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17218 18912 17224 18964
rect 17276 18952 17282 18964
rect 17589 18955 17647 18961
rect 17589 18952 17601 18955
rect 17276 18924 17601 18952
rect 17276 18912 17282 18924
rect 17589 18921 17601 18924
rect 17635 18921 17647 18955
rect 17589 18915 17647 18921
rect 17678 18912 17684 18964
rect 17736 18912 17742 18964
rect 17770 18912 17776 18964
rect 17828 18912 17834 18964
rect 18322 18952 18328 18964
rect 17880 18924 18328 18952
rect 11517 18887 11575 18893
rect 11517 18853 11529 18887
rect 11563 18853 11575 18887
rect 11517 18847 11575 18853
rect 12986 18844 12992 18896
rect 13044 18884 13050 18896
rect 16666 18884 16672 18896
rect 13044 18856 16672 18884
rect 13044 18844 13050 18856
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 17696 18884 17724 18912
rect 17144 18856 17724 18884
rect 8895 18788 9076 18816
rect 9677 18819 9735 18825
rect 8895 18785 8907 18788
rect 8849 18779 8907 18785
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 10318 18816 10324 18828
rect 9723 18788 10324 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11241 18819 11299 18825
rect 11241 18816 11253 18819
rect 11112 18788 11253 18816
rect 11112 18776 11118 18788
rect 11241 18785 11253 18788
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 6972 18720 7052 18748
rect 8113 18751 8171 18757
rect 6972 18708 6978 18720
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8159 18720 8692 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8664 18680 8692 18720
rect 9030 18708 9036 18760
rect 9088 18708 9094 18760
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9950 18748 9956 18760
rect 9539 18720 9956 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 10686 18708 10692 18760
rect 10744 18708 10750 18760
rect 10962 18680 10968 18692
rect 8664 18652 10968 18680
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 11054 18640 11060 18692
rect 11112 18640 11118 18692
rect 11256 18680 11284 18779
rect 11606 18776 11612 18828
rect 11664 18776 11670 18828
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 11882 18816 11888 18828
rect 11839 18788 11888 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 11882 18776 11888 18788
rect 11940 18816 11946 18828
rect 13354 18816 13360 18828
rect 11940 18788 13360 18816
rect 11940 18776 11946 18788
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 13722 18776 13728 18828
rect 13780 18776 13786 18828
rect 13906 18776 13912 18828
rect 13964 18776 13970 18828
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 17144 18825 17172 18856
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18785 17187 18819
rect 17129 18779 17187 18785
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18816 17371 18819
rect 17880 18816 17908 18924
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 19518 18952 19524 18964
rect 18472 18924 19524 18952
rect 18472 18912 18478 18924
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 20898 18952 20904 18964
rect 20364 18924 20904 18952
rect 18138 18844 18144 18896
rect 18196 18884 18202 18896
rect 18196 18856 20024 18884
rect 18196 18844 18202 18856
rect 19996 18828 20024 18856
rect 17359 18788 17908 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 17954 18776 17960 18828
rect 18012 18776 18018 18828
rect 19058 18776 19064 18828
rect 19116 18776 19122 18828
rect 19150 18776 19156 18828
rect 19208 18776 19214 18828
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11471 18720 11713 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 13648 18748 13676 18776
rect 15562 18748 15568 18760
rect 13648 18720 15568 18748
rect 11701 18711 11759 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 18049 18751 18107 18757
rect 16632 18720 17816 18748
rect 16632 18708 16638 18720
rect 11256 18652 13768 18680
rect 5040 18584 6040 18612
rect 5040 18572 5046 18584
rect 6454 18572 6460 18624
rect 6512 18572 6518 18624
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18612 6699 18615
rect 7374 18612 7380 18624
rect 6687 18584 7380 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 7374 18572 7380 18584
rect 7432 18612 7438 18624
rect 8662 18612 8668 18624
rect 7432 18584 8668 18612
rect 7432 18572 7438 18584
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 10137 18615 10195 18621
rect 10137 18612 10149 18615
rect 9180 18584 10149 18612
rect 9180 18572 9186 18584
rect 10137 18581 10149 18584
rect 10183 18581 10195 18615
rect 10137 18575 10195 18581
rect 11517 18615 11575 18621
rect 11517 18581 11529 18615
rect 11563 18612 11575 18615
rect 11790 18612 11796 18624
rect 11563 18584 11796 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13078 18612 13084 18624
rect 12676 18584 13084 18612
rect 12676 18572 12682 18584
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 13740 18612 13768 18652
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 15194 18680 15200 18692
rect 14608 18652 15200 18680
rect 14608 18640 14614 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17678 18680 17684 18692
rect 16908 18652 17684 18680
rect 16908 18640 16914 18652
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 17788 18680 17816 18720
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18414 18748 18420 18760
rect 18279 18720 18420 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18064 18680 18092 18711
rect 17788 18652 18092 18680
rect 18156 18680 18184 18711
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 19168 18680 19196 18776
rect 19260 18748 19288 18779
rect 19334 18776 19340 18828
rect 19392 18776 19398 18828
rect 19426 18776 19432 18828
rect 19484 18776 19490 18828
rect 19794 18776 19800 18828
rect 19852 18776 19858 18828
rect 19978 18776 19984 18828
rect 20036 18776 20042 18828
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18816 20131 18819
rect 20364 18816 20392 18924
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21634 18952 21640 18964
rect 21048 18924 21640 18952
rect 21048 18912 21054 18924
rect 21634 18912 21640 18924
rect 21692 18952 21698 18964
rect 22370 18952 22376 18964
rect 21692 18924 22376 18952
rect 21692 18912 21698 18924
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 22465 18955 22523 18961
rect 22465 18921 22477 18955
rect 22511 18952 22523 18955
rect 22554 18952 22560 18964
rect 22511 18924 22560 18952
rect 22511 18921 22523 18924
rect 22465 18915 22523 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 22922 18912 22928 18964
rect 22980 18912 22986 18964
rect 23014 18912 23020 18964
rect 23072 18952 23078 18964
rect 23072 18924 23888 18952
rect 23072 18912 23078 18924
rect 21729 18887 21787 18893
rect 21729 18884 21741 18887
rect 20468 18856 21741 18884
rect 20468 18825 20496 18856
rect 21729 18853 21741 18856
rect 21775 18853 21787 18887
rect 23750 18884 23756 18896
rect 21729 18847 21787 18853
rect 21836 18856 23756 18884
rect 20119 18788 20392 18816
rect 20441 18819 20499 18825
rect 20119 18785 20131 18788
rect 20073 18779 20131 18785
rect 20441 18785 20453 18819
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 20530 18776 20536 18828
rect 20588 18776 20594 18828
rect 21174 18776 21180 18828
rect 21232 18776 21238 18828
rect 21450 18776 21456 18828
rect 21508 18816 21514 18828
rect 21836 18825 21864 18856
rect 23750 18844 23756 18856
rect 23808 18844 23814 18896
rect 23860 18884 23888 18924
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24728 18924 24777 18952
rect 24728 18912 24734 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 26878 18912 26884 18964
rect 26936 18912 26942 18964
rect 29270 18912 29276 18964
rect 29328 18952 29334 18964
rect 29365 18955 29423 18961
rect 29365 18952 29377 18955
rect 29328 18924 29377 18952
rect 29328 18912 29334 18924
rect 29365 18921 29377 18924
rect 29411 18921 29423 18955
rect 29365 18915 29423 18921
rect 30650 18912 30656 18964
rect 30708 18912 30714 18964
rect 26896 18884 26924 18912
rect 30668 18884 30696 18912
rect 23860 18856 26648 18884
rect 26896 18856 27016 18884
rect 26620 18828 26648 18856
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21508 18788 21649 18816
rect 21508 18776 21514 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18816 22155 18819
rect 22741 18819 22799 18825
rect 22741 18816 22753 18819
rect 22143 18788 22753 18816
rect 22143 18785 22155 18788
rect 22097 18779 22155 18785
rect 22741 18785 22753 18788
rect 22787 18785 22799 18819
rect 22741 18779 22799 18785
rect 19812 18748 19840 18776
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19260 18720 19472 18748
rect 19812 18720 20177 18748
rect 18156 18652 19196 18680
rect 14182 18612 14188 18624
rect 13740 18584 14188 18612
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 14826 18612 14832 18624
rect 14424 18584 14832 18612
rect 14424 18572 14430 18584
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 17770 18612 17776 18624
rect 15068 18584 17776 18612
rect 15068 18572 15074 18584
rect 17770 18572 17776 18584
rect 17828 18572 17834 18624
rect 18064 18612 18092 18652
rect 19334 18612 19340 18624
rect 18064 18584 19340 18612
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 19444 18612 19472 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20257 18751 20315 18757
rect 20257 18717 20269 18751
rect 20303 18748 20315 18751
rect 20303 18720 20496 18748
rect 20303 18717 20315 18720
rect 20257 18711 20315 18717
rect 19705 18683 19763 18689
rect 19705 18649 19717 18683
rect 19751 18680 19763 18683
rect 20468 18680 20496 18720
rect 20622 18708 20628 18760
rect 20680 18708 20686 18760
rect 21192 18748 21220 18776
rect 20916 18720 21220 18748
rect 20916 18689 20944 18720
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21600 18720 22017 18748
rect 21600 18708 21606 18720
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 20901 18683 20959 18689
rect 19751 18652 20392 18680
rect 20468 18652 20668 18680
rect 19751 18649 19763 18652
rect 19705 18643 19763 18649
rect 19797 18615 19855 18621
rect 19797 18612 19809 18615
rect 19444 18584 19809 18612
rect 19797 18581 19809 18584
rect 19843 18581 19855 18615
rect 19797 18575 19855 18581
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20254 18612 20260 18624
rect 20036 18584 20260 18612
rect 20036 18572 20042 18584
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20364 18612 20392 18652
rect 20533 18615 20591 18621
rect 20533 18612 20545 18615
rect 20364 18584 20545 18612
rect 20533 18581 20545 18584
rect 20579 18581 20591 18615
rect 20640 18612 20668 18652
rect 20901 18649 20913 18683
rect 20947 18649 20959 18683
rect 20901 18643 20959 18649
rect 21174 18640 21180 18692
rect 21232 18680 21238 18692
rect 22112 18680 22140 18779
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23256 18788 25176 18816
rect 23256 18776 23262 18788
rect 25148 18760 25176 18788
rect 26602 18776 26608 18828
rect 26660 18816 26666 18828
rect 26988 18825 27016 18856
rect 29012 18856 30696 18884
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 26660 18788 26709 18816
rect 26660 18776 26666 18788
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 26881 18819 26939 18825
rect 26881 18785 26893 18819
rect 26927 18785 26939 18819
rect 26881 18779 26939 18785
rect 26973 18819 27031 18825
rect 26973 18785 26985 18819
rect 27019 18785 27031 18819
rect 26973 18779 27031 18785
rect 27065 18819 27123 18825
rect 27065 18785 27077 18819
rect 27111 18816 27123 18819
rect 27111 18788 28856 18816
rect 27111 18785 27123 18788
rect 27065 18779 27123 18785
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18748 22615 18751
rect 22922 18748 22928 18760
rect 22603 18720 22928 18748
rect 22603 18717 22615 18720
rect 22557 18711 22615 18717
rect 21232 18652 22140 18680
rect 21232 18640 21238 18652
rect 20990 18612 20996 18624
rect 20640 18584 20996 18612
rect 20533 18575 20591 18581
rect 20990 18572 20996 18584
rect 21048 18572 21054 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 22094 18612 22100 18624
rect 21324 18584 22100 18612
rect 21324 18572 21330 18584
rect 22094 18572 22100 18584
rect 22152 18612 22158 18624
rect 22204 18612 22232 18711
rect 22296 18680 22324 18711
rect 22922 18708 22928 18720
rect 22980 18708 22986 18760
rect 24118 18708 24124 18760
rect 24176 18708 24182 18760
rect 24946 18708 24952 18760
rect 25004 18708 25010 18760
rect 25038 18708 25044 18760
rect 25096 18708 25102 18760
rect 25130 18708 25136 18760
rect 25188 18708 25194 18760
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 22646 18680 22652 18692
rect 22296 18652 22652 18680
rect 22646 18640 22652 18652
rect 22704 18680 22710 18692
rect 24136 18680 24164 18708
rect 22704 18652 24164 18680
rect 25240 18680 25268 18711
rect 26142 18708 26148 18760
rect 26200 18748 26206 18760
rect 26896 18748 26924 18779
rect 26200 18720 26924 18748
rect 27249 18751 27307 18757
rect 26200 18708 26206 18720
rect 27249 18717 27261 18751
rect 27295 18717 27307 18751
rect 28828 18748 28856 18788
rect 28902 18776 28908 18828
rect 28960 18776 28966 18828
rect 29012 18825 29040 18856
rect 28997 18819 29055 18825
rect 28997 18785 29009 18819
rect 29043 18785 29055 18819
rect 28997 18779 29055 18785
rect 29086 18776 29092 18828
rect 29144 18816 29150 18828
rect 29181 18819 29239 18825
rect 29181 18816 29193 18819
rect 29144 18788 29193 18816
rect 29144 18776 29150 18788
rect 29181 18785 29193 18788
rect 29227 18785 29239 18819
rect 29181 18779 29239 18785
rect 29914 18748 29920 18760
rect 28828 18720 29920 18748
rect 27249 18711 27307 18717
rect 27157 18683 27215 18689
rect 27157 18680 27169 18683
rect 25240 18652 27169 18680
rect 22704 18640 22710 18652
rect 27157 18649 27169 18652
rect 27203 18649 27215 18683
rect 27157 18643 27215 18649
rect 22152 18584 22232 18612
rect 22152 18572 22158 18584
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 24026 18612 24032 18624
rect 23532 18584 24032 18612
rect 23532 18572 23538 18584
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 26970 18612 26976 18624
rect 24912 18584 26976 18612
rect 24912 18572 24918 18584
rect 26970 18572 26976 18584
rect 27028 18612 27034 18624
rect 27264 18612 27292 18711
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 29089 18683 29147 18689
rect 29089 18649 29101 18683
rect 29135 18649 29147 18683
rect 29089 18643 29147 18649
rect 28166 18612 28172 18624
rect 27028 18584 28172 18612
rect 27028 18572 27034 18584
rect 28166 18572 28172 18584
rect 28224 18572 28230 18624
rect 28902 18572 28908 18624
rect 28960 18612 28966 18624
rect 29104 18612 29132 18643
rect 28960 18584 29132 18612
rect 28960 18572 28966 18584
rect 552 18522 31648 18544
rect 552 18470 4285 18522
rect 4337 18470 4349 18522
rect 4401 18470 4413 18522
rect 4465 18470 4477 18522
rect 4529 18470 4541 18522
rect 4593 18470 12059 18522
rect 12111 18470 12123 18522
rect 12175 18470 12187 18522
rect 12239 18470 12251 18522
rect 12303 18470 12315 18522
rect 12367 18470 19833 18522
rect 19885 18470 19897 18522
rect 19949 18470 19961 18522
rect 20013 18470 20025 18522
rect 20077 18470 20089 18522
rect 20141 18470 27607 18522
rect 27659 18470 27671 18522
rect 27723 18470 27735 18522
rect 27787 18470 27799 18522
rect 27851 18470 27863 18522
rect 27915 18470 31648 18522
rect 552 18448 31648 18470
rect 2590 18368 2596 18420
rect 2648 18408 2654 18420
rect 2774 18408 2780 18420
rect 2648 18380 2780 18408
rect 2648 18368 2654 18380
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3050 18368 3056 18420
rect 3108 18368 3114 18420
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 3789 18411 3847 18417
rect 3789 18408 3801 18411
rect 3568 18380 3801 18408
rect 3568 18368 3574 18380
rect 3789 18377 3801 18380
rect 3835 18377 3847 18411
rect 4890 18408 4896 18420
rect 3789 18371 3847 18377
rect 3896 18380 4896 18408
rect 2869 18343 2927 18349
rect 2869 18340 2881 18343
rect 2746 18312 2881 18340
rect 1026 18232 1032 18284
rect 1084 18232 1090 18284
rect 1305 18275 1363 18281
rect 1305 18241 1317 18275
rect 1351 18272 1363 18275
rect 2746 18272 2774 18312
rect 2869 18309 2881 18312
rect 2915 18309 2927 18343
rect 2869 18303 2927 18309
rect 1351 18244 2774 18272
rect 1351 18241 1363 18244
rect 1305 18235 1363 18241
rect 3068 18213 3096 18368
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 3896 18340 3924 18380
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 4982 18368 4988 18420
rect 5040 18368 5046 18420
rect 5442 18408 5448 18420
rect 5092 18380 5448 18408
rect 3292 18312 3924 18340
rect 3292 18300 3298 18312
rect 3436 18213 3464 18312
rect 4154 18300 4160 18352
rect 4212 18300 4218 18352
rect 5000 18340 5028 18368
rect 4264 18312 5028 18340
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3053 18167 3111 18173
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18173 3479 18207
rect 3528 18204 3556 18235
rect 3602 18232 3608 18284
rect 3660 18272 3666 18284
rect 3660 18244 3924 18272
rect 3660 18232 3666 18244
rect 3896 18213 3924 18244
rect 4264 18213 4292 18312
rect 4982 18272 4988 18284
rect 4356 18244 4988 18272
rect 3881 18207 3939 18213
rect 3528 18176 3648 18204
rect 3421 18167 3479 18173
rect 2682 18136 2688 18148
rect 2530 18108 2688 18136
rect 2682 18096 2688 18108
rect 2740 18096 2746 18148
rect 3326 18096 3332 18148
rect 3384 18136 3390 18148
rect 3620 18136 3648 18176
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 3927 18176 4261 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 4249 18173 4261 18176
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 3384 18108 3648 18136
rect 3384 18096 3390 18108
rect 3620 18068 3648 18108
rect 3786 18096 3792 18148
rect 3844 18136 3850 18148
rect 3973 18139 4031 18145
rect 3973 18136 3985 18139
rect 3844 18108 3985 18136
rect 3844 18096 3850 18108
rect 3973 18105 3985 18108
rect 4019 18105 4031 18139
rect 3973 18099 4031 18105
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 4157 18139 4215 18145
rect 4157 18136 4169 18139
rect 4120 18108 4169 18136
rect 4120 18096 4126 18108
rect 4157 18105 4169 18108
rect 4203 18136 4215 18139
rect 4356 18136 4384 18244
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5092 18281 5120 18380
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 5626 18368 5632 18420
rect 5684 18368 5690 18420
rect 5718 18368 5724 18420
rect 5776 18368 5782 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 10502 18408 10508 18420
rect 8251 18380 10508 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 10962 18368 10968 18420
rect 11020 18368 11026 18420
rect 11054 18368 11060 18420
rect 11112 18368 11118 18420
rect 11241 18411 11299 18417
rect 11241 18377 11253 18411
rect 11287 18408 11299 18411
rect 11606 18408 11612 18420
rect 11287 18380 11612 18408
rect 11287 18377 11299 18380
rect 11241 18371 11299 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 15838 18408 15844 18420
rect 12268 18380 15844 18408
rect 5184 18312 6040 18340
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5077 18235 5135 18241
rect 5184 18204 5212 18312
rect 6012 18272 6040 18312
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 8352 18312 8708 18340
rect 8352 18300 8358 18312
rect 6012 18244 8248 18272
rect 4540 18176 5212 18204
rect 4203 18108 4384 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4430 18096 4436 18148
rect 4488 18096 4494 18148
rect 4540 18068 4568 18176
rect 5350 18164 5356 18216
rect 5408 18204 5414 18216
rect 6012 18213 6040 18244
rect 5905 18207 5963 18213
rect 5905 18204 5917 18207
rect 5408 18176 5917 18204
rect 5408 18164 5414 18176
rect 5905 18173 5917 18176
rect 5951 18173 5963 18207
rect 5905 18167 5963 18173
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18173 6055 18207
rect 5997 18167 6055 18173
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 6178 18164 6184 18216
rect 6236 18164 6242 18216
rect 8220 18213 8248 18244
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8444 18244 8585 18272
rect 8444 18232 8450 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8680 18272 8708 18312
rect 10318 18300 10324 18352
rect 10376 18300 10382 18352
rect 11072 18340 11100 18368
rect 11422 18340 11428 18352
rect 11072 18312 11428 18340
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11790 18300 11796 18352
rect 11848 18300 11854 18352
rect 12268 18281 12296 18380
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 17034 18368 17040 18420
rect 17092 18368 17098 18420
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 17405 18411 17463 18417
rect 17405 18408 17417 18411
rect 17276 18380 17417 18408
rect 17276 18368 17282 18380
rect 17405 18377 17417 18380
rect 17451 18377 17463 18411
rect 17405 18371 17463 18377
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 17552 18380 19472 18408
rect 17552 18368 17558 18380
rect 12618 18340 12624 18352
rect 12544 18312 12624 18340
rect 12544 18281 12572 18312
rect 12618 18300 12624 18312
rect 12676 18300 12682 18352
rect 12986 18340 12992 18352
rect 12728 18312 12992 18340
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 8680 18244 11192 18272
rect 8573 18235 8631 18241
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18173 8079 18207
rect 8021 18167 8079 18173
rect 8205 18207 8263 18213
rect 8205 18173 8217 18207
rect 8251 18173 8263 18207
rect 8205 18167 8263 18173
rect 5711 18139 5769 18145
rect 5711 18105 5723 18139
rect 5757 18136 5769 18139
rect 6104 18136 6132 18164
rect 6457 18139 6515 18145
rect 6457 18136 6469 18139
rect 5757 18108 6040 18136
rect 6104 18108 6469 18136
rect 5757 18105 5769 18108
rect 5711 18099 5769 18105
rect 6012 18080 6040 18108
rect 6457 18105 6469 18108
rect 6503 18105 6515 18139
rect 6457 18099 6515 18105
rect 7466 18096 7472 18148
rect 7524 18096 7530 18148
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 8036 18136 8064 18167
rect 7800 18108 8064 18136
rect 8220 18136 8248 18167
rect 9950 18164 9956 18216
rect 10008 18164 10014 18216
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18204 10655 18207
rect 10686 18204 10692 18216
rect 10643 18176 10692 18204
rect 10643 18173 10655 18176
rect 10597 18167 10655 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11164 18213 11192 18244
rect 11900 18244 12173 18272
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 11149 18207 11207 18213
rect 10919 18176 11008 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 8570 18136 8576 18148
rect 8220 18108 8576 18136
rect 7800 18096 7806 18108
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18105 8907 18139
rect 10336 18136 10364 18164
rect 10781 18139 10839 18145
rect 10781 18136 10793 18139
rect 10336 18108 10793 18136
rect 8849 18099 8907 18105
rect 3620 18040 4568 18068
rect 4614 18028 4620 18080
rect 4672 18028 4678 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5169 18071 5227 18077
rect 5169 18068 5181 18071
rect 4856 18040 5181 18068
rect 4856 18028 4862 18040
rect 5169 18037 5181 18040
rect 5215 18037 5227 18071
rect 5169 18031 5227 18037
rect 5258 18028 5264 18080
rect 5316 18028 5322 18080
rect 5994 18028 6000 18080
rect 6052 18028 6058 18080
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 7834 18068 7840 18080
rect 7248 18040 7840 18068
rect 7248 18028 7254 18040
rect 7834 18028 7840 18040
rect 7892 18068 7898 18080
rect 7929 18071 7987 18077
rect 7929 18068 7941 18071
rect 7892 18040 7941 18068
rect 7892 18028 7898 18040
rect 7929 18037 7941 18040
rect 7975 18037 7987 18071
rect 8864 18068 8892 18099
rect 10612 18080 10640 18108
rect 10781 18105 10793 18108
rect 10827 18105 10839 18139
rect 10781 18099 10839 18105
rect 10980 18080 11008 18176
rect 11149 18173 11161 18207
rect 11195 18173 11207 18207
rect 11149 18167 11207 18173
rect 11422 18164 11428 18216
rect 11480 18164 11486 18216
rect 11606 18164 11612 18216
rect 11664 18164 11670 18216
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 11790 18204 11796 18216
rect 11747 18176 11796 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11900 18136 11928 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 12544 18204 12572 18235
rect 12023 18176 12572 18204
rect 12621 18207 12679 18213
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 12728 18204 12756 18312
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 14829 18343 14887 18349
rect 14829 18340 14841 18343
rect 13096 18312 14841 18340
rect 13096 18272 13124 18312
rect 14829 18309 14841 18312
rect 14875 18309 14887 18343
rect 14829 18303 14887 18309
rect 15102 18300 15108 18352
rect 15160 18300 15166 18352
rect 15194 18300 15200 18352
rect 15252 18340 15258 18352
rect 19444 18340 19472 18380
rect 19518 18368 19524 18420
rect 19576 18368 19582 18420
rect 19610 18368 19616 18420
rect 19668 18368 19674 18420
rect 20438 18368 20444 18420
rect 20496 18368 20502 18420
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 22370 18408 22376 18420
rect 20772 18380 22376 18408
rect 20772 18368 20778 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 24029 18411 24087 18417
rect 24029 18408 24041 18411
rect 22480 18380 24041 18408
rect 22480 18352 22508 18380
rect 24029 18377 24041 18380
rect 24075 18408 24087 18411
rect 24118 18408 24124 18420
rect 24075 18380 24124 18408
rect 24075 18377 24087 18380
rect 24029 18371 24087 18377
rect 24118 18368 24124 18380
rect 24176 18368 24182 18420
rect 24486 18368 24492 18420
rect 24544 18408 24550 18420
rect 24765 18411 24823 18417
rect 24765 18408 24777 18411
rect 24544 18380 24777 18408
rect 24544 18368 24550 18380
rect 24765 18377 24777 18380
rect 24811 18377 24823 18411
rect 24765 18371 24823 18377
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 24949 18411 25007 18417
rect 24949 18408 24961 18411
rect 24912 18380 24961 18408
rect 24912 18368 24918 18380
rect 24949 18377 24961 18380
rect 24995 18408 25007 18411
rect 26142 18408 26148 18420
rect 24995 18380 26148 18408
rect 24995 18377 25007 18380
rect 24949 18371 25007 18377
rect 26142 18368 26148 18380
rect 26200 18368 26206 18420
rect 26694 18368 26700 18420
rect 26752 18408 26758 18420
rect 27525 18411 27583 18417
rect 27525 18408 27537 18411
rect 26752 18380 27537 18408
rect 26752 18368 26758 18380
rect 27525 18377 27537 18380
rect 27571 18377 27583 18411
rect 27525 18371 27583 18377
rect 29270 18368 29276 18420
rect 29328 18408 29334 18420
rect 29365 18411 29423 18417
rect 29365 18408 29377 18411
rect 29328 18380 29377 18408
rect 29328 18368 29334 18380
rect 29365 18377 29377 18380
rect 29411 18408 29423 18411
rect 29546 18408 29552 18420
rect 29411 18380 29552 18408
rect 29411 18377 29423 18380
rect 29365 18371 29423 18377
rect 29546 18368 29552 18380
rect 29604 18368 29610 18420
rect 30190 18368 30196 18420
rect 30248 18368 30254 18420
rect 30466 18368 30472 18420
rect 30524 18368 30530 18420
rect 20254 18340 20260 18352
rect 15252 18312 19272 18340
rect 19444 18312 20260 18340
rect 15252 18300 15258 18312
rect 12667 18176 12756 18204
rect 12820 18244 13124 18272
rect 13173 18275 13231 18281
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 12342 18136 12348 18148
rect 11900 18108 12348 18136
rect 12342 18096 12348 18108
rect 12400 18136 12406 18148
rect 12820 18136 12848 18244
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 13219 18244 14105 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18272 14427 18275
rect 15120 18272 15148 18300
rect 14415 18244 15148 18272
rect 14415 18241 14427 18244
rect 14369 18235 14427 18241
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13262 18204 13268 18216
rect 13035 18176 13268 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 12400 18108 12848 18136
rect 12912 18136 12940 18167
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13906 18164 13912 18216
rect 13964 18164 13970 18216
rect 14001 18207 14059 18213
rect 14001 18173 14013 18207
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18204 14243 18207
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14231 18176 14473 18204
rect 14231 18173 14243 18176
rect 14185 18167 14243 18173
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 14016 18136 14044 18167
rect 14642 18164 14648 18216
rect 14700 18164 14706 18216
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 14752 18136 14780 18167
rect 14918 18164 14924 18216
rect 14976 18164 14982 18216
rect 15010 18164 15016 18216
rect 15068 18164 15074 18216
rect 15212 18213 15240 18300
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15378 18164 15384 18216
rect 15436 18164 15442 18216
rect 15470 18164 15476 18216
rect 15528 18164 15534 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 15654 18204 15660 18216
rect 15611 18176 15660 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 15856 18204 15884 18235
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16172 18244 18920 18272
rect 16172 18232 16178 18244
rect 15933 18207 15991 18213
rect 15933 18204 15945 18207
rect 15856 18176 15945 18204
rect 15933 18173 15945 18176
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 16022 18164 16028 18216
rect 16080 18164 16086 18216
rect 16209 18207 16267 18213
rect 16209 18173 16221 18207
rect 16255 18204 16267 18207
rect 16255 18176 16804 18204
rect 16255 18173 16267 18176
rect 16209 18167 16267 18173
rect 15028 18136 15056 18164
rect 12912 18108 13492 18136
rect 14016 18108 14504 18136
rect 14752 18108 15056 18136
rect 15396 18136 15424 18164
rect 16776 18148 16804 18176
rect 16850 18164 16856 18216
rect 16908 18164 16914 18216
rect 16942 18164 16948 18216
rect 17000 18204 17006 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 17000 18176 17141 18204
rect 17000 18164 17006 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 17218 18164 17224 18216
rect 17276 18204 17282 18216
rect 17862 18204 17868 18216
rect 17276 18176 17868 18204
rect 17276 18164 17282 18176
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 18690 18164 18696 18216
rect 18748 18204 18754 18216
rect 18892 18213 18920 18244
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19024 18244 19196 18272
rect 19024 18232 19030 18244
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 18748 18176 18797 18204
rect 18748 18164 18754 18176
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 18877 18207 18935 18213
rect 18877 18173 18889 18207
rect 18923 18173 18935 18207
rect 18877 18167 18935 18173
rect 19058 18164 19064 18216
rect 19116 18164 19122 18216
rect 19168 18213 19196 18244
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19244 18204 19272 18312
rect 20254 18300 20260 18312
rect 20312 18340 20318 18352
rect 20312 18312 20484 18340
rect 20312 18300 20318 18312
rect 20456 18281 20484 18312
rect 20622 18300 20628 18352
rect 20680 18300 20686 18352
rect 20806 18300 20812 18352
rect 20864 18300 20870 18352
rect 21266 18300 21272 18352
rect 21324 18340 21330 18352
rect 22462 18340 22468 18352
rect 21324 18312 22468 18340
rect 21324 18300 21330 18312
rect 22462 18300 22468 18312
rect 22520 18300 22526 18352
rect 23014 18340 23020 18352
rect 22664 18312 23020 18340
rect 19337 18280 19395 18281
rect 19425 18280 19483 18281
rect 19337 18275 19483 18280
rect 19337 18241 19349 18275
rect 19383 18252 19437 18275
rect 19383 18241 19395 18252
rect 19337 18235 19395 18241
rect 19425 18241 19437 18252
rect 19471 18241 19483 18275
rect 20441 18275 20499 18281
rect 19425 18235 19483 18241
rect 19536 18244 20024 18272
rect 19536 18204 19564 18244
rect 19702 18204 19708 18216
rect 19244 18176 19564 18204
rect 19628 18176 19708 18204
rect 19153 18167 19211 18173
rect 15396 18108 16620 18136
rect 12400 18096 12406 18108
rect 13464 18080 13492 18108
rect 9674 18068 9680 18080
rect 8864 18040 9680 18068
rect 7929 18031 7987 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10410 18028 10416 18080
rect 10468 18028 10474 18080
rect 10594 18028 10600 18080
rect 10652 18028 10658 18080
rect 10962 18028 10968 18080
rect 11020 18028 11026 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12032 18040 12725 18068
rect 12032 18028 12038 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12713 18031 12771 18037
rect 13446 18028 13452 18080
rect 13504 18028 13510 18080
rect 14476 18068 14504 18108
rect 16592 18080 16620 18108
rect 16758 18096 16764 18148
rect 16816 18096 16822 18148
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 17736 18108 19272 18136
rect 17736 18096 17742 18108
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 14476 18040 15945 18068
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16482 18068 16488 18080
rect 16080 18040 16488 18068
rect 16080 18028 16086 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 16574 18028 16580 18080
rect 16632 18028 16638 18080
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17586 18068 17592 18080
rect 17276 18040 17592 18068
rect 17276 18028 17282 18040
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 18506 18028 18512 18080
rect 18564 18068 18570 18080
rect 19150 18068 19156 18080
rect 18564 18040 19156 18068
rect 18564 18028 18570 18040
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 19244 18068 19272 18108
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 19628 18136 19656 18176
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 19996 18204 20024 18244
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20640 18272 20668 18300
rect 20640 18244 20760 18272
rect 20441 18235 20499 18241
rect 20548 18213 20668 18214
rect 20548 18207 20683 18213
rect 20548 18206 20637 18207
rect 20468 18204 20637 18206
rect 19996 18186 20637 18204
rect 19996 18178 20576 18186
rect 19996 18176 20496 18178
rect 19392 18108 19656 18136
rect 19392 18096 19398 18108
rect 20070 18096 20076 18148
rect 20128 18136 20134 18148
rect 20349 18139 20407 18145
rect 20349 18136 20361 18139
rect 20128 18108 20361 18136
rect 20128 18096 20134 18108
rect 20349 18105 20361 18108
rect 20395 18105 20407 18139
rect 20548 18136 20576 18178
rect 20625 18173 20637 18186
rect 20671 18173 20683 18207
rect 20732 18204 20760 18244
rect 22664 18213 22692 18312
rect 23014 18300 23020 18312
rect 23072 18300 23078 18352
rect 23201 18343 23259 18349
rect 23201 18309 23213 18343
rect 23247 18340 23259 18343
rect 25866 18340 25872 18352
rect 23247 18312 25872 18340
rect 23247 18309 23259 18312
rect 23201 18303 23259 18309
rect 25866 18300 25872 18312
rect 25924 18300 25930 18352
rect 26234 18300 26240 18352
rect 26292 18340 26298 18352
rect 28074 18340 28080 18352
rect 26292 18312 28080 18340
rect 26292 18300 26298 18312
rect 22738 18232 22744 18284
rect 22796 18232 22802 18284
rect 23106 18232 23112 18284
rect 23164 18272 23170 18284
rect 24302 18272 24308 18284
rect 23164 18244 24308 18272
rect 23164 18232 23170 18244
rect 24302 18232 24308 18244
rect 24360 18232 24366 18284
rect 24486 18232 24492 18284
rect 24544 18272 24550 18284
rect 24673 18275 24731 18281
rect 24673 18272 24685 18275
rect 24544 18244 24685 18272
rect 24544 18232 24550 18244
rect 24673 18241 24685 18244
rect 24719 18272 24731 18275
rect 25041 18275 25099 18281
rect 25041 18272 25053 18275
rect 24719 18244 25053 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 25041 18241 25053 18244
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 26697 18275 26755 18281
rect 26697 18241 26709 18275
rect 26743 18272 26755 18275
rect 27246 18272 27252 18284
rect 26743 18244 27252 18272
rect 26743 18241 26755 18244
rect 26697 18235 26755 18241
rect 27246 18232 27252 18244
rect 27304 18232 27310 18284
rect 27338 18232 27344 18284
rect 27396 18272 27402 18284
rect 27396 18244 27522 18272
rect 27396 18232 27402 18244
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 20732 18176 22661 18204
rect 20625 18167 20683 18173
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 22830 18164 22836 18216
rect 22888 18204 22894 18216
rect 22925 18207 22983 18213
rect 22925 18204 22937 18207
rect 22888 18176 22937 18204
rect 22888 18164 22894 18176
rect 22925 18173 22937 18176
rect 22971 18173 22983 18207
rect 22925 18167 22983 18173
rect 23014 18164 23020 18216
rect 23072 18164 23078 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 23750 18204 23756 18216
rect 23532 18176 23756 18204
rect 23532 18164 23538 18176
rect 23750 18164 23756 18176
rect 23808 18204 23814 18216
rect 23937 18207 23995 18213
rect 23937 18204 23949 18207
rect 23808 18176 23949 18204
rect 23808 18164 23814 18176
rect 23937 18173 23949 18176
rect 23983 18173 23995 18207
rect 23937 18167 23995 18173
rect 24026 18164 24032 18216
rect 24084 18204 24090 18216
rect 24397 18207 24455 18213
rect 24397 18204 24409 18207
rect 24084 18176 24409 18204
rect 24084 18164 24090 18176
rect 24397 18173 24409 18176
rect 24443 18173 24455 18207
rect 24397 18167 24455 18173
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 24949 18207 25007 18213
rect 24949 18204 24961 18207
rect 24912 18176 24961 18204
rect 24912 18164 24918 18176
rect 24949 18173 24961 18176
rect 24995 18173 25007 18207
rect 24949 18167 25007 18173
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25271 18176 27384 18204
rect 27494 18179 27522 18244
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 24044 18136 24072 18164
rect 20548 18108 24072 18136
rect 24213 18139 24271 18145
rect 20349 18099 20407 18105
rect 24213 18105 24225 18139
rect 24259 18136 24271 18139
rect 24670 18136 24676 18148
rect 24259 18108 24676 18136
rect 24259 18105 24271 18108
rect 24213 18099 24271 18105
rect 24670 18096 24676 18108
rect 24728 18096 24734 18148
rect 25406 18136 25412 18148
rect 24872 18108 25412 18136
rect 20990 18068 20996 18080
rect 19244 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18068 21054 18080
rect 21910 18068 21916 18080
rect 21048 18040 21916 18068
rect 21048 18028 21054 18040
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 24872 18068 24900 18108
rect 25406 18096 25412 18108
rect 25464 18136 25470 18148
rect 25682 18136 25688 18148
rect 25464 18108 25688 18136
rect 25464 18096 25470 18108
rect 25682 18096 25688 18108
rect 25740 18096 25746 18148
rect 25866 18096 25872 18148
rect 25924 18136 25930 18148
rect 26697 18139 26755 18145
rect 26697 18136 26709 18139
rect 25924 18108 26709 18136
rect 25924 18096 25930 18108
rect 26697 18105 26709 18108
rect 26743 18105 26755 18139
rect 26697 18099 26755 18105
rect 26789 18139 26847 18145
rect 26789 18105 26801 18139
rect 26835 18136 26847 18139
rect 26970 18136 26976 18148
rect 26835 18108 26976 18136
rect 26835 18105 26847 18108
rect 26789 18099 26847 18105
rect 26970 18096 26976 18108
rect 27028 18096 27034 18148
rect 24351 18040 24900 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 27356 18077 27384 18176
rect 27479 18173 27537 18179
rect 27479 18139 27491 18173
rect 27525 18139 27537 18173
rect 27479 18133 27537 18139
rect 27632 18136 27660 18312
rect 28074 18300 28080 18312
rect 28132 18300 28138 18352
rect 30208 18272 30236 18368
rect 30377 18275 30435 18281
rect 30377 18272 30389 18275
rect 30208 18244 30389 18272
rect 30377 18241 30389 18244
rect 30423 18241 30435 18275
rect 30484 18272 30512 18368
rect 30561 18275 30619 18281
rect 30561 18272 30573 18275
rect 30484 18244 30573 18272
rect 30377 18235 30435 18241
rect 30561 18241 30573 18244
rect 30607 18241 30619 18275
rect 30561 18235 30619 18241
rect 28626 18164 28632 18216
rect 28684 18204 28690 18216
rect 30098 18204 30104 18216
rect 28684 18176 30104 18204
rect 28684 18164 28690 18176
rect 30098 18164 30104 18176
rect 30156 18204 30162 18216
rect 30469 18207 30527 18213
rect 30469 18204 30481 18207
rect 30156 18176 30481 18204
rect 30156 18164 30162 18176
rect 30469 18173 30481 18176
rect 30515 18173 30527 18207
rect 30469 18167 30527 18173
rect 30650 18164 30656 18216
rect 30708 18164 30714 18216
rect 27709 18139 27767 18145
rect 27709 18136 27721 18139
rect 27632 18108 27721 18136
rect 27709 18105 27721 18108
rect 27755 18105 27767 18139
rect 27709 18099 27767 18105
rect 27798 18096 27804 18148
rect 27856 18136 27862 18148
rect 29089 18139 29147 18145
rect 29089 18136 29101 18139
rect 27856 18108 29101 18136
rect 27856 18096 27862 18108
rect 29089 18105 29101 18108
rect 29135 18136 29147 18139
rect 30006 18136 30012 18148
rect 29135 18108 30012 18136
rect 29135 18105 29147 18108
rect 29089 18099 29147 18105
rect 30006 18096 30012 18108
rect 30064 18096 30070 18148
rect 26219 18071 26277 18077
rect 26219 18068 26231 18071
rect 25280 18040 26231 18068
rect 25280 18028 25286 18040
rect 26219 18037 26231 18040
rect 26265 18037 26277 18071
rect 26219 18031 26277 18037
rect 27341 18071 27399 18077
rect 27341 18037 27353 18071
rect 27387 18037 27399 18071
rect 27341 18031 27399 18037
rect 30193 18071 30251 18077
rect 30193 18037 30205 18071
rect 30239 18068 30251 18071
rect 30466 18068 30472 18080
rect 30239 18040 30472 18068
rect 30239 18037 30251 18040
rect 30193 18031 30251 18037
rect 30466 18028 30472 18040
rect 30524 18028 30530 18080
rect 552 17978 31808 18000
rect 552 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 15946 17978
rect 15998 17926 16010 17978
rect 16062 17926 16074 17978
rect 16126 17926 16138 17978
rect 16190 17926 16202 17978
rect 16254 17926 23720 17978
rect 23772 17926 23784 17978
rect 23836 17926 23848 17978
rect 23900 17926 23912 17978
rect 23964 17926 23976 17978
rect 24028 17926 31494 17978
rect 31546 17926 31558 17978
rect 31610 17926 31622 17978
rect 31674 17926 31686 17978
rect 31738 17926 31750 17978
rect 31802 17926 31808 17978
rect 552 17904 31808 17926
rect 860 17836 2728 17864
rect 860 17737 888 17836
rect 2590 17796 2596 17808
rect 2346 17768 2596 17796
rect 2590 17756 2596 17768
rect 2648 17756 2654 17808
rect 2700 17740 2728 17836
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3786 17864 3792 17876
rect 2832 17836 3792 17864
rect 2832 17824 2838 17836
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 3970 17824 3976 17876
rect 4028 17864 4034 17876
rect 4028 17836 4108 17864
rect 4028 17824 4034 17836
rect 845 17731 903 17737
rect 845 17697 857 17731
rect 891 17697 903 17731
rect 845 17691 903 17697
rect 2682 17688 2688 17740
rect 2740 17688 2746 17740
rect 4080 17714 4108 17836
rect 5810 17824 5816 17876
rect 5868 17864 5874 17876
rect 6273 17867 6331 17873
rect 6273 17864 6285 17867
rect 5868 17836 6285 17864
rect 5868 17824 5874 17836
rect 6273 17833 6285 17836
rect 6319 17833 6331 17867
rect 6822 17864 6828 17876
rect 6273 17827 6331 17833
rect 6380 17836 6828 17864
rect 4522 17756 4528 17808
rect 4580 17796 4586 17808
rect 4580 17768 5120 17796
rect 4580 17756 4586 17768
rect 4430 17688 4436 17740
rect 4488 17728 4494 17740
rect 5092 17737 5120 17768
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 6380 17796 6408 17836
rect 6822 17824 6828 17836
rect 6880 17864 6886 17876
rect 7742 17864 7748 17876
rect 6880 17836 7748 17864
rect 6880 17824 6886 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 7837 17867 7895 17873
rect 7837 17833 7849 17867
rect 7883 17864 7895 17867
rect 8018 17864 8024 17876
rect 7883 17836 8024 17864
rect 7883 17833 7895 17836
rect 7837 17827 7895 17833
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 8662 17864 8668 17876
rect 8404 17836 8668 17864
rect 5684 17768 6408 17796
rect 6641 17799 6699 17805
rect 5684 17756 5690 17768
rect 6641 17765 6653 17799
rect 6687 17796 6699 17799
rect 7190 17796 7196 17808
rect 6687 17768 7196 17796
rect 6687 17765 6699 17768
rect 6641 17759 6699 17765
rect 7190 17756 7196 17768
rect 7248 17756 7254 17808
rect 8189 17799 8247 17805
rect 8189 17765 8201 17799
rect 8235 17796 8247 17799
rect 8294 17796 8300 17808
rect 8235 17768 8300 17796
rect 8235 17765 8247 17768
rect 8189 17759 8247 17765
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 8404 17805 8432 17836
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 9030 17864 9036 17876
rect 8869 17836 9036 17864
rect 8869 17805 8897 17836
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9140 17836 9720 17864
rect 8389 17799 8447 17805
rect 8389 17765 8401 17799
rect 8435 17765 8447 17799
rect 8849 17799 8907 17805
rect 8389 17759 8447 17765
rect 8496 17768 8708 17796
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4488 17700 4813 17728
rect 4488 17688 4494 17700
rect 4801 17697 4813 17700
rect 4847 17697 4859 17731
rect 4801 17691 4859 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17697 4951 17731
rect 4893 17691 4951 17697
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 6733 17731 6791 17737
rect 6733 17697 6745 17731
rect 6779 17728 6791 17731
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 6779 17700 7389 17728
rect 6779 17697 6791 17700
rect 6733 17691 6791 17697
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 1118 17620 1124 17672
rect 1176 17620 1182 17672
rect 2958 17620 2964 17672
rect 3016 17620 3022 17672
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4908 17660 4936 17691
rect 4028 17632 4936 17660
rect 4028 17620 4034 17632
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 5537 17663 5595 17669
rect 5537 17660 5549 17663
rect 5500 17632 5549 17660
rect 5500 17620 5506 17632
rect 5537 17629 5549 17632
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 6104 17592 6132 17691
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 6748 17660 6776 17691
rect 7466 17688 7472 17740
rect 7524 17688 7530 17740
rect 8496 17737 8524 17768
rect 8481 17731 8539 17737
rect 8128 17700 8340 17728
rect 6512 17632 6776 17660
rect 6825 17663 6883 17669
rect 6512 17620 6518 17632
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 7098 17660 7104 17672
rect 6871 17632 7104 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 8128 17592 8156 17700
rect 3988 17564 4936 17592
rect 6104 17564 8156 17592
rect 2593 17527 2651 17533
rect 2593 17493 2605 17527
rect 2639 17524 2651 17527
rect 3050 17524 3056 17536
rect 2639 17496 3056 17524
rect 2639 17493 2651 17496
rect 2593 17487 2651 17493
rect 3050 17484 3056 17496
rect 3108 17524 3114 17536
rect 3694 17524 3700 17536
rect 3108 17496 3700 17524
rect 3108 17484 3114 17496
rect 3694 17484 3700 17496
rect 3752 17524 3758 17536
rect 3988 17524 4016 17564
rect 4908 17536 4936 17564
rect 3752 17496 4016 17524
rect 4433 17527 4491 17533
rect 3752 17484 3758 17496
rect 4433 17493 4445 17527
rect 4479 17524 4491 17527
rect 4706 17524 4712 17536
rect 4479 17496 4712 17524
rect 4479 17493 4491 17496
rect 4433 17487 4491 17493
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 4890 17484 4896 17536
rect 4948 17484 4954 17536
rect 5902 17484 5908 17536
rect 5960 17484 5966 17536
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7834 17524 7840 17536
rect 6788 17496 7840 17524
rect 6788 17484 6794 17496
rect 7834 17484 7840 17496
rect 7892 17524 7898 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7892 17496 8033 17524
rect 7892 17484 7898 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 8202 17484 8208 17536
rect 8260 17484 8266 17536
rect 8312 17524 8340 17700
rect 8481 17697 8493 17731
rect 8527 17697 8539 17731
rect 8481 17691 8539 17697
rect 8574 17731 8632 17737
rect 8574 17697 8586 17731
rect 8620 17697 8632 17731
rect 8574 17691 8632 17697
rect 8588 17660 8616 17691
rect 8497 17632 8616 17660
rect 8680 17660 8708 17768
rect 8849 17765 8861 17799
rect 8895 17765 8907 17799
rect 8849 17759 8907 17765
rect 8754 17688 8760 17740
rect 8812 17688 8818 17740
rect 8987 17731 9045 17737
rect 8987 17697 8999 17731
rect 9033 17728 9045 17731
rect 9140 17728 9168 17836
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 9493 17799 9551 17805
rect 9493 17796 9505 17799
rect 9456 17768 9505 17796
rect 9456 17756 9462 17768
rect 9493 17765 9505 17768
rect 9539 17765 9551 17799
rect 9493 17759 9551 17765
rect 9033 17700 9168 17728
rect 9033 17697 9045 17700
rect 8987 17691 9045 17697
rect 9214 17688 9220 17740
rect 9272 17688 9278 17740
rect 9310 17731 9368 17737
rect 9310 17697 9322 17731
rect 9356 17697 9368 17731
rect 9310 17691 9368 17697
rect 9232 17660 9260 17688
rect 8680 17632 9260 17660
rect 9325 17660 9353 17691
rect 9582 17688 9588 17740
rect 9640 17688 9646 17740
rect 9692 17737 9720 17836
rect 9950 17824 9956 17876
rect 10008 17824 10014 17876
rect 10410 17864 10416 17876
rect 10336 17836 10416 17864
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 10336 17805 10364 17836
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 12342 17873 12348 17876
rect 11885 17867 11943 17873
rect 11885 17864 11897 17867
rect 10652 17836 11897 17864
rect 10652 17824 10658 17836
rect 10321 17799 10379 17805
rect 9916 17768 10272 17796
rect 9916 17756 9922 17768
rect 10134 17737 10140 17740
rect 9682 17731 9740 17737
rect 9682 17697 9694 17731
rect 9728 17718 9740 17731
rect 10132 17728 10140 17737
rect 9876 17718 10140 17728
rect 9728 17700 10140 17718
rect 9728 17697 9904 17700
rect 9682 17691 9904 17697
rect 10132 17691 10140 17700
rect 9692 17690 9904 17691
rect 10134 17688 10140 17691
rect 10192 17688 10198 17740
rect 10244 17737 10272 17768
rect 10321 17765 10333 17799
rect 10367 17765 10379 17799
rect 10321 17759 10379 17765
rect 10962 17756 10968 17808
rect 11020 17796 11026 17808
rect 11348 17805 11376 17836
rect 11885 17833 11897 17836
rect 11931 17833 11943 17867
rect 12338 17864 12348 17873
rect 12303 17836 12348 17864
rect 11885 17827 11943 17833
rect 12338 17827 12348 17836
rect 12342 17824 12348 17827
rect 12400 17824 12406 17876
rect 16574 17864 16580 17876
rect 15166 17836 16580 17864
rect 11117 17799 11175 17805
rect 11117 17796 11129 17799
rect 11020 17768 11129 17796
rect 11020 17756 11026 17768
rect 11117 17765 11129 17768
rect 11163 17765 11175 17799
rect 11117 17759 11175 17765
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17765 11391 17799
rect 11333 17759 11391 17765
rect 11422 17756 11428 17808
rect 11480 17796 11486 17808
rect 12253 17799 12311 17805
rect 11480 17768 12204 17796
rect 11480 17756 11486 17768
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10502 17728 10508 17740
rect 10463 17700 10508 17728
rect 10229 17691 10287 17697
rect 10502 17688 10508 17700
rect 10560 17688 10566 17740
rect 10594 17688 10600 17740
rect 10652 17688 10658 17740
rect 10778 17688 10784 17740
rect 10836 17728 10842 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 10836 17700 11713 17728
rect 10836 17688 10842 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 11790 17688 11796 17740
rect 11848 17688 11854 17740
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12176 17737 12204 17768
rect 12253 17765 12265 17799
rect 12299 17796 12311 17799
rect 12618 17796 12624 17808
rect 12299 17768 12624 17796
rect 12299 17765 12311 17768
rect 12253 17759 12311 17765
rect 12618 17756 12624 17768
rect 12676 17796 12682 17808
rect 15166 17796 15194 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16942 17824 16948 17876
rect 17000 17824 17006 17876
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17833 17371 17867
rect 17313 17827 17371 17833
rect 17328 17796 17356 17827
rect 17770 17824 17776 17876
rect 17828 17864 17834 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17828 17836 17877 17864
rect 17828 17824 17834 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 18506 17864 18512 17876
rect 17865 17827 17923 17833
rect 17972 17836 18512 17864
rect 17972 17796 18000 17836
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 18748 17836 19564 17864
rect 18748 17824 18754 17836
rect 12676 17768 15194 17796
rect 16776 17768 18000 17796
rect 12676 17756 12682 17768
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 12032 17700 12081 17728
rect 12032 17688 12038 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17697 12219 17731
rect 12161 17691 12219 17697
rect 9325 17632 12112 17660
rect 8497 17604 8525 17632
rect 8478 17552 8484 17604
rect 8536 17552 8542 17604
rect 9125 17595 9183 17601
rect 9125 17561 9137 17595
rect 9171 17592 9183 17595
rect 9490 17592 9496 17604
rect 9171 17564 9496 17592
rect 9171 17561 9183 17564
rect 9125 17555 9183 17561
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 10226 17592 10232 17604
rect 9876 17564 10232 17592
rect 8662 17524 8668 17536
rect 8312 17496 8668 17524
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 9876 17533 9904 17564
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 10686 17552 10692 17604
rect 10744 17592 10750 17604
rect 10744 17564 11192 17592
rect 10744 17552 10750 17564
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11164 17533 11192 17564
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 12084 17601 12112 17632
rect 11517 17595 11575 17601
rect 11517 17592 11529 17595
rect 11296 17564 11529 17592
rect 11296 17552 11302 17564
rect 11517 17561 11529 17564
rect 11563 17561 11575 17595
rect 11517 17555 11575 17561
rect 12069 17595 12127 17601
rect 12069 17561 12081 17595
rect 12115 17561 12127 17595
rect 12069 17555 12127 17561
rect 10965 17527 11023 17533
rect 10965 17524 10977 17527
rect 10928 17496 10977 17524
rect 10928 17484 10934 17496
rect 10965 17493 10977 17496
rect 11011 17493 11023 17527
rect 10965 17487 11023 17493
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11974 17484 11980 17536
rect 12032 17524 12038 17536
rect 12176 17524 12204 17691
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 13538 17728 13544 17740
rect 12492 17700 13544 17728
rect 12492 17688 12498 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 16666 17728 16672 17740
rect 13688 17700 16672 17728
rect 13688 17688 13694 17700
rect 16666 17688 16672 17700
rect 16724 17728 16730 17740
rect 16776 17728 16804 17768
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 19024 17768 19288 17796
rect 19024 17756 19030 17768
rect 16724 17700 16804 17728
rect 17221 17731 17279 17737
rect 16724 17688 16730 17700
rect 17221 17697 17233 17731
rect 17267 17697 17279 17731
rect 17221 17691 17279 17697
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13354 17660 13360 17672
rect 12860 17632 13360 17660
rect 12860 17620 12866 17632
rect 13354 17620 13360 17632
rect 13412 17660 13418 17672
rect 16206 17660 16212 17672
rect 13412 17632 16212 17660
rect 13412 17620 13418 17632
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 17236 17660 17264 17691
rect 17310 17688 17316 17740
rect 17368 17728 17374 17740
rect 17405 17731 17463 17737
rect 17405 17728 17417 17731
rect 17368 17700 17417 17728
rect 17368 17688 17374 17700
rect 17405 17697 17417 17700
rect 17451 17697 17463 17731
rect 17405 17691 17463 17697
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 17552 17700 17601 17728
rect 17552 17688 17558 17700
rect 17589 17697 17601 17700
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 17862 17728 17868 17740
rect 17727 17700 17868 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 17957 17731 18015 17737
rect 17957 17697 17969 17731
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 18141 17731 18199 17737
rect 18141 17697 18153 17731
rect 18187 17728 18199 17731
rect 18874 17728 18880 17740
rect 18187 17700 18880 17728
rect 18187 17697 18199 17700
rect 18141 17691 18199 17697
rect 17972 17660 18000 17691
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 19150 17728 19156 17740
rect 18984 17700 19156 17728
rect 18984 17660 19012 17700
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 19260 17737 19288 17768
rect 19426 17756 19432 17808
rect 19484 17756 19490 17808
rect 19536 17805 19564 17836
rect 19794 17824 19800 17876
rect 19852 17824 19858 17876
rect 21542 17864 21548 17876
rect 19950 17836 21548 17864
rect 19521 17799 19579 17805
rect 19521 17765 19533 17799
rect 19567 17796 19579 17799
rect 19950 17796 19978 17836
rect 21542 17824 21548 17836
rect 21600 17864 21606 17876
rect 23290 17864 23296 17876
rect 21600 17836 23296 17864
rect 21600 17824 21606 17836
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 23953 17867 24011 17873
rect 23953 17864 23965 17867
rect 23532 17836 23965 17864
rect 23532 17824 23538 17836
rect 23953 17833 23965 17836
rect 23999 17833 24011 17867
rect 23953 17827 24011 17833
rect 24121 17867 24179 17873
rect 24121 17833 24133 17867
rect 24167 17833 24179 17867
rect 24121 17827 24179 17833
rect 19567 17768 19978 17796
rect 19567 17765 19579 17768
rect 19521 17759 19579 17765
rect 20162 17756 20168 17808
rect 20220 17796 20226 17808
rect 20220 17768 20760 17796
rect 20220 17756 20226 17768
rect 20732 17740 20760 17768
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 20864 17768 21496 17796
rect 20864 17756 20870 17768
rect 19245 17731 19303 17737
rect 19245 17697 19257 17731
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 19610 17688 19616 17740
rect 19668 17688 19674 17740
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 19852 17700 19901 17728
rect 19852 17688 19858 17700
rect 19889 17697 19901 17700
rect 19935 17697 19947 17731
rect 19889 17691 19947 17697
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20088 17700 20668 17728
rect 17236 17632 17540 17660
rect 17972 17632 18276 17660
rect 17512 17604 17540 17632
rect 18248 17604 18276 17632
rect 18892 17632 19012 17660
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 14056 17564 17448 17592
rect 14056 17552 14062 17564
rect 12032 17496 12204 17524
rect 12032 17484 12038 17496
rect 14090 17484 14096 17536
rect 14148 17524 14154 17536
rect 15194 17524 15200 17536
rect 14148 17496 15200 17524
rect 14148 17484 14154 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 17420 17524 17448 17564
rect 17494 17552 17500 17604
rect 17552 17552 17558 17604
rect 18230 17552 18236 17604
rect 18288 17552 18294 17604
rect 18892 17524 18920 17632
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19996 17660 20024 17691
rect 19484 17632 20024 17660
rect 19484 17620 19490 17632
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 20088 17592 20116 17700
rect 20530 17620 20536 17672
rect 20588 17620 20594 17672
rect 20640 17660 20668 17700
rect 20714 17688 20720 17740
rect 20772 17688 20778 17740
rect 21468 17737 21496 17768
rect 21634 17756 21640 17808
rect 21692 17756 21698 17808
rect 23198 17756 23204 17808
rect 23256 17756 23262 17808
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 23753 17799 23811 17805
rect 23753 17796 23765 17799
rect 23624 17768 23765 17796
rect 23624 17756 23630 17768
rect 23753 17765 23765 17768
rect 23799 17765 23811 17799
rect 23753 17759 23811 17765
rect 21453 17731 21511 17737
rect 21453 17697 21465 17731
rect 21499 17697 21511 17731
rect 21453 17691 21511 17697
rect 21545 17731 21603 17737
rect 21545 17697 21557 17731
rect 21591 17697 21603 17731
rect 21545 17691 21603 17697
rect 20806 17660 20812 17672
rect 20640 17632 20812 17660
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21560 17660 21588 17691
rect 21818 17688 21824 17740
rect 21876 17688 21882 17740
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 23216 17728 23244 17756
rect 21959 17700 23244 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 21048 17632 21588 17660
rect 23968 17660 23996 17827
rect 24136 17796 24164 17827
rect 25038 17824 25044 17876
rect 25096 17864 25102 17876
rect 25133 17867 25191 17873
rect 25133 17864 25145 17867
rect 25096 17836 25145 17864
rect 25096 17824 25102 17836
rect 25133 17833 25145 17836
rect 25179 17833 25191 17867
rect 25133 17827 25191 17833
rect 27062 17824 27068 17876
rect 27120 17864 27126 17876
rect 28074 17864 28080 17876
rect 27120 17836 28080 17864
rect 27120 17824 27126 17836
rect 28074 17824 28080 17836
rect 28132 17864 28138 17876
rect 28132 17836 28672 17864
rect 28132 17824 28138 17836
rect 24213 17799 24271 17805
rect 24213 17796 24225 17799
rect 24136 17768 24225 17796
rect 24213 17765 24225 17768
rect 24259 17765 24271 17799
rect 24213 17759 24271 17765
rect 24397 17799 24455 17805
rect 24397 17765 24409 17799
rect 24443 17796 24455 17799
rect 24673 17799 24731 17805
rect 24673 17796 24685 17799
rect 24443 17768 24685 17796
rect 24443 17765 24455 17768
rect 24397 17759 24455 17765
rect 24673 17765 24685 17768
rect 24719 17765 24731 17799
rect 26050 17796 26056 17808
rect 24673 17759 24731 17765
rect 24872 17768 26056 17796
rect 24872 17740 24900 17768
rect 26050 17756 26056 17768
rect 26108 17756 26114 17808
rect 28442 17796 28448 17808
rect 26436 17768 28448 17796
rect 26436 17740 26464 17768
rect 28442 17756 28448 17768
rect 28500 17796 28506 17808
rect 28537 17799 28595 17805
rect 28537 17796 28549 17799
rect 28500 17768 28549 17796
rect 28500 17756 28506 17768
rect 28537 17765 28549 17768
rect 28583 17765 28595 17799
rect 28644 17796 28672 17836
rect 28902 17824 28908 17876
rect 28960 17824 28966 17876
rect 29914 17824 29920 17876
rect 29972 17824 29978 17876
rect 29089 17799 29147 17805
rect 29089 17796 29101 17799
rect 28644 17768 29101 17796
rect 28537 17759 28595 17765
rect 29089 17765 29101 17768
rect 29135 17765 29147 17799
rect 29089 17759 29147 17765
rect 29178 17756 29184 17808
rect 29236 17796 29242 17808
rect 29273 17799 29331 17805
rect 29273 17796 29285 17799
rect 29236 17768 29285 17796
rect 29236 17756 29242 17768
rect 29273 17765 29285 17768
rect 29319 17765 29331 17799
rect 29273 17759 29331 17765
rect 24486 17688 24492 17740
rect 24544 17688 24550 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 24302 17660 24308 17672
rect 23968 17632 24308 17660
rect 21048 17620 21054 17632
rect 24302 17620 24308 17632
rect 24360 17660 24366 17672
rect 24596 17660 24624 17691
rect 24854 17688 24860 17740
rect 24912 17688 24918 17740
rect 25314 17688 25320 17740
rect 25372 17728 25378 17740
rect 25685 17731 25743 17737
rect 25685 17728 25697 17731
rect 25372 17700 25697 17728
rect 25372 17688 25378 17700
rect 25685 17697 25697 17700
rect 25731 17697 25743 17731
rect 25685 17691 25743 17697
rect 25774 17688 25780 17740
rect 25832 17728 25838 17740
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 25832 17700 25973 17728
rect 25832 17688 25838 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 26418 17688 26424 17740
rect 26476 17688 26482 17740
rect 26510 17688 26516 17740
rect 26568 17688 26574 17740
rect 26602 17688 26608 17740
rect 26660 17728 26666 17740
rect 26660 17700 27108 17728
rect 26660 17688 26666 17700
rect 24360 17632 24624 17660
rect 25133 17663 25191 17669
rect 24360 17620 24366 17632
rect 25133 17629 25145 17663
rect 25179 17660 25191 17663
rect 25501 17663 25559 17669
rect 25501 17660 25513 17663
rect 25179 17632 25513 17660
rect 25179 17629 25191 17632
rect 25133 17623 25191 17629
rect 25501 17629 25513 17632
rect 25547 17629 25559 17663
rect 26528 17660 26556 17688
rect 26881 17663 26939 17669
rect 26881 17660 26893 17663
rect 25501 17623 25559 17629
rect 25592 17632 26893 17660
rect 19392 17564 20116 17592
rect 20165 17595 20223 17601
rect 19392 17552 19398 17564
rect 20165 17561 20177 17595
rect 20211 17592 20223 17595
rect 20548 17592 20576 17620
rect 22922 17592 22928 17604
rect 20211 17564 20576 17592
rect 20640 17564 22928 17592
rect 20211 17561 20223 17564
rect 20165 17555 20223 17561
rect 17420 17496 18920 17524
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 20640 17524 20668 17564
rect 22922 17552 22928 17564
rect 22980 17552 22986 17604
rect 24213 17595 24271 17601
rect 24213 17561 24225 17595
rect 24259 17592 24271 17595
rect 24949 17595 25007 17601
rect 24949 17592 24961 17595
rect 24259 17564 24961 17592
rect 24259 17561 24271 17564
rect 24213 17555 24271 17561
rect 24949 17561 24961 17564
rect 24995 17561 25007 17595
rect 24949 17555 25007 17561
rect 19208 17496 20668 17524
rect 19208 17484 19214 17496
rect 21266 17484 21272 17536
rect 21324 17484 21330 17536
rect 22278 17484 22284 17536
rect 22336 17524 22342 17536
rect 23934 17524 23940 17536
rect 22336 17496 23940 17524
rect 22336 17484 22342 17496
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 25592 17524 25620 17632
rect 26881 17629 26893 17632
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 25774 17552 25780 17604
rect 25832 17552 25838 17604
rect 25869 17595 25927 17601
rect 25869 17561 25881 17595
rect 25915 17592 25927 17595
rect 26421 17595 26479 17601
rect 26421 17592 26433 17595
rect 25915 17564 26433 17592
rect 25915 17561 25927 17564
rect 25869 17555 25927 17561
rect 26421 17561 26433 17564
rect 26467 17561 26479 17595
rect 27080 17592 27108 17700
rect 28350 17688 28356 17740
rect 28408 17688 28414 17740
rect 28629 17731 28687 17737
rect 28629 17728 28641 17731
rect 28552 17700 28641 17728
rect 28552 17672 28580 17700
rect 28629 17697 28641 17700
rect 28675 17697 28687 17731
rect 28629 17691 28687 17697
rect 28718 17688 28724 17740
rect 28776 17688 28782 17740
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17697 29055 17731
rect 28997 17691 29055 17697
rect 28534 17620 28540 17672
rect 28592 17620 28598 17672
rect 28626 17592 28632 17604
rect 27080 17564 28632 17592
rect 26421 17555 26479 17561
rect 28626 17552 28632 17564
rect 28684 17552 28690 17604
rect 24912 17496 25620 17524
rect 24912 17484 24918 17496
rect 26510 17484 26516 17536
rect 26568 17524 26574 17536
rect 26789 17527 26847 17533
rect 26789 17524 26801 17527
rect 26568 17496 26801 17524
rect 26568 17484 26574 17496
rect 26789 17493 26801 17496
rect 26835 17524 26847 17527
rect 26970 17524 26976 17536
rect 26835 17496 26976 17524
rect 26835 17493 26847 17496
rect 26789 17487 26847 17493
rect 26970 17484 26976 17496
rect 27028 17484 27034 17536
rect 29012 17524 29040 17691
rect 30190 17688 30196 17740
rect 30248 17688 30254 17740
rect 30285 17731 30343 17737
rect 30285 17697 30297 17731
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 30377 17731 30435 17737
rect 30377 17697 30389 17731
rect 30423 17697 30435 17731
rect 30377 17691 30435 17697
rect 30300 17660 30328 17691
rect 29288 17632 30328 17660
rect 29288 17601 29316 17632
rect 29273 17595 29331 17601
rect 29273 17561 29285 17595
rect 29319 17561 29331 17595
rect 29273 17555 29331 17561
rect 30282 17552 30288 17604
rect 30340 17592 30346 17604
rect 30392 17592 30420 17691
rect 30466 17688 30472 17740
rect 30524 17728 30530 17740
rect 30561 17731 30619 17737
rect 30561 17728 30573 17731
rect 30524 17700 30573 17728
rect 30524 17688 30530 17700
rect 30561 17697 30573 17700
rect 30607 17697 30619 17731
rect 30561 17691 30619 17697
rect 30340 17564 30420 17592
rect 30340 17552 30346 17564
rect 29454 17524 29460 17536
rect 29012 17496 29460 17524
rect 29454 17484 29460 17496
rect 29512 17484 29518 17536
rect 552 17434 31648 17456
rect 552 17382 4285 17434
rect 4337 17382 4349 17434
rect 4401 17382 4413 17434
rect 4465 17382 4477 17434
rect 4529 17382 4541 17434
rect 4593 17382 12059 17434
rect 12111 17382 12123 17434
rect 12175 17382 12187 17434
rect 12239 17382 12251 17434
rect 12303 17382 12315 17434
rect 12367 17382 19833 17434
rect 19885 17382 19897 17434
rect 19949 17382 19961 17434
rect 20013 17382 20025 17434
rect 20077 17382 20089 17434
rect 20141 17382 27607 17434
rect 27659 17382 27671 17434
rect 27723 17382 27735 17434
rect 27787 17382 27799 17434
rect 27851 17382 27863 17434
rect 27915 17382 31648 17434
rect 552 17360 31648 17382
rect 1118 17280 1124 17332
rect 1176 17320 1182 17332
rect 1213 17323 1271 17329
rect 1213 17320 1225 17323
rect 1176 17292 1225 17320
rect 1176 17280 1182 17292
rect 1213 17289 1225 17292
rect 1259 17289 1271 17323
rect 1213 17283 1271 17289
rect 2958 17280 2964 17332
rect 3016 17320 3022 17332
rect 3237 17323 3295 17329
rect 3237 17320 3249 17323
rect 3016 17292 3249 17320
rect 3016 17280 3022 17292
rect 3237 17289 3249 17292
rect 3283 17289 3295 17323
rect 3237 17283 3295 17289
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 3476 17292 4905 17320
rect 3476 17280 3482 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 5353 17323 5411 17329
rect 5353 17289 5365 17323
rect 5399 17320 5411 17323
rect 5626 17320 5632 17332
rect 5399 17292 5632 17320
rect 5399 17289 5411 17292
rect 5353 17283 5411 17289
rect 2866 17212 2872 17264
rect 2924 17252 2930 17264
rect 4706 17252 4712 17264
rect 2924 17224 4712 17252
rect 2924 17212 2930 17224
rect 4706 17212 4712 17224
rect 4764 17212 4770 17264
rect 2130 17144 2136 17196
rect 2188 17144 2194 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 4062 17184 4068 17196
rect 2547 17156 4068 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 5368 17184 5396 17283
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5800 17323 5858 17329
rect 5800 17289 5812 17323
rect 5846 17320 5858 17323
rect 5902 17320 5908 17332
rect 5846 17292 5908 17320
rect 5846 17289 5858 17292
rect 5800 17283 5858 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 8110 17280 8116 17332
rect 8168 17280 8174 17332
rect 8202 17280 8208 17332
rect 8260 17280 8266 17332
rect 8754 17280 8760 17332
rect 8812 17280 8818 17332
rect 8849 17323 8907 17329
rect 8849 17289 8861 17323
rect 8895 17320 8907 17323
rect 8938 17320 8944 17332
rect 8895 17292 8944 17320
rect 8895 17289 8907 17292
rect 8849 17283 8907 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9674 17280 9680 17332
rect 9732 17280 9738 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10410 17320 10416 17332
rect 10192 17292 10416 17320
rect 10192 17280 10198 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 11238 17320 11244 17332
rect 11112 17292 11244 17320
rect 11112 17280 11118 17292
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 13964 17292 14381 17320
rect 13964 17280 13970 17292
rect 14369 17289 14381 17292
rect 14415 17289 14427 17323
rect 14369 17283 14427 17289
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15470 17320 15476 17332
rect 14792 17292 15476 17320
rect 14792 17280 14798 17292
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 16117 17323 16175 17329
rect 16117 17320 16129 17323
rect 15896 17292 16129 17320
rect 15896 17280 15902 17292
rect 16117 17289 16129 17292
rect 16163 17289 16175 17323
rect 16117 17283 16175 17289
rect 16942 17280 16948 17332
rect 17000 17320 17006 17332
rect 17037 17323 17095 17329
rect 17037 17320 17049 17323
rect 17000 17292 17049 17320
rect 17000 17280 17006 17292
rect 17037 17289 17049 17292
rect 17083 17289 17095 17323
rect 17037 17283 17095 17289
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 17862 17320 17868 17332
rect 17736 17292 17868 17320
rect 17736 17280 17742 17292
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 18380 17292 19073 17320
rect 18380 17280 18386 17292
rect 19061 17289 19073 17292
rect 19107 17289 19119 17323
rect 19061 17283 19119 17289
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19886 17320 19892 17332
rect 19300 17292 19892 17320
rect 19300 17280 19306 17292
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 20901 17323 20959 17329
rect 20901 17289 20913 17323
rect 20947 17320 20959 17323
rect 20990 17320 20996 17332
rect 20947 17292 20996 17320
rect 20947 17289 20959 17292
rect 20901 17283 20959 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 21100 17292 23796 17320
rect 6178 17184 6184 17196
rect 4724 17156 5396 17184
rect 5552 17156 6184 17184
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2685 17119 2743 17125
rect 1443 17088 1532 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1504 16989 1532 17088
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 2866 17116 2872 17128
rect 2731 17088 2872 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 3068 17088 3433 17116
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 2958 17048 2964 17060
rect 1903 17020 2964 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 1489 16983 1547 16989
rect 1489 16949 1501 16983
rect 1535 16949 1547 16983
rect 1489 16943 1547 16949
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 2498 16980 2504 16992
rect 1995 16952 2504 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 2498 16940 2504 16952
rect 2556 16980 2562 16992
rect 3068 16989 3096 17088
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 3421 17079 3479 17085
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4724 17125 4752 17156
rect 4341 17119 4399 17125
rect 4341 17116 4353 17119
rect 4212 17088 4353 17116
rect 4212 17076 4218 17088
rect 4341 17085 4353 17088
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 5074 17076 5080 17128
rect 5132 17076 5138 17128
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5552 17125 5580 17156
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7650 17184 7656 17196
rect 7607 17156 7656 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5224 17088 5549 17116
rect 5224 17076 5230 17088
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 6914 17076 6920 17128
rect 6972 17076 6978 17128
rect 7926 17116 7932 17128
rect 7116 17088 7932 17116
rect 3973 17051 4031 17057
rect 3973 17048 3985 17051
rect 3620 17020 3985 17048
rect 3620 16992 3648 17020
rect 3973 17017 3985 17020
rect 4019 17017 4031 17051
rect 3973 17011 4031 17017
rect 4522 17008 4528 17060
rect 4580 17008 4586 17060
rect 4617 17051 4675 17057
rect 4617 17017 4629 17051
rect 4663 17017 4675 17051
rect 4617 17011 4675 17017
rect 2593 16983 2651 16989
rect 2593 16980 2605 16983
rect 2556 16952 2605 16980
rect 2556 16940 2562 16952
rect 2593 16949 2605 16952
rect 2639 16949 2651 16983
rect 2593 16943 2651 16949
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16949 3111 16983
rect 3053 16943 3111 16949
rect 3510 16940 3516 16992
rect 3568 16940 3574 16992
rect 3602 16940 3608 16992
rect 3660 16940 3666 16992
rect 3878 16940 3884 16992
rect 3936 16940 3942 16992
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4632 16980 4660 17011
rect 4212 16952 4660 16980
rect 4212 16940 4218 16952
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 7116 16980 7144 17088
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 7653 17051 7711 17057
rect 7653 17017 7665 17051
rect 7699 17048 7711 17051
rect 7699 17020 7880 17048
rect 7699 17017 7711 17020
rect 7653 17011 7711 17017
rect 7852 16992 7880 17020
rect 5684 16952 7144 16980
rect 7285 16983 7343 16989
rect 5684 16940 5690 16952
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7742 16980 7748 16992
rect 7331 16952 7748 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 7834 16940 7840 16992
rect 7892 16940 7898 16992
rect 8220 16980 8248 17280
rect 9858 17252 9864 17264
rect 9232 17224 9864 17252
rect 9232 17193 9260 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 10226 17212 10232 17264
rect 10284 17212 10290 17264
rect 11790 17252 11796 17264
rect 11348 17224 11796 17252
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9766 17184 9772 17196
rect 9217 17147 9275 17153
rect 9600 17156 9772 17184
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 8352 17088 8401 17116
rect 8352 17076 8358 17088
rect 8389 17085 8401 17088
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17116 9091 17119
rect 9122 17116 9128 17128
rect 9079 17088 9128 17116
rect 9079 17085 9091 17088
rect 9033 17079 9091 17085
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 8570 17008 8576 17060
rect 8628 17048 8634 17060
rect 8754 17048 8760 17060
rect 8628 17020 8760 17048
rect 8628 17008 8634 17020
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 9324 17048 9352 17079
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 9600 17125 9628 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10244 17184 10272 17212
rect 10505 17187 10563 17193
rect 10244 17156 10456 17184
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 9766 17048 9772 17060
rect 9324 17020 9772 17048
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 9876 17048 9904 17079
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10045 17119 10103 17125
rect 10045 17116 10057 17119
rect 10008 17088 10057 17116
rect 10008 17076 10014 17088
rect 10045 17085 10057 17088
rect 10091 17085 10103 17119
rect 10045 17079 10103 17085
rect 10134 17076 10140 17128
rect 10192 17076 10198 17128
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 10318 17076 10324 17128
rect 10376 17076 10382 17128
rect 10428 17125 10456 17156
rect 10505 17153 10517 17187
rect 10551 17184 10563 17187
rect 10686 17184 10692 17196
rect 10551 17156 10692 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 11348 17184 11376 17224
rect 11790 17212 11796 17224
rect 11848 17212 11854 17264
rect 12526 17252 12532 17264
rect 12176 17224 12532 17252
rect 11020 17156 11376 17184
rect 11020 17144 11026 17156
rect 11348 17125 11376 17156
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17085 10471 17119
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10413 17079 10471 17085
rect 10617 17088 11161 17116
rect 10336 17048 10364 17076
rect 10617 17048 10645 17088
rect 11149 17085 11161 17088
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 11333 17079 11391 17085
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 11572 17088 11713 17116
rect 11572 17076 11578 17088
rect 11701 17085 11713 17088
rect 11747 17116 11759 17119
rect 11790 17116 11796 17128
rect 11747 17088 11796 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12176 17125 12204 17224
rect 12526 17212 12532 17224
rect 12584 17252 12590 17264
rect 20622 17252 20628 17264
rect 12584 17224 20628 17252
rect 12584 17212 12590 17224
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 21100 17252 21128 17292
rect 23768 17264 23796 17292
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24670 17320 24676 17332
rect 24176 17292 24676 17320
rect 24176 17280 24182 17292
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 27065 17323 27123 17329
rect 25516 17292 26786 17320
rect 25516 17264 25544 17292
rect 20916 17224 21128 17252
rect 13630 17184 13636 17196
rect 13004 17156 13636 17184
rect 12161 17119 12219 17125
rect 12161 17085 12173 17119
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12526 17116 12532 17128
rect 12483 17088 12532 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17116 12771 17119
rect 13004 17116 13032 17156
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 13906 17184 13912 17196
rect 13833 17156 13912 17184
rect 12759 17088 13032 17116
rect 12759 17085 12771 17088
rect 12713 17079 12771 17085
rect 13078 17076 13084 17128
rect 13136 17076 13142 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13833 17125 13861 17156
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14016 17156 14473 17184
rect 14016 17125 14044 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 16298 17184 16304 17196
rect 14461 17147 14519 17153
rect 15488 17156 16304 17184
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13228 17088 13737 17116
rect 13228 17076 13234 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 13818 17119 13876 17125
rect 13818 17085 13830 17119
rect 13864 17085 13876 17119
rect 13818 17079 13876 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14231 17119 14289 17125
rect 14231 17085 14243 17119
rect 14277 17116 14289 17119
rect 14550 17116 14556 17128
rect 14277 17088 14556 17116
rect 14277 17085 14289 17088
rect 14231 17079 14289 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 14642 17076 14648 17128
rect 14700 17076 14706 17128
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 15194 17116 15200 17128
rect 14967 17088 15200 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 15286 17076 15292 17128
rect 15344 17076 15350 17128
rect 15488 17125 15516 17156
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 18785 17192 18843 17193
rect 18616 17187 18843 17192
rect 18616 17184 18797 17187
rect 17460 17164 18797 17184
rect 17460 17156 18644 17164
rect 17460 17144 17466 17156
rect 18785 17153 18797 17164
rect 18831 17153 18843 17187
rect 18785 17147 18843 17153
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 20254 17184 20260 17196
rect 19760 17156 20260 17184
rect 19760 17144 19766 17156
rect 20254 17144 20260 17156
rect 20312 17184 20318 17196
rect 20312 17156 20760 17184
rect 20312 17144 20318 17156
rect 18693 17129 18751 17135
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17085 15531 17119
rect 15636 17119 15694 17125
rect 15636 17116 15648 17119
rect 15473 17079 15531 17085
rect 15579 17088 15648 17116
rect 9876 17020 10645 17048
rect 10689 17051 10747 17057
rect 10689 17017 10701 17051
rect 10735 17017 10747 17051
rect 10689 17011 10747 17017
rect 10704 16980 10732 17011
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 10836 17020 10885 17048
rect 10836 17008 10842 17020
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 10873 17011 10931 17017
rect 10962 17008 10968 17060
rect 11020 17008 11026 17060
rect 11974 17008 11980 17060
rect 12032 17008 12038 17060
rect 12802 17008 12808 17060
rect 12860 17008 12866 17060
rect 12897 17051 12955 17057
rect 12897 17017 12909 17051
rect 12943 17048 12955 17051
rect 14093 17051 14151 17057
rect 12943 17020 13308 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 11054 16980 11060 16992
rect 8220 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 11480 16952 11529 16980
rect 11480 16940 11486 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 11517 16943 11575 16949
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12158 16980 12164 16992
rect 11664 16952 12164 16980
rect 11664 16940 11670 16952
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 12529 16983 12587 16989
rect 12529 16980 12541 16983
rect 12391 16952 12541 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 12529 16949 12541 16952
rect 12575 16949 12587 16983
rect 12529 16943 12587 16949
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13170 16980 13176 16992
rect 12768 16952 13176 16980
rect 12768 16940 12774 16952
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 13280 16980 13308 17020
rect 14093 17017 14105 17051
rect 14139 17048 14151 17051
rect 15010 17048 15016 17060
rect 14139 17020 15016 17048
rect 14139 17017 14151 17020
rect 14093 17011 14151 17017
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 15304 17048 15332 17076
rect 15579 17048 15607 17088
rect 15636 17085 15648 17088
rect 15682 17085 15694 17119
rect 15636 17079 15694 17085
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 15887 17119 15945 17125
rect 15804 17088 15849 17116
rect 15804 17076 15810 17088
rect 15887 17085 15899 17119
rect 15933 17116 15945 17119
rect 16390 17116 16396 17128
rect 15933 17088 16396 17116
rect 15933 17085 15945 17088
rect 15887 17079 15945 17085
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17184 17088 17233 17116
rect 17184 17076 17190 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17497 17119 17555 17125
rect 17359 17088 17448 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17420 17060 17448 17088
rect 17497 17085 17509 17119
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 15304 17020 15607 17048
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 16540 17020 17356 17048
rect 16540 17008 16546 17020
rect 13446 16980 13452 16992
rect 13280 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16980 13510 16992
rect 14829 16983 14887 16989
rect 14829 16980 14841 16983
rect 13504 16952 14841 16980
rect 13504 16940 13510 16952
rect 14829 16949 14841 16952
rect 14875 16980 14887 16983
rect 17218 16980 17224 16992
rect 14875 16952 17224 16980
rect 14875 16949 14887 16952
rect 14829 16943 14887 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17328 16980 17356 17020
rect 17402 17008 17408 17060
rect 17460 17008 17466 17060
rect 17512 16980 17540 17079
rect 17954 17076 17960 17128
rect 18012 17076 18018 17128
rect 18046 17076 18052 17128
rect 18104 17076 18110 17128
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18279 17088 18368 17116
rect 18693 17095 18705 17129
rect 18739 17095 18751 17129
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18693 17089 18751 17095
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 17972 17048 18000 17076
rect 17972 17020 18092 17048
rect 17954 16980 17960 16992
rect 17328 16952 17960 16980
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18064 16989 18092 17020
rect 18049 16983 18107 16989
rect 18049 16949 18061 16983
rect 18095 16949 18107 16983
rect 18340 16980 18368 17088
rect 18708 17060 18736 17089
rect 18800 17088 18889 17116
rect 18800 17060 18828 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19116 17088 19380 17116
rect 19116 17076 19122 17088
rect 18690 17008 18696 17060
rect 18748 17008 18754 17060
rect 18782 17008 18788 17060
rect 18840 17008 18846 17060
rect 19242 17057 19248 17060
rect 19229 17051 19248 17057
rect 19229 17017 19241 17051
rect 19229 17011 19248 17017
rect 19242 17008 19248 17011
rect 19300 17008 19306 17060
rect 19352 17048 19380 17088
rect 20530 17076 20536 17128
rect 20588 17076 20594 17128
rect 20732 17125 20760 17156
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17085 20775 17119
rect 20717 17079 20775 17085
rect 20806 17076 20812 17128
rect 20864 17076 20870 17128
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 19352 17020 19441 17048
rect 19429 17017 19441 17020
rect 19475 17048 19487 17051
rect 20548 17048 20576 17076
rect 19475 17020 20576 17048
rect 19475 17017 19487 17020
rect 19429 17011 19487 17017
rect 18506 16980 18512 16992
rect 18340 16952 18512 16980
rect 18049 16943 18107 16949
rect 18506 16940 18512 16952
rect 18564 16980 18570 16992
rect 20916 16980 20944 17224
rect 22278 17212 22284 17264
rect 22336 17212 22342 17264
rect 22370 17212 22376 17264
rect 22428 17252 22434 17264
rect 23474 17252 23480 17264
rect 22428 17224 23480 17252
rect 22428 17212 22434 17224
rect 23474 17212 23480 17224
rect 23532 17212 23538 17264
rect 23750 17212 23756 17264
rect 23808 17212 23814 17264
rect 24210 17212 24216 17264
rect 24268 17252 24274 17264
rect 25314 17252 25320 17264
rect 24268 17224 25320 17252
rect 24268 17212 24274 17224
rect 25314 17212 25320 17224
rect 25372 17212 25378 17264
rect 25498 17212 25504 17264
rect 25556 17212 25562 17264
rect 26758 17252 26786 17292
rect 27065 17289 27077 17323
rect 27111 17320 27123 17323
rect 27154 17320 27160 17332
rect 27111 17292 27160 17320
rect 27111 17289 27123 17292
rect 27065 17283 27123 17289
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 27801 17323 27859 17329
rect 27801 17289 27813 17323
rect 27847 17320 27859 17323
rect 27982 17320 27988 17332
rect 27847 17292 27988 17320
rect 27847 17289 27859 17292
rect 27801 17283 27859 17289
rect 27982 17280 27988 17292
rect 28040 17280 28046 17332
rect 30650 17280 30656 17332
rect 30708 17320 30714 17332
rect 30745 17323 30803 17329
rect 30745 17320 30757 17323
rect 30708 17292 30757 17320
rect 30708 17280 30714 17292
rect 30745 17289 30757 17292
rect 30791 17289 30803 17323
rect 30745 17283 30803 17289
rect 28258 17252 28264 17264
rect 26758 17224 28264 17252
rect 28258 17212 28264 17224
rect 28316 17252 28322 17264
rect 29178 17252 29184 17264
rect 28316 17224 29184 17252
rect 28316 17212 28322 17224
rect 29178 17212 29184 17224
rect 29236 17212 29242 17264
rect 30834 17252 30840 17264
rect 30392 17224 30840 17252
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17184 21051 17187
rect 23566 17184 23572 17196
rect 21039 17156 21588 17184
rect 21039 17153 21051 17156
rect 20993 17147 21051 17153
rect 21082 17008 21088 17060
rect 21140 17008 21146 17060
rect 21266 17008 21272 17060
rect 21324 17008 21330 17060
rect 21560 17048 21588 17156
rect 22112 17156 23572 17184
rect 21637 17119 21695 17125
rect 21637 17085 21649 17119
rect 21683 17116 21695 17119
rect 22002 17116 22008 17128
rect 21683 17088 22008 17116
rect 21683 17085 21695 17088
rect 21637 17079 21695 17085
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 22112 17125 22140 17156
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 26234 17184 26240 17196
rect 23992 17156 26240 17184
rect 23992 17144 23998 17156
rect 26234 17144 26240 17156
rect 26292 17184 26298 17196
rect 26602 17184 26608 17196
rect 26292 17156 26608 17184
rect 26292 17144 26298 17156
rect 26602 17144 26608 17156
rect 26660 17184 26666 17196
rect 26660 17156 26740 17184
rect 26660 17144 26666 17156
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17085 22155 17119
rect 22097 17079 22155 17085
rect 22189 17119 22247 17125
rect 22189 17085 22201 17119
rect 22235 17116 22247 17119
rect 22278 17116 22284 17128
rect 22235 17088 22284 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 22373 17119 22431 17125
rect 22373 17085 22385 17119
rect 22419 17085 22431 17119
rect 22373 17079 22431 17085
rect 22388 17048 22416 17079
rect 22922 17076 22928 17128
rect 22980 17076 22986 17128
rect 26712 17125 26740 17156
rect 26970 17144 26976 17196
rect 27028 17184 27034 17196
rect 27183 17184 27384 17192
rect 28626 17184 28632 17196
rect 27028 17164 27936 17184
rect 27028 17156 27211 17164
rect 27356 17156 27936 17164
rect 27028 17144 27034 17156
rect 27249 17129 27307 17135
rect 26422 17119 26480 17125
rect 26422 17116 26434 17119
rect 23032 17088 26434 17116
rect 22940 17048 22968 17076
rect 21560 17020 21956 17048
rect 22388 17020 22968 17048
rect 18564 16952 20944 16980
rect 18564 16940 18570 16952
rect 21358 16940 21364 16992
rect 21416 16940 21422 16992
rect 21453 16983 21511 16989
rect 21453 16949 21465 16983
rect 21499 16980 21511 16983
rect 21634 16980 21640 16992
rect 21499 16952 21640 16980
rect 21499 16949 21511 16952
rect 21453 16943 21511 16949
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 21928 16989 21956 17020
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 23032 16980 23060 17088
rect 26422 17085 26434 17088
rect 26468 17085 26480 17119
rect 26422 17079 26480 17085
rect 26513 17119 26571 17125
rect 26513 17085 26525 17119
rect 26559 17085 26571 17119
rect 26513 17079 26571 17085
rect 26697 17119 26755 17125
rect 26697 17085 26709 17119
rect 26743 17085 26755 17119
rect 26697 17079 26755 17085
rect 23750 17008 23756 17060
rect 23808 17048 23814 17060
rect 25133 17051 25191 17057
rect 25133 17048 25145 17051
rect 23808 17020 25145 17048
rect 23808 17008 23814 17020
rect 25133 17017 25145 17020
rect 25179 17048 25191 17051
rect 26528 17048 26556 17079
rect 26878 17076 26884 17128
rect 26936 17116 26942 17128
rect 27062 17116 27068 17128
rect 26936 17088 27068 17116
rect 26936 17076 26942 17088
rect 27062 17076 27068 17088
rect 27120 17076 27126 17128
rect 27249 17095 27261 17129
rect 27295 17095 27307 17129
rect 27249 17089 27307 17095
rect 27341 17119 27399 17125
rect 27264 17060 27292 17089
rect 27341 17085 27353 17119
rect 27387 17085 27399 17119
rect 27341 17079 27399 17085
rect 25179 17020 26556 17048
rect 26789 17051 26847 17057
rect 25179 17017 25191 17020
rect 25133 17011 25191 17017
rect 26436 16992 26464 17020
rect 26789 17017 26801 17051
rect 26835 17048 26847 17051
rect 26970 17048 26976 17060
rect 26835 17020 26976 17048
rect 26835 17017 26847 17020
rect 26789 17011 26847 17017
rect 26970 17008 26976 17020
rect 27028 17048 27034 17060
rect 27154 17048 27160 17060
rect 27028 17020 27160 17048
rect 27028 17008 27034 17020
rect 27154 17008 27160 17020
rect 27212 17008 27218 17060
rect 27246 17008 27252 17060
rect 27304 17008 27310 17060
rect 27356 17048 27384 17079
rect 27430 17076 27436 17128
rect 27488 17116 27494 17128
rect 27525 17119 27583 17125
rect 27525 17116 27537 17119
rect 27488 17088 27537 17116
rect 27488 17076 27494 17088
rect 27525 17085 27537 17088
rect 27571 17085 27583 17119
rect 27525 17079 27583 17085
rect 27614 17076 27620 17128
rect 27672 17076 27678 17128
rect 27908 17125 27936 17156
rect 28092 17156 28632 17184
rect 28092 17125 28120 17156
rect 28626 17144 28632 17156
rect 28684 17144 28690 17196
rect 28902 17144 28908 17196
rect 28960 17184 28966 17196
rect 29086 17184 29092 17196
rect 28960 17156 29092 17184
rect 28960 17144 28966 17156
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 27893 17119 27951 17125
rect 27893 17085 27905 17119
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17085 28135 17119
rect 28077 17079 28135 17085
rect 29362 17076 29368 17128
rect 29420 17116 29426 17128
rect 30101 17119 30159 17125
rect 30101 17116 30113 17119
rect 29420 17088 30113 17116
rect 29420 17076 29426 17088
rect 30101 17085 30113 17088
rect 30147 17085 30159 17119
rect 30101 17079 30159 17085
rect 30194 17119 30252 17125
rect 30194 17085 30206 17119
rect 30240 17116 30252 17119
rect 30392 17116 30420 17224
rect 30834 17212 30840 17224
rect 30892 17212 30898 17264
rect 30466 17144 30472 17196
rect 30524 17144 30530 17196
rect 30240 17088 30420 17116
rect 30484 17116 30512 17144
rect 30566 17119 30624 17125
rect 30566 17116 30578 17119
rect 30484 17088 30578 17116
rect 30240 17085 30252 17088
rect 30194 17079 30252 17085
rect 30566 17085 30578 17088
rect 30612 17085 30624 17119
rect 30566 17079 30624 17085
rect 27985 17051 28043 17057
rect 27985 17048 27997 17051
rect 27356 17020 27997 17048
rect 27985 17017 27997 17020
rect 28031 17017 28043 17051
rect 27985 17011 28043 17017
rect 28350 17008 28356 17060
rect 28408 17048 28414 17060
rect 30208 17048 30236 17079
rect 28408 17020 30236 17048
rect 28408 17008 28414 17020
rect 30374 17008 30380 17060
rect 30432 17008 30438 17060
rect 30469 17051 30527 17057
rect 30469 17017 30481 17051
rect 30515 17017 30527 17051
rect 30469 17011 30527 17017
rect 21959 16952 23060 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 25314 16980 25320 16992
rect 23164 16952 25320 16980
rect 23164 16940 23170 16952
rect 25314 16940 25320 16952
rect 25372 16940 25378 16992
rect 26418 16940 26424 16992
rect 26476 16940 26482 16992
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 30190 16980 30196 16992
rect 27120 16952 30196 16980
rect 27120 16940 27126 16952
rect 30190 16940 30196 16952
rect 30248 16940 30254 16992
rect 30484 16980 30512 17011
rect 30558 16980 30564 16992
rect 30484 16952 30564 16980
rect 30558 16940 30564 16952
rect 30616 16940 30622 16992
rect 552 16890 31808 16912
rect 552 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 15946 16890
rect 15998 16838 16010 16890
rect 16062 16838 16074 16890
rect 16126 16838 16138 16890
rect 16190 16838 16202 16890
rect 16254 16838 23720 16890
rect 23772 16838 23784 16890
rect 23836 16838 23848 16890
rect 23900 16838 23912 16890
rect 23964 16838 23976 16890
rect 24028 16838 31494 16890
rect 31546 16838 31558 16890
rect 31610 16838 31622 16890
rect 31674 16838 31686 16890
rect 31738 16838 31750 16890
rect 31802 16838 31808 16890
rect 552 16816 31808 16838
rect 3694 16776 3700 16788
rect 860 16748 3700 16776
rect 860 16649 888 16748
rect 845 16643 903 16649
rect 845 16609 857 16643
rect 891 16609 903 16643
rect 2774 16640 2780 16652
rect 2254 16612 2780 16640
rect 845 16603 903 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 3068 16649 3096 16748
rect 3694 16736 3700 16748
rect 3752 16776 3758 16788
rect 5166 16776 5172 16788
rect 3752 16748 5172 16776
rect 3752 16736 3758 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 5815 16748 7665 16776
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 4706 16640 4712 16652
rect 4462 16612 4712 16640
rect 3053 16603 3111 16609
rect 4706 16600 4712 16612
rect 4764 16640 4770 16652
rect 4893 16643 4951 16649
rect 4893 16640 4905 16643
rect 4764 16612 4905 16640
rect 4764 16600 4770 16612
rect 4893 16609 4905 16612
rect 4939 16609 4951 16643
rect 5184 16640 5212 16736
rect 5261 16711 5319 16717
rect 5261 16677 5273 16711
rect 5307 16708 5319 16711
rect 5626 16708 5632 16720
rect 5307 16680 5632 16708
rect 5307 16677 5319 16680
rect 5261 16671 5319 16677
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 5445 16643 5503 16649
rect 5184 16612 5396 16640
rect 4893 16603 4951 16609
rect 1118 16532 1124 16584
rect 1176 16532 1182 16584
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16572 3387 16575
rect 3418 16572 3424 16584
rect 3375 16544 3424 16572
rect 3375 16541 3387 16544
rect 3329 16535 3387 16541
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 5368 16572 5396 16612
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 5815 16640 5843 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8570 16776 8576 16788
rect 7800 16748 8576 16776
rect 7800 16736 7806 16748
rect 8570 16736 8576 16748
rect 8628 16776 8634 16788
rect 9582 16776 9588 16788
rect 8628 16748 9588 16776
rect 8628 16736 8634 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10042 16776 10048 16788
rect 9824 16748 10048 16776
rect 9824 16736 9830 16748
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 7374 16708 7380 16720
rect 7314 16680 7380 16708
rect 7374 16668 7380 16680
rect 7432 16708 7438 16720
rect 10152 16708 10180 16739
rect 10594 16736 10600 16788
rect 10652 16736 10658 16788
rect 11808 16748 13032 16776
rect 7432 16680 9352 16708
rect 7432 16668 7438 16680
rect 7834 16640 7840 16652
rect 5491 16638 5672 16640
rect 5736 16638 5843 16640
rect 5491 16612 5843 16638
rect 7576 16612 7840 16640
rect 5491 16609 5503 16612
rect 5644 16610 5764 16612
rect 5445 16603 5503 16609
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 3844 16544 5304 16572
rect 5368 16544 5825 16572
rect 3844 16532 3850 16544
rect 5276 16516 5304 16544
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5813 16535 5871 16541
rect 5920 16544 6101 16572
rect 5258 16464 5264 16516
rect 5316 16464 5322 16516
rect 5629 16507 5687 16513
rect 5629 16473 5641 16507
rect 5675 16504 5687 16507
rect 5920 16504 5948 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 7098 16532 7104 16584
rect 7156 16532 7162 16584
rect 7576 16581 7604 16612
rect 7834 16600 7840 16612
rect 7892 16640 7898 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 7892 16612 8033 16640
rect 7892 16600 7898 16612
rect 8021 16609 8033 16612
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8159 16612 8340 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 5675 16476 5948 16504
rect 7116 16504 7144 16532
rect 8220 16504 8248 16535
rect 7116 16476 8248 16504
rect 8312 16504 8340 16612
rect 9324 16584 9352 16680
rect 10060 16680 10180 16708
rect 10612 16708 10640 16736
rect 11422 16708 11428 16720
rect 10612 16680 11428 16708
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16642 9919 16643
rect 9950 16642 9956 16652
rect 9907 16614 9956 16642
rect 9907 16609 9919 16614
rect 9861 16603 9919 16609
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8754 16572 8760 16584
rect 8619 16544 8760 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 8938 16532 8944 16584
rect 8996 16532 9002 16584
rect 9306 16532 9312 16584
rect 9364 16532 9370 16584
rect 8956 16504 8984 16532
rect 8312 16476 8984 16504
rect 5675 16473 5687 16476
rect 5629 16467 5687 16473
rect 2590 16396 2596 16448
rect 2648 16436 2654 16448
rect 3786 16436 3792 16448
rect 2648 16408 3792 16436
rect 2648 16396 2654 16408
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4798 16436 4804 16448
rect 3936 16408 4804 16436
rect 3936 16396 3942 16408
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 5166 16396 5172 16448
rect 5224 16436 5230 16448
rect 5350 16436 5356 16448
rect 5224 16408 5356 16436
rect 5224 16396 5230 16408
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9398 16436 9404 16448
rect 9355 16408 9404 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 9508 16436 9536 16603
rect 9950 16600 9956 16614
rect 10008 16600 10014 16652
rect 10060 16649 10088 16680
rect 10318 16649 10324 16652
rect 10045 16643 10103 16649
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 10316 16640 10324 16649
rect 10279 16612 10324 16640
rect 10045 16603 10103 16609
rect 10316 16603 10324 16612
rect 10318 16600 10324 16603
rect 10376 16600 10382 16652
rect 10410 16600 10416 16652
rect 10468 16600 10474 16652
rect 10502 16600 10508 16652
rect 10560 16600 10566 16652
rect 10594 16600 10600 16652
rect 10652 16649 10658 16652
rect 10796 16649 10824 16680
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 10652 16643 10691 16649
rect 10679 16609 10691 16643
rect 10652 16603 10691 16609
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 10652 16600 10658 16603
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 9766 16532 9772 16584
rect 9824 16532 9830 16584
rect 10980 16572 11008 16603
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11808 16649 11836 16748
rect 11882 16668 11888 16720
rect 11940 16668 11946 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 13004 16708 13032 16748
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 13136 16748 14381 16776
rect 13136 16736 13142 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 15562 16776 15568 16788
rect 14516 16748 15568 16776
rect 14516 16736 14522 16748
rect 15562 16736 15568 16748
rect 15620 16776 15626 16788
rect 18414 16776 18420 16788
rect 15620 16748 18420 16776
rect 15620 16736 15626 16748
rect 13906 16708 13912 16720
rect 12216 16680 12388 16708
rect 13004 16680 13912 16708
rect 12216 16668 12222 16680
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11112 16612 11529 16640
rect 11112 16600 11118 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 9968 16544 11008 16572
rect 11716 16572 11744 16603
rect 11900 16572 11928 16668
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 11716 16544 11928 16572
rect 11992 16572 12020 16603
rect 12066 16600 12072 16652
rect 12124 16600 12130 16652
rect 12360 16649 12388 16680
rect 13906 16668 13912 16680
rect 13964 16708 13970 16720
rect 13964 16680 14228 16708
rect 13964 16668 13970 16680
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 12529 16643 12587 16649
rect 12529 16609 12541 16643
rect 12575 16640 12587 16643
rect 13354 16640 13360 16652
rect 12575 16612 13360 16640
rect 12575 16609 12587 16612
rect 12529 16603 12587 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 12618 16572 12624 16584
rect 11992 16544 12624 16572
rect 9968 16504 9996 16544
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16541 12955 16575
rect 12897 16535 12955 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 9789 16476 9996 16504
rect 9789 16436 9817 16476
rect 10226 16464 10232 16516
rect 10284 16504 10290 16516
rect 10962 16504 10968 16516
rect 10284 16476 10968 16504
rect 10284 16464 10290 16476
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 12437 16507 12495 16513
rect 12437 16473 12449 16507
rect 12483 16504 12495 16507
rect 12912 16504 12940 16535
rect 12483 16476 12940 16504
rect 13004 16504 13032 16535
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16572 13231 16575
rect 13219 16544 13400 16572
rect 13219 16541 13231 16544
rect 13173 16535 13231 16541
rect 13372 16516 13400 16544
rect 13004 16476 13308 16504
rect 12483 16473 12495 16476
rect 12437 16467 12495 16473
rect 9508 16408 9817 16436
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 13170 16436 13176 16448
rect 12299 16408 13176 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13280 16436 13308 16476
rect 13354 16464 13360 16516
rect 13412 16464 13418 16516
rect 14108 16504 14136 16603
rect 14200 16572 14228 16680
rect 14292 16680 14780 16708
rect 14292 16649 14320 16680
rect 14752 16652 14780 16680
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14424 16612 14565 16640
rect 14424 16600 14430 16612
rect 14553 16609 14565 16612
rect 14599 16640 14611 16643
rect 14642 16640 14648 16652
rect 14599 16612 14648 16640
rect 14599 16609 14611 16612
rect 14553 16603 14611 16609
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 14734 16600 14740 16652
rect 14792 16600 14798 16652
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 14918 16640 14924 16652
rect 14875 16612 14924 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 16316 16649 16344 16748
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19705 16779 19763 16785
rect 19705 16745 19717 16779
rect 19751 16776 19763 16779
rect 20165 16779 20223 16785
rect 20165 16776 20177 16779
rect 19751 16748 20177 16776
rect 19751 16745 19763 16748
rect 19705 16739 19763 16745
rect 20165 16745 20177 16748
rect 20211 16745 20223 16779
rect 20165 16739 20223 16745
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 21266 16776 21272 16788
rect 20680 16748 21272 16776
rect 20680 16736 20686 16748
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 21692 16748 24624 16776
rect 21692 16736 21698 16748
rect 16574 16668 16580 16720
rect 16632 16668 16638 16720
rect 16684 16680 17632 16708
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16684 16640 16712 16680
rect 16960 16649 16988 16680
rect 16448 16612 16712 16640
rect 16761 16643 16819 16649
rect 16448 16600 16454 16612
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 16117 16575 16175 16581
rect 14200 16544 14964 16572
rect 14936 16516 14964 16544
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16408 16572 16436 16600
rect 16163 16544 16436 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 16776 16572 16804 16603
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 17494 16640 17500 16652
rect 17451 16612 17500 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17604 16640 17632 16680
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 17920 16680 22048 16708
rect 17920 16668 17926 16680
rect 19521 16643 19579 16649
rect 17604 16612 19472 16640
rect 16850 16572 16856 16584
rect 16776 16544 16856 16572
rect 14458 16504 14464 16516
rect 14108 16476 14464 16504
rect 14458 16464 14464 16476
rect 14516 16464 14522 16516
rect 14645 16507 14703 16513
rect 14645 16473 14657 16507
rect 14691 16473 14703 16507
rect 14645 16467 14703 16473
rect 14090 16436 14096 16448
rect 13280 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 14366 16436 14372 16448
rect 14323 16408 14372 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14660 16436 14688 16467
rect 14734 16464 14740 16516
rect 14792 16464 14798 16516
rect 14918 16464 14924 16516
rect 14976 16464 14982 16516
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 16776 16504 16804 16544
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 18598 16572 18604 16584
rect 17420 16544 18604 16572
rect 17420 16504 17448 16544
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 19444 16572 19472 16612
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 19702 16640 19708 16652
rect 19567 16612 19708 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19444 16544 19748 16572
rect 19720 16516 19748 16544
rect 16356 16476 17448 16504
rect 16356 16464 16362 16476
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 19150 16504 19156 16516
rect 18104 16476 19156 16504
rect 18104 16464 18110 16476
rect 19150 16464 19156 16476
rect 19208 16464 19214 16516
rect 19337 16507 19395 16513
rect 19337 16473 19349 16507
rect 19383 16504 19395 16507
rect 19426 16504 19432 16516
rect 19383 16476 19432 16504
rect 19383 16473 19395 16476
rect 19337 16467 19395 16473
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 19822 16504 19850 16603
rect 19886 16600 19892 16652
rect 19944 16600 19950 16652
rect 20088 16649 20116 16680
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16609 20131 16643
rect 20073 16603 20131 16609
rect 20162 16600 20168 16652
rect 20220 16600 20226 16652
rect 20349 16643 20407 16649
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 20530 16640 20536 16652
rect 20395 16612 20536 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21542 16640 21548 16652
rect 20956 16612 21548 16640
rect 20956 16600 20962 16612
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 22020 16649 22048 16680
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 22373 16711 22431 16717
rect 22373 16708 22385 16711
rect 22336 16680 22385 16708
rect 22336 16668 22342 16680
rect 22373 16677 22385 16680
rect 22419 16677 22431 16711
rect 22373 16671 22431 16677
rect 22738 16668 22744 16720
rect 22796 16708 22802 16720
rect 24210 16708 24216 16720
rect 22796 16680 23428 16708
rect 22796 16668 22802 16680
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 23017 16643 23075 16649
rect 23017 16640 23029 16643
rect 22612 16612 23029 16640
rect 22612 16600 22618 16612
rect 23017 16609 23029 16612
rect 23063 16609 23075 16643
rect 23017 16603 23075 16609
rect 23106 16600 23112 16652
rect 23164 16600 23170 16652
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23290 16640 23296 16652
rect 23247 16612 23296 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 23290 16600 23296 16612
rect 23348 16600 23354 16652
rect 23400 16649 23428 16680
rect 23492 16680 24216 16708
rect 23492 16649 23520 16680
rect 24210 16668 24216 16680
rect 24268 16668 24274 16720
rect 24302 16668 24308 16720
rect 24360 16668 24366 16720
rect 24394 16668 24400 16720
rect 24452 16668 24458 16720
rect 23385 16643 23443 16649
rect 23385 16609 23397 16643
rect 23431 16609 23443 16643
rect 23385 16603 23443 16609
rect 23477 16643 23535 16649
rect 23477 16609 23489 16643
rect 23523 16609 23535 16643
rect 24320 16639 24348 16668
rect 24489 16643 24547 16649
rect 23477 16603 23535 16609
rect 24305 16633 24363 16639
rect 24305 16599 24317 16633
rect 24351 16599 24363 16633
rect 24489 16609 24501 16643
rect 24535 16609 24547 16643
rect 24596 16640 24624 16748
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 24728 16748 25329 16776
rect 24728 16736 24734 16748
rect 25317 16745 25329 16748
rect 25363 16745 25375 16779
rect 25317 16739 25375 16745
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 26421 16779 26479 16785
rect 26421 16776 26433 16779
rect 25832 16748 26433 16776
rect 25832 16736 25838 16748
rect 26421 16745 26433 16748
rect 26467 16745 26479 16779
rect 26421 16739 26479 16745
rect 26602 16736 26608 16788
rect 26660 16776 26666 16788
rect 26970 16776 26976 16788
rect 26660 16748 26976 16776
rect 26660 16736 26666 16748
rect 26970 16736 26976 16748
rect 27028 16736 27034 16788
rect 27154 16736 27160 16788
rect 27212 16736 27218 16788
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 28169 16779 28227 16785
rect 28169 16776 28181 16779
rect 27488 16748 28181 16776
rect 27488 16736 27494 16748
rect 28169 16745 28181 16748
rect 28215 16776 28227 16779
rect 30558 16776 30564 16788
rect 28215 16748 30564 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 30558 16736 30564 16748
rect 30616 16736 30622 16788
rect 24949 16711 25007 16717
rect 24949 16677 24961 16711
rect 24995 16708 25007 16711
rect 25038 16708 25044 16720
rect 24995 16680 25044 16708
rect 24995 16677 25007 16680
rect 24949 16671 25007 16677
rect 25038 16668 25044 16680
rect 25096 16708 25102 16720
rect 25133 16711 25191 16717
rect 25133 16708 25145 16711
rect 25096 16680 25145 16708
rect 25096 16668 25102 16680
rect 25133 16677 25145 16680
rect 25179 16677 25191 16711
rect 25133 16671 25191 16677
rect 25222 16668 25228 16720
rect 25280 16708 25286 16720
rect 25685 16711 25743 16717
rect 25280 16680 25544 16708
rect 25280 16668 25286 16680
rect 25516 16640 25544 16680
rect 25685 16677 25697 16711
rect 25731 16708 25743 16711
rect 25731 16680 28212 16708
rect 25731 16677 25743 16680
rect 25685 16671 25743 16677
rect 25961 16643 26019 16649
rect 25961 16640 25973 16643
rect 24596 16612 25452 16640
rect 25516 16612 25973 16640
rect 24489 16603 24547 16609
rect 24305 16593 24363 16599
rect 19978 16532 19984 16584
rect 20036 16532 20042 16584
rect 21358 16532 21364 16584
rect 21416 16572 21422 16584
rect 24504 16572 24532 16603
rect 25424 16572 25452 16612
rect 25961 16609 25973 16612
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26697 16643 26755 16649
rect 26697 16640 26709 16643
rect 26292 16612 26709 16640
rect 26292 16600 26298 16612
rect 26697 16609 26709 16612
rect 26743 16609 26755 16643
rect 26697 16603 26755 16609
rect 26789 16643 26847 16649
rect 26789 16609 26801 16643
rect 26835 16609 26847 16643
rect 26789 16603 26847 16609
rect 25685 16575 25743 16581
rect 25685 16572 25697 16575
rect 21416 16544 24256 16572
rect 21416 16532 21422 16544
rect 20162 16504 20168 16516
rect 19822 16476 20168 16504
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 22922 16504 22928 16516
rect 20772 16476 22928 16504
rect 20772 16464 20778 16476
rect 22922 16464 22928 16476
rect 22980 16464 22986 16516
rect 23566 16464 23572 16516
rect 23624 16464 23630 16516
rect 24228 16504 24256 16544
rect 24504 16544 25360 16572
rect 25424 16544 25697 16572
rect 24504 16504 24532 16544
rect 24228 16476 24532 16504
rect 16758 16436 16764 16448
rect 14660 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 16942 16436 16948 16448
rect 16899 16408 16948 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 16942 16396 16948 16408
rect 17000 16436 17006 16448
rect 17126 16436 17132 16448
rect 17000 16408 17132 16436
rect 17000 16396 17006 16408
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17402 16396 17408 16448
rect 17460 16396 17466 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18598 16436 18604 16448
rect 18012 16408 18604 16436
rect 18012 16396 18018 16408
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 21266 16436 21272 16448
rect 19668 16408 21272 16436
rect 19668 16396 19674 16408
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22373 16439 22431 16445
rect 22373 16436 22385 16439
rect 22244 16408 22385 16436
rect 22244 16396 22250 16408
rect 22373 16405 22385 16408
rect 22419 16405 22431 16439
rect 22373 16399 22431 16405
rect 22557 16439 22615 16445
rect 22557 16405 22569 16439
rect 22603 16436 22615 16439
rect 22738 16436 22744 16448
rect 22603 16408 22744 16436
rect 22603 16405 22615 16408
rect 22557 16399 22615 16405
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 22830 16396 22836 16448
rect 22888 16396 22894 16448
rect 23584 16436 23612 16464
rect 24578 16436 24584 16448
rect 23584 16408 24584 16436
rect 24578 16396 24584 16408
rect 24636 16436 24642 16448
rect 24673 16439 24731 16445
rect 24673 16436 24685 16439
rect 24636 16408 24685 16436
rect 24636 16396 24642 16408
rect 24673 16405 24685 16408
rect 24719 16436 24731 16439
rect 25222 16436 25228 16448
rect 24719 16408 25228 16436
rect 24719 16405 24731 16408
rect 24673 16399 24731 16405
rect 25222 16396 25228 16408
rect 25280 16396 25286 16448
rect 25332 16445 25360 16544
rect 25685 16541 25697 16544
rect 25731 16541 25743 16575
rect 26804 16572 26832 16603
rect 26878 16600 26884 16652
rect 26936 16600 26942 16652
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 27028 16612 27077 16640
rect 27028 16600 27034 16612
rect 27065 16609 27077 16612
rect 27111 16609 27123 16643
rect 27065 16603 27123 16609
rect 27157 16643 27215 16649
rect 27157 16609 27169 16643
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 27183 16572 27211 16603
rect 27246 16600 27252 16652
rect 27304 16640 27310 16652
rect 27341 16643 27399 16649
rect 27341 16640 27353 16643
rect 27304 16612 27353 16640
rect 27304 16600 27310 16612
rect 27341 16609 27353 16612
rect 27387 16609 27399 16643
rect 27341 16603 27399 16609
rect 27985 16643 28043 16649
rect 27985 16609 27997 16643
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 26804 16544 27211 16572
rect 25685 16535 25743 16541
rect 26988 16516 27016 16544
rect 25498 16464 25504 16516
rect 25556 16464 25562 16516
rect 25774 16464 25780 16516
rect 25832 16504 25838 16516
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 25832 16476 25881 16504
rect 25832 16464 25838 16476
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 26970 16464 26976 16516
rect 27028 16464 27034 16516
rect 27154 16464 27160 16516
rect 27212 16504 27218 16516
rect 27614 16504 27620 16516
rect 27212 16476 27620 16504
rect 27212 16464 27218 16476
rect 27614 16464 27620 16476
rect 27672 16464 27678 16516
rect 25317 16439 25375 16445
rect 25317 16405 25329 16439
rect 25363 16436 25375 16439
rect 28000 16436 28028 16603
rect 28184 16572 28212 16680
rect 28276 16680 28856 16708
rect 28276 16652 28304 16680
rect 28258 16600 28264 16652
rect 28316 16600 28322 16652
rect 28534 16600 28540 16652
rect 28592 16640 28598 16652
rect 28828 16649 28856 16680
rect 28920 16680 29316 16708
rect 28629 16643 28687 16649
rect 28629 16640 28641 16643
rect 28592 16612 28641 16640
rect 28592 16600 28598 16612
rect 28629 16609 28641 16612
rect 28675 16609 28687 16643
rect 28629 16603 28687 16609
rect 28813 16643 28871 16649
rect 28813 16609 28825 16643
rect 28859 16609 28871 16643
rect 28813 16603 28871 16609
rect 28920 16572 28948 16680
rect 29089 16643 29147 16649
rect 29089 16609 29101 16643
rect 29135 16609 29147 16643
rect 29089 16603 29147 16609
rect 28184 16544 28948 16572
rect 28810 16464 28816 16516
rect 28868 16464 28874 16516
rect 28902 16464 28908 16516
rect 28960 16464 28966 16516
rect 28350 16436 28356 16448
rect 25363 16408 28356 16436
rect 25363 16405 25375 16408
rect 25317 16399 25375 16405
rect 28350 16396 28356 16408
rect 28408 16396 28414 16448
rect 29104 16436 29132 16603
rect 29178 16600 29184 16652
rect 29236 16600 29242 16652
rect 29288 16649 29316 16680
rect 29273 16643 29331 16649
rect 29273 16609 29285 16643
rect 29319 16609 29331 16643
rect 29273 16603 29331 16609
rect 29362 16600 29368 16652
rect 29420 16600 29426 16652
rect 29546 16600 29552 16652
rect 29604 16600 29610 16652
rect 30374 16600 30380 16652
rect 30432 16640 30438 16652
rect 30650 16640 30656 16652
rect 30432 16612 30656 16640
rect 30432 16600 30438 16612
rect 30650 16600 30656 16612
rect 30708 16600 30714 16652
rect 29196 16513 29224 16600
rect 29181 16507 29239 16513
rect 29181 16473 29193 16507
rect 29227 16473 29239 16507
rect 29181 16467 29239 16473
rect 29270 16436 29276 16448
rect 29104 16408 29276 16436
rect 29270 16396 29276 16408
rect 29328 16396 29334 16448
rect 552 16346 31648 16368
rect 552 16294 4285 16346
rect 4337 16294 4349 16346
rect 4401 16294 4413 16346
rect 4465 16294 4477 16346
rect 4529 16294 4541 16346
rect 4593 16294 12059 16346
rect 12111 16294 12123 16346
rect 12175 16294 12187 16346
rect 12239 16294 12251 16346
rect 12303 16294 12315 16346
rect 12367 16294 19833 16346
rect 19885 16294 19897 16346
rect 19949 16294 19961 16346
rect 20013 16294 20025 16346
rect 20077 16294 20089 16346
rect 20141 16294 27607 16346
rect 27659 16294 27671 16346
rect 27723 16294 27735 16346
rect 27787 16294 27799 16346
rect 27851 16294 27863 16346
rect 27915 16294 31648 16346
rect 552 16272 31648 16294
rect 1118 16192 1124 16244
rect 1176 16232 1182 16244
rect 1213 16235 1271 16241
rect 1213 16232 1225 16235
rect 1176 16204 1225 16232
rect 1176 16192 1182 16204
rect 1213 16201 1225 16204
rect 1259 16201 1271 16235
rect 7561 16235 7619 16241
rect 1213 16195 1271 16201
rect 2424 16204 4200 16232
rect 1026 16124 1032 16176
rect 1084 16164 1090 16176
rect 2317 16167 2375 16173
rect 2317 16164 2329 16167
rect 1084 16136 2329 16164
rect 1084 16124 1090 16136
rect 2317 16133 2329 16136
rect 2363 16133 2375 16167
rect 2317 16127 2375 16133
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 2424 16096 2452 16204
rect 4062 16164 4068 16176
rect 2976 16136 4068 16164
rect 2976 16105 3004 16136
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 2188 16068 2452 16096
rect 2961 16099 3019 16105
rect 2188 16056 2194 16068
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3142 16056 3148 16108
rect 3200 16096 3206 16108
rect 3973 16099 4031 16105
rect 3200 16068 3740 16096
rect 3200 16056 3206 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1857 16031 1915 16037
rect 1443 16000 1532 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1504 15901 1532 16000
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2590 16028 2596 16040
rect 1903 16000 2596 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 2866 16028 2872 16040
rect 2731 16000 2872 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3602 16028 3608 16040
rect 3160 16000 3608 16028
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 3160 15960 3188 16000
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 3712 16037 3740 16068
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4172 16096 4200 16204
rect 4913 16204 7328 16232
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 4019 16068 4353 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 4341 16065 4353 16068
rect 4387 16096 4399 16099
rect 4913 16096 4941 16204
rect 5000 16136 5304 16164
rect 5000 16108 5028 16136
rect 4387 16068 4941 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 4982 16056 4988 16108
rect 5040 16056 5046 16108
rect 5166 16056 5172 16108
rect 5224 16056 5230 16108
rect 5276 16105 5304 16136
rect 7300 16108 7328 16204
rect 7561 16201 7573 16235
rect 7607 16232 7619 16235
rect 8754 16232 8760 16244
rect 7607 16204 8760 16232
rect 7607 16201 7619 16204
rect 7561 16195 7619 16201
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5592 16068 5825 16096
rect 5592 16056 5598 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7742 16096 7748 16108
rect 7340 16068 7748 16096
rect 7340 16056 7346 16068
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 7852 16105 7880 16204
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 8869 16204 9076 16232
rect 8389 16167 8447 16173
rect 8389 16133 8401 16167
rect 8435 16164 8447 16167
rect 8662 16164 8668 16176
rect 8435 16136 8668 16164
rect 8435 16133 8447 16136
rect 8389 16127 8447 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16065 7895 16099
rect 8869 16096 8897 16204
rect 9048 16105 9076 16204
rect 9306 16192 9312 16244
rect 9364 16192 9370 16244
rect 9398 16192 9404 16244
rect 9456 16192 9462 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9858 16232 9864 16244
rect 9732 16204 9864 16232
rect 9732 16192 9738 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10870 16192 10876 16244
rect 10928 16192 10934 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11425 16235 11483 16241
rect 11425 16232 11437 16235
rect 11388 16204 11437 16232
rect 11388 16192 11394 16204
rect 11425 16201 11437 16204
rect 11471 16201 11483 16235
rect 11425 16195 11483 16201
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12253 16235 12311 16241
rect 12253 16232 12265 16235
rect 12032 16204 12265 16232
rect 12032 16192 12038 16204
rect 12253 16201 12265 16204
rect 12299 16201 12311 16235
rect 12253 16195 12311 16201
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 13412 16204 14504 16232
rect 13412 16192 13418 16204
rect 9416 16164 9444 16192
rect 10888 16164 10916 16192
rect 9416 16136 9674 16164
rect 10888 16136 12296 16164
rect 7837 16059 7895 16065
rect 7944 16068 8897 16096
rect 9033 16099 9091 16105
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 5350 16028 5356 16040
rect 3743 16000 5356 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 7374 16028 7380 16040
rect 7222 16000 7380 16028
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 7760 16028 7788 16056
rect 7944 16028 7972 16068
rect 9033 16065 9045 16099
rect 9079 16065 9091 16099
rect 9646 16096 9674 16136
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9646 16068 9873 16096
rect 9033 16059 9091 16065
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11112 16068 11345 16096
rect 11112 16056 11118 16068
rect 11333 16065 11345 16068
rect 11379 16096 11391 16099
rect 11379 16068 11836 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 7760 16000 7972 16028
rect 8018 15988 8024 16040
rect 8076 15988 8082 16040
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8478 16028 8484 16040
rect 8251 16000 8484 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 9306 15988 9312 16040
rect 9364 16038 9370 16040
rect 9364 16028 9444 16038
rect 9582 16028 9588 16040
rect 9364 16010 9588 16028
rect 9364 15988 9370 16010
rect 9416 16000 9588 16010
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 11808 16037 11836 16068
rect 11882 16056 11888 16108
rect 11940 16096 11946 16108
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11940 16068 11989 16096
rect 11940 16056 11946 16068
rect 11977 16065 11989 16068
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12268 16037 12296 16136
rect 12802 16124 12808 16176
rect 12860 16164 12866 16176
rect 13998 16164 14004 16176
rect 12860 16136 14004 16164
rect 12860 16124 12866 16136
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 13044 16068 13093 16096
rect 13044 16056 13050 16068
rect 13081 16065 13093 16068
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13630 16096 13636 16108
rect 13403 16068 13636 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 1995 15932 3188 15960
rect 3252 15932 3801 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 3252 15904 3280 15932
rect 3789 15929 3801 15932
rect 3835 15929 3847 15963
rect 3789 15923 3847 15929
rect 4433 15963 4491 15969
rect 4433 15929 4445 15963
rect 4479 15960 4491 15963
rect 5626 15960 5632 15972
rect 4479 15932 5632 15960
rect 4479 15929 4491 15932
rect 4433 15923 4491 15929
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 6086 15920 6092 15972
rect 6144 15920 6150 15972
rect 8496 15932 9352 15960
rect 1489 15895 1547 15901
rect 1489 15861 1501 15895
rect 1535 15861 1547 15895
rect 1489 15855 1547 15861
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 3234 15892 3240 15904
rect 2823 15864 3240 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 3326 15852 3332 15904
rect 3384 15852 3390 15904
rect 4525 15895 4583 15901
rect 4525 15861 4537 15895
rect 4571 15892 4583 15895
rect 4614 15892 4620 15904
rect 4571 15864 4620 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 4893 15895 4951 15901
rect 4893 15861 4905 15895
rect 4939 15892 4951 15895
rect 5166 15892 5172 15904
rect 4939 15864 5172 15892
rect 4939 15861 4951 15864
rect 4893 15855 4951 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5721 15895 5779 15901
rect 5721 15861 5733 15895
rect 5767 15892 5779 15895
rect 8496 15892 8524 15932
rect 5767 15864 8524 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8628 15864 8769 15892
rect 8628 15852 8634 15864
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 8757 15855 8815 15861
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 8938 15892 8944 15904
rect 8895 15864 8944 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9324 15892 9352 15932
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 9950 15960 9956 15972
rect 9456 15932 9956 15960
rect 9456 15920 9462 15932
rect 9950 15920 9956 15932
rect 10008 15960 10014 15972
rect 11885 15963 11943 15969
rect 11885 15960 11897 15963
rect 10008 15932 10350 15960
rect 11164 15932 11897 15960
rect 10008 15920 10014 15932
rect 11164 15892 11192 15932
rect 11885 15929 11897 15932
rect 11931 15929 11943 15963
rect 11885 15923 11943 15929
rect 9324 15864 11192 15892
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 12452 15892 12480 15991
rect 12872 15963 12930 15969
rect 12872 15929 12884 15963
rect 12918 15960 12930 15963
rect 14366 15960 14372 15972
rect 12918 15932 14372 15960
rect 12918 15929 12930 15932
rect 12872 15923 12930 15929
rect 14366 15920 14372 15932
rect 14424 15920 14430 15972
rect 14476 15960 14504 16204
rect 14550 16192 14556 16244
rect 14608 16232 14614 16244
rect 14645 16235 14703 16241
rect 14645 16232 14657 16235
rect 14608 16204 14657 16232
rect 14608 16192 14614 16204
rect 14645 16201 14657 16204
rect 14691 16201 14703 16235
rect 14645 16195 14703 16201
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 14918 16232 14924 16244
rect 14875 16204 14924 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 17310 16232 17316 16244
rect 16356 16204 17316 16232
rect 16356 16192 16362 16204
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 17911 16204 18920 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 15378 16164 15384 16176
rect 14568 16136 15384 16164
rect 14568 16037 14596 16136
rect 15378 16124 15384 16136
rect 15436 16164 15442 16176
rect 16390 16164 16396 16176
rect 15436 16136 16396 16164
rect 15436 16124 15442 16136
rect 16390 16124 16396 16136
rect 16448 16124 16454 16176
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 17402 16164 17408 16176
rect 16816 16136 17408 16164
rect 16816 16124 16822 16136
rect 17402 16124 17408 16136
rect 17460 16164 17466 16176
rect 17589 16167 17647 16173
rect 17589 16164 17601 16167
rect 17460 16136 17601 16164
rect 17460 16124 17466 16136
rect 17589 16133 17601 16136
rect 17635 16133 17647 16167
rect 17589 16127 17647 16133
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18138 16164 18144 16176
rect 18012 16136 18144 16164
rect 18012 16124 18018 16136
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 18690 16124 18696 16176
rect 18748 16124 18754 16176
rect 15746 16096 15752 16108
rect 14844 16068 15752 16096
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 14844 16037 14872 16068
rect 15746 16056 15752 16068
rect 15804 16096 15810 16108
rect 18708 16096 18736 16124
rect 15804 16068 18736 16096
rect 15804 16056 15810 16068
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15286 16028 15292 16040
rect 15059 16000 15292 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17310 16028 17316 16040
rect 17267 16000 17316 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 17402 15988 17408 16040
rect 17460 15988 17466 16040
rect 17494 15988 17500 16040
rect 17552 15988 17558 16040
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 16028 17739 16031
rect 17770 16028 17776 16040
rect 17727 16000 17776 16028
rect 17727 15997 17739 16000
rect 17681 15991 17739 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18598 16028 18604 16040
rect 18012 16000 18604 16028
rect 18012 15988 18018 16000
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 18892 16037 18920 16204
rect 18966 16192 18972 16244
rect 19024 16192 19030 16244
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 19300 16204 19441 16232
rect 19300 16192 19306 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 21177 16235 21235 16241
rect 21177 16232 21189 16235
rect 20956 16204 21189 16232
rect 20956 16192 20962 16204
rect 21177 16201 21189 16204
rect 21223 16201 21235 16235
rect 21818 16232 21824 16244
rect 21177 16195 21235 16201
rect 21284 16204 21824 16232
rect 18984 16096 19012 16192
rect 19337 16167 19395 16173
rect 19337 16133 19349 16167
rect 19383 16164 19395 16167
rect 21284 16164 21312 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 21910 16192 21916 16244
rect 21968 16232 21974 16244
rect 22925 16235 22983 16241
rect 21968 16204 22692 16232
rect 21968 16192 21974 16204
rect 19383 16136 21312 16164
rect 21637 16167 21695 16173
rect 19383 16133 19395 16136
rect 19337 16127 19395 16133
rect 21637 16133 21649 16167
rect 21683 16164 21695 16167
rect 22664 16164 22692 16204
rect 22925 16201 22937 16235
rect 22971 16232 22983 16235
rect 23014 16232 23020 16244
rect 22971 16204 23020 16232
rect 22971 16201 22983 16204
rect 22925 16195 22983 16201
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 23382 16232 23388 16244
rect 23164 16204 23388 16232
rect 23164 16192 23170 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 24210 16192 24216 16244
rect 24268 16192 24274 16244
rect 24394 16192 24400 16244
rect 24452 16232 24458 16244
rect 25774 16232 25780 16244
rect 24452 16204 25780 16232
rect 24452 16192 24458 16204
rect 25774 16192 25780 16204
rect 25832 16192 25838 16244
rect 26050 16192 26056 16244
rect 26108 16232 26114 16244
rect 29362 16232 29368 16244
rect 26108 16204 29368 16232
rect 26108 16192 26114 16204
rect 29362 16192 29368 16204
rect 29420 16232 29426 16244
rect 29638 16232 29644 16244
rect 29420 16204 29644 16232
rect 29420 16192 29426 16204
rect 29638 16192 29644 16204
rect 29696 16192 29702 16244
rect 30190 16192 30196 16244
rect 30248 16192 30254 16244
rect 30377 16235 30435 16241
rect 30377 16201 30389 16235
rect 30423 16201 30435 16235
rect 30377 16195 30435 16201
rect 24228 16164 24256 16192
rect 21683 16136 22600 16164
rect 22664 16136 24256 16164
rect 21683 16133 21695 16136
rect 21637 16127 21695 16133
rect 19242 16096 19248 16108
rect 18984 16068 19248 16096
rect 19242 16056 19248 16068
rect 19300 16096 19306 16108
rect 19300 16068 19748 16096
rect 19300 16056 19306 16068
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 18877 16031 18935 16037
rect 18877 15997 18889 16031
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 18322 15960 18328 15972
rect 14476 15932 18328 15960
rect 18322 15920 18328 15932
rect 18380 15960 18386 15972
rect 18708 15960 18736 15991
rect 18966 15988 18972 16040
rect 19024 15988 19030 16040
rect 19058 15988 19064 16040
rect 19116 15988 19122 16040
rect 19720 16037 19748 16068
rect 20070 16056 20076 16108
rect 20128 16096 20134 16108
rect 20128 16068 20760 16096
rect 20128 16056 20134 16068
rect 19705 16031 19763 16037
rect 19614 16009 19672 16015
rect 19614 15975 19626 16009
rect 19660 15975 19672 16009
rect 19705 15997 19717 16031
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 16028 19855 16031
rect 20533 16031 20591 16037
rect 19843 16000 20392 16028
rect 19843 15997 19855 16000
rect 19797 15991 19855 15997
rect 19614 15972 19672 15975
rect 19426 15960 19432 15972
rect 18380 15932 18736 15960
rect 18800 15932 19432 15960
rect 18380 15920 18386 15932
rect 11296 15864 12480 15892
rect 11296 15852 11302 15864
rect 12710 15852 12716 15904
rect 12768 15852 12774 15904
rect 12989 15895 13047 15901
rect 12989 15861 13001 15895
rect 13035 15892 13047 15895
rect 13078 15892 13084 15904
rect 13035 15864 13084 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13078 15852 13084 15864
rect 13136 15892 13142 15904
rect 13446 15892 13452 15904
rect 13136 15864 13452 15892
rect 13136 15852 13142 15864
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 18800 15892 18828 15932
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 19610 15920 19616 15972
rect 19668 15920 19674 15972
rect 17644 15864 18828 15892
rect 17644 15852 17650 15864
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19812 15892 19840 15991
rect 20364 15972 20392 16000
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 19935 15963 19993 15969
rect 19935 15929 19947 15963
rect 19981 15960 19993 15963
rect 20162 15960 20168 15972
rect 19981 15932 20168 15960
rect 19981 15929 19993 15932
rect 19935 15923 19993 15929
rect 20162 15920 20168 15932
rect 20220 15920 20226 15972
rect 20346 15920 20352 15972
rect 20404 15920 20410 15972
rect 20548 15960 20576 15991
rect 20622 15988 20628 16040
rect 20680 15988 20686 16040
rect 20732 16028 20760 16068
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 20990 16056 20996 16108
rect 21048 16056 21054 16108
rect 21174 16056 21180 16108
rect 21232 16056 21238 16108
rect 21266 16056 21272 16108
rect 21324 16056 21330 16108
rect 21008 16028 21036 16056
rect 21192 16028 21220 16056
rect 20732 16000 21036 16028
rect 21100 16000 21220 16028
rect 21453 16031 21511 16037
rect 20548 15932 20668 15960
rect 18932 15864 19840 15892
rect 20640 15892 20668 15932
rect 20990 15892 20996 15904
rect 20640 15864 20996 15892
rect 18932 15852 18938 15864
rect 20990 15852 20996 15864
rect 21048 15892 21054 15904
rect 21100 15892 21128 16000
rect 21453 15997 21465 16031
rect 21499 16028 21511 16031
rect 21910 16028 21916 16040
rect 21499 16000 21916 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 22572 16037 22600 16136
rect 27062 16124 27068 16176
rect 27120 16124 27126 16176
rect 28626 16164 28632 16176
rect 27172 16136 28632 16164
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16096 22799 16099
rect 22830 16096 22836 16108
rect 22787 16068 22836 16096
rect 22787 16065 22799 16068
rect 22741 16059 22799 16065
rect 22830 16056 22836 16068
rect 22888 16056 22894 16108
rect 25682 16096 25688 16108
rect 23032 16068 25688 16096
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22922 15988 22928 16040
rect 22980 16037 22986 16040
rect 22980 16031 22995 16037
rect 22983 16028 22995 16031
rect 23032 16028 23060 16068
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 25774 16056 25780 16108
rect 25832 16096 25838 16108
rect 27172 16096 27200 16136
rect 28626 16124 28632 16136
rect 28684 16124 28690 16176
rect 25832 16068 27200 16096
rect 25832 16056 25838 16068
rect 27522 16056 27528 16108
rect 27580 16056 27586 16108
rect 27617 16099 27675 16105
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 28166 16096 28172 16108
rect 27663 16068 28172 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 28166 16056 28172 16068
rect 28224 16056 28230 16108
rect 30190 16056 30196 16108
rect 30248 16096 30254 16108
rect 30392 16096 30420 16195
rect 30248 16068 30420 16096
rect 30248 16056 30254 16068
rect 22983 16000 23060 16028
rect 22983 15997 22995 16000
rect 22980 15991 22995 15997
rect 22980 15988 22986 15991
rect 23566 15988 23572 16040
rect 23624 16028 23630 16040
rect 24029 16031 24087 16037
rect 24029 16028 24041 16031
rect 23624 16000 24041 16028
rect 23624 15988 23630 16000
rect 24029 15997 24041 16000
rect 24075 15997 24087 16031
rect 24029 15991 24087 15997
rect 24121 16031 24179 16037
rect 24121 15997 24133 16031
rect 24167 16028 24179 16031
rect 28718 16028 28724 16040
rect 24167 16000 28724 16028
rect 24167 15997 24179 16000
rect 24121 15991 24179 15997
rect 21174 15920 21180 15972
rect 21232 15960 21238 15972
rect 21542 15960 21548 15972
rect 21232 15932 21548 15960
rect 21232 15920 21238 15932
rect 21542 15920 21548 15932
rect 21600 15920 21606 15972
rect 22649 15963 22707 15969
rect 22649 15929 22661 15963
rect 22695 15960 22707 15963
rect 22695 15932 23888 15960
rect 22695 15929 22707 15932
rect 22649 15923 22707 15929
rect 21048 15864 21128 15892
rect 21048 15852 21054 15864
rect 21266 15852 21272 15904
rect 21324 15892 21330 15904
rect 23290 15892 23296 15904
rect 21324 15864 23296 15892
rect 21324 15852 21330 15864
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 23860 15901 23888 15932
rect 23934 15920 23940 15972
rect 23992 15960 23998 15972
rect 24136 15960 24164 15991
rect 28718 15988 28724 16000
rect 28776 15988 28782 16040
rect 30374 15988 30380 16040
rect 30432 15988 30438 16040
rect 30469 16031 30527 16037
rect 30469 15997 30481 16031
rect 30515 16028 30527 16031
rect 30742 16028 30748 16040
rect 30515 16000 30748 16028
rect 30515 15997 30527 16000
rect 30469 15991 30527 15997
rect 23992 15932 24164 15960
rect 24305 15963 24363 15969
rect 23992 15920 23998 15932
rect 24305 15929 24317 15963
rect 24351 15960 24363 15963
rect 24351 15932 24440 15960
rect 24351 15929 24363 15932
rect 24305 15923 24363 15929
rect 24412 15904 24440 15932
rect 26694 15920 26700 15972
rect 26752 15960 26758 15972
rect 27430 15960 27436 15972
rect 26752 15932 27436 15960
rect 26752 15920 26758 15932
rect 27430 15920 27436 15932
rect 27488 15920 27494 15972
rect 29730 15920 29736 15972
rect 29788 15960 29794 15972
rect 30484 15960 30512 15991
rect 30742 15988 30748 16000
rect 30800 15988 30806 16040
rect 29788 15932 30512 15960
rect 30653 15963 30711 15969
rect 29788 15920 29794 15932
rect 30653 15929 30665 15963
rect 30699 15929 30711 15963
rect 30653 15923 30711 15929
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15861 23903 15895
rect 23845 15855 23903 15861
rect 24394 15852 24400 15904
rect 24452 15852 24458 15904
rect 27522 15852 27528 15904
rect 27580 15852 27586 15904
rect 30466 15852 30472 15904
rect 30524 15892 30530 15904
rect 30668 15892 30696 15923
rect 30524 15864 30696 15892
rect 30524 15852 30530 15864
rect 552 15802 31808 15824
rect 552 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 15946 15802
rect 15998 15750 16010 15802
rect 16062 15750 16074 15802
rect 16126 15750 16138 15802
rect 16190 15750 16202 15802
rect 16254 15750 23720 15802
rect 23772 15750 23784 15802
rect 23836 15750 23848 15802
rect 23900 15750 23912 15802
rect 23964 15750 23976 15802
rect 24028 15750 31494 15802
rect 31546 15750 31558 15802
rect 31610 15750 31622 15802
rect 31674 15750 31686 15802
rect 31738 15750 31750 15802
rect 31802 15750 31808 15802
rect 552 15728 31808 15750
rect 1026 15648 1032 15700
rect 1084 15648 1090 15700
rect 1121 15691 1179 15697
rect 1121 15657 1133 15691
rect 1167 15657 1179 15691
rect 5169 15691 5227 15697
rect 1121 15651 1179 15657
rect 3344 15660 4844 15688
rect 937 15555 995 15561
rect 937 15521 949 15555
rect 983 15552 995 15555
rect 1044 15552 1072 15648
rect 1136 15620 1164 15651
rect 1489 15623 1547 15629
rect 1489 15620 1501 15623
rect 1136 15592 1501 15620
rect 1489 15589 1501 15592
rect 1535 15589 1547 15623
rect 2774 15620 2780 15632
rect 2714 15592 2780 15620
rect 1489 15583 1547 15589
rect 2774 15580 2780 15592
rect 2832 15620 2838 15632
rect 3344 15620 3372 15660
rect 2832 15592 3372 15620
rect 2832 15580 2838 15592
rect 4816 15564 4844 15660
rect 5169 15657 5181 15691
rect 5215 15688 5227 15691
rect 5350 15688 5356 15700
rect 5215 15660 5356 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 6086 15648 6092 15700
rect 6144 15648 6150 15700
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 6638 15688 6644 15700
rect 6595 15660 6644 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 9306 15688 9312 15700
rect 7300 15660 9312 15688
rect 983 15524 1072 15552
rect 3145 15555 3203 15561
rect 983 15521 995 15524
rect 937 15515 995 15521
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 3326 15552 3332 15564
rect 3191 15524 3332 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4798 15512 4804 15564
rect 4856 15512 4862 15564
rect 1213 15487 1271 15493
rect 1213 15484 1225 15487
rect 952 15456 1225 15484
rect 952 15360 980 15456
rect 1213 15453 1225 15456
rect 1259 15484 1271 15487
rect 2682 15484 2688 15496
rect 1259 15456 2688 15484
rect 1259 15453 1271 15456
rect 1213 15447 1271 15453
rect 2682 15444 2688 15456
rect 2740 15484 2746 15496
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 2740 15456 3433 15484
rect 2740 15444 2746 15456
rect 3421 15453 3433 15456
rect 3467 15453 3479 15487
rect 3697 15487 3755 15493
rect 3697 15484 3709 15487
rect 3421 15447 3479 15453
rect 3528 15456 3709 15484
rect 3329 15419 3387 15425
rect 3329 15385 3341 15419
rect 3375 15416 3387 15419
rect 3528 15416 3556 15456
rect 3697 15453 3709 15456
rect 3743 15453 3755 15487
rect 3697 15447 3755 15453
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4062 15484 4068 15496
rect 3844 15456 4068 15484
rect 3844 15444 3850 15456
rect 4062 15444 4068 15456
rect 4120 15484 4126 15496
rect 4120 15456 5120 15484
rect 4120 15444 4126 15456
rect 3375 15388 3556 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 934 15308 940 15360
rect 992 15308 998 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2924 15320 2973 15348
rect 2924 15308 2930 15320
rect 2961 15317 2973 15320
rect 3007 15348 3019 15351
rect 4982 15348 4988 15360
rect 3007 15320 4988 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5092 15348 5120 15456
rect 6104 15416 6132 15648
rect 6196 15620 6224 15648
rect 7300 15629 7328 15660
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9398 15648 9404 15700
rect 9456 15648 9462 15700
rect 9490 15648 9496 15700
rect 9548 15648 9554 15700
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 11054 15688 11060 15700
rect 9640 15660 11060 15688
rect 9640 15648 9646 15660
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11756 15660 11989 15688
rect 11756 15648 11762 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 11977 15651 12035 15657
rect 12526 15648 12532 15700
rect 12584 15648 12590 15700
rect 12710 15648 12716 15700
rect 12768 15648 12774 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 14182 15688 14188 15700
rect 13679 15660 14188 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 14424 15660 15301 15688
rect 14424 15648 14430 15660
rect 15289 15657 15301 15660
rect 15335 15688 15347 15691
rect 16298 15688 16304 15700
rect 15335 15660 16304 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 16540 15660 17233 15688
rect 16540 15648 16546 15660
rect 17221 15657 17233 15660
rect 17267 15688 17279 15691
rect 17494 15688 17500 15700
rect 17267 15660 17500 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 17586 15648 17592 15700
rect 17644 15688 17650 15700
rect 18233 15691 18291 15697
rect 18233 15688 18245 15691
rect 17644 15660 18245 15688
rect 17644 15648 17650 15660
rect 18233 15657 18245 15660
rect 18279 15657 18291 15691
rect 18233 15651 18291 15657
rect 18322 15648 18328 15700
rect 18380 15648 18386 15700
rect 18506 15648 18512 15700
rect 18564 15648 18570 15700
rect 18785 15691 18843 15697
rect 18785 15657 18797 15691
rect 18831 15688 18843 15691
rect 18966 15688 18972 15700
rect 18831 15660 18972 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19426 15688 19432 15700
rect 19168 15660 19432 15688
rect 7285 15623 7343 15629
rect 7285 15620 7297 15623
rect 6196 15592 7297 15620
rect 7285 15589 7297 15592
rect 7331 15589 7343 15623
rect 7285 15583 7343 15589
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 9416 15620 9444 15648
rect 7984 15592 9444 15620
rect 9508 15620 9536 15648
rect 9508 15592 9904 15620
rect 7984 15580 7990 15592
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 6730 15552 6736 15564
rect 6687 15524 6736 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 6472 15484 6500 15515
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15552 6975 15555
rect 7006 15552 7012 15564
rect 6963 15524 7012 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8536 15524 9045 15552
rect 8536 15512 8542 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 9122 15512 9128 15564
rect 9180 15552 9186 15564
rect 9876 15561 9904 15592
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10870 15620 10876 15632
rect 10008 15592 10876 15620
rect 10008 15580 10014 15592
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 12221 15623 12279 15629
rect 12221 15620 12233 15623
rect 11848 15592 12233 15620
rect 11848 15580 11854 15592
rect 12221 15589 12233 15592
rect 12267 15589 12279 15623
rect 12221 15583 12279 15589
rect 12437 15623 12495 15629
rect 12437 15589 12449 15623
rect 12483 15589 12495 15623
rect 12728 15620 12756 15648
rect 16206 15620 16212 15632
rect 12728 15592 12848 15620
rect 12437 15583 12495 15589
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 9180 15524 9321 15552
rect 9180 15512 9186 15524
rect 9309 15521 9321 15524
rect 9355 15521 9367 15555
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9309 15515 9367 15521
rect 9416 15524 9689 15552
rect 6840 15484 6868 15512
rect 6472 15456 6868 15484
rect 8036 15484 8064 15512
rect 8036 15456 9352 15484
rect 9324 15428 9352 15456
rect 9416 15428 9444 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15521 9919 15555
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 9861 15515 9919 15521
rect 9968 15524 10977 15552
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 9766 15484 9772 15496
rect 9631 15456 9772 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9125 15419 9183 15425
rect 9125 15416 9137 15419
rect 6104 15388 9137 15416
rect 9125 15385 9137 15388
rect 9171 15385 9183 15419
rect 9125 15379 9183 15385
rect 9306 15376 9312 15428
rect 9364 15376 9370 15428
rect 9398 15376 9404 15428
rect 9456 15376 9462 15428
rect 9508 15416 9536 15447
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9858 15416 9864 15428
rect 9508 15388 9864 15416
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 5092 15320 6837 15348
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 9968 15348 9996 15524
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 11146 15512 11152 15564
rect 11204 15512 11210 15564
rect 11606 15512 11612 15564
rect 11664 15552 11670 15564
rect 12452 15552 12480 15583
rect 12710 15552 12716 15564
rect 11664 15524 12480 15552
rect 12674 15524 12716 15552
rect 11664 15512 11670 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12820 15561 12848 15592
rect 15396 15592 16212 15620
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15521 12863 15555
rect 12805 15515 12863 15521
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 13354 15512 13360 15564
rect 13412 15512 13418 15564
rect 14182 15512 14188 15564
rect 14240 15512 14246 15564
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 14700 15524 14749 15552
rect 14700 15512 14706 15524
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 15396 15561 15424 15592
rect 16206 15580 16212 15592
rect 16264 15620 16270 15632
rect 16853 15623 16911 15629
rect 16264 15592 16712 15620
rect 16264 15580 16270 15592
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14884 15524 14933 15552
rect 14884 15512 14890 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15521 15439 15555
rect 15381 15515 15439 15521
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 16022 15552 16028 15564
rect 15611 15524 16028 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 10836 15456 11345 15484
rect 10836 15444 10842 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 10502 15376 10508 15428
rect 10560 15416 10566 15428
rect 10965 15419 11023 15425
rect 10965 15416 10977 15419
rect 10560 15388 10977 15416
rect 10560 15376 10566 15388
rect 10965 15385 10977 15388
rect 11011 15385 11023 15419
rect 10965 15379 11023 15385
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 11348 15416 11376 15447
rect 11514 15444 11520 15496
rect 11572 15444 11578 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 13096 15456 16129 15484
rect 11882 15416 11888 15428
rect 11348 15388 11888 15416
rect 11882 15376 11888 15388
rect 11940 15376 11946 15428
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 12032 15388 12296 15416
rect 12032 15376 12038 15388
rect 8720 15320 9996 15348
rect 8720 15308 8726 15320
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10744 15320 10793 15348
rect 10744 15308 10750 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 11072 15348 11100 15376
rect 12268 15357 12296 15388
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 11072 15320 12081 15348
rect 10781 15311 10839 15317
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12986 15348 12992 15360
rect 12299 15320 12992 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 13096 15357 13124 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16316 15484 16344 15515
rect 16482 15512 16488 15564
rect 16540 15512 16546 15564
rect 16574 15512 16580 15564
rect 16632 15512 16638 15564
rect 16684 15552 16712 15592
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 16942 15620 16948 15632
rect 16899 15592 16948 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 16942 15580 16948 15592
rect 17000 15580 17006 15632
rect 17069 15623 17127 15629
rect 17069 15589 17081 15623
rect 17115 15620 17127 15623
rect 17402 15620 17408 15632
rect 17115 15592 17408 15620
rect 17115 15589 17127 15592
rect 17069 15583 17127 15589
rect 17402 15580 17408 15592
rect 17460 15580 17466 15632
rect 18524 15620 18552 15648
rect 18874 15620 18880 15632
rect 17880 15592 18552 15620
rect 18800 15592 18880 15620
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16684 15524 16773 15552
rect 16761 15521 16773 15524
rect 16807 15552 16819 15555
rect 17880 15552 17908 15592
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 16807 15524 17908 15552
rect 17972 15524 18521 15552
rect 16807 15521 16819 15524
rect 16761 15515 16819 15521
rect 17972 15484 18000 15524
rect 18509 15521 18521 15524
rect 18555 15552 18567 15555
rect 18800 15552 18828 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 19168 15620 19196 15660
rect 19426 15648 19432 15660
rect 19484 15688 19490 15700
rect 22554 15688 22560 15700
rect 19484 15660 22560 15688
rect 19484 15648 19490 15660
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23198 15648 23204 15700
rect 23256 15648 23262 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 24026 15688 24032 15700
rect 23440 15660 24032 15688
rect 23440 15648 23446 15660
rect 24026 15648 24032 15660
rect 24084 15648 24090 15700
rect 24302 15688 24308 15700
rect 24136 15660 24308 15688
rect 19168 15592 19272 15620
rect 19244 15561 19272 15592
rect 19702 15580 19708 15632
rect 19760 15620 19766 15632
rect 21542 15620 21548 15632
rect 19760 15592 21548 15620
rect 19760 15580 19766 15592
rect 21542 15580 21548 15592
rect 21600 15580 21606 15632
rect 22833 15623 22891 15629
rect 22833 15620 22845 15623
rect 21652 15592 22845 15620
rect 18555 15524 18828 15552
rect 19061 15555 19119 15561
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 19061 15521 19073 15555
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 19153 15555 19211 15561
rect 19153 15521 19165 15555
rect 19199 15521 19211 15555
rect 19244 15555 19308 15561
rect 19244 15524 19262 15555
rect 19153 15515 19211 15521
rect 19250 15521 19262 15524
rect 19296 15521 19308 15555
rect 19250 15515 19308 15521
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15550 19487 15555
rect 19518 15550 19524 15564
rect 19475 15522 19524 15550
rect 19475 15521 19487 15522
rect 19429 15515 19487 15521
rect 16316 15456 18000 15484
rect 16117 15447 16175 15453
rect 16776 15428 16804 15456
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18598 15493 18604 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 18104 15456 18153 15484
rect 18104 15444 18110 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18597 15447 18604 15493
rect 18656 15484 18662 15496
rect 18656 15456 18697 15484
rect 16393 15419 16451 15425
rect 16393 15385 16405 15419
rect 16439 15385 16451 15419
rect 16393 15379 16451 15385
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15317 13139 15351
rect 13081 15311 13139 15317
rect 14366 15308 14372 15360
rect 14424 15308 14430 15360
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 15746 15348 15752 15360
rect 15151 15320 15752 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 16408 15348 16436 15379
rect 16758 15376 16764 15428
rect 16816 15376 16822 15428
rect 17770 15416 17776 15428
rect 16970 15388 17776 15416
rect 16970 15348 16998 15388
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 18156 15416 18184 15447
rect 18598 15444 18604 15447
rect 18656 15444 18662 15456
rect 18966 15444 18972 15496
rect 19024 15444 19030 15496
rect 19076 15416 19104 15515
rect 18156 15388 19104 15416
rect 19168 15416 19196 15515
rect 19518 15512 19524 15522
rect 19576 15512 19582 15564
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19629 15484 19657 15515
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 20717 15555 20775 15561
rect 20717 15552 20729 15555
rect 20680 15524 20729 15552
rect 20680 15512 20686 15524
rect 20717 15521 20729 15524
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 20990 15512 20996 15564
rect 21048 15512 21054 15564
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21652 15552 21680 15592
rect 22833 15589 22845 15592
rect 22879 15589 22891 15623
rect 22833 15583 22891 15589
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 23216 15620 23244 15648
rect 23072 15592 23704 15620
rect 23072 15580 23078 15592
rect 21508 15524 21680 15552
rect 21508 15512 21514 15524
rect 22186 15512 22192 15564
rect 22244 15512 22250 15564
rect 22738 15512 22744 15564
rect 22796 15512 22802 15564
rect 22925 15555 22983 15561
rect 22925 15552 22937 15555
rect 22848 15524 22937 15552
rect 20438 15484 20444 15496
rect 19629 15456 20444 15484
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 21376 15484 21404 15512
rect 20588 15456 21404 15484
rect 20588 15444 20594 15456
rect 19521 15419 19579 15425
rect 19521 15416 19533 15419
rect 19168 15388 19533 15416
rect 16408 15320 16998 15348
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15348 17095 15351
rect 17586 15348 17592 15360
rect 17083 15320 17592 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17586 15308 17592 15320
rect 17644 15348 17650 15360
rect 17862 15348 17868 15360
rect 17644 15320 17868 15348
rect 17644 15308 17650 15320
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 19168 15348 19196 15388
rect 19521 15385 19533 15388
rect 19567 15385 19579 15419
rect 20806 15416 20812 15428
rect 19521 15379 19579 15385
rect 19628 15388 20812 15416
rect 18380 15320 19196 15348
rect 18380 15308 18386 15320
rect 19242 15308 19248 15360
rect 19300 15348 19306 15360
rect 19628 15348 19656 15388
rect 20806 15376 20812 15388
rect 20864 15416 20870 15428
rect 20901 15419 20959 15425
rect 20901 15416 20913 15419
rect 20864 15388 20913 15416
rect 20864 15376 20870 15388
rect 20901 15385 20913 15388
rect 20947 15385 20959 15419
rect 21468 15416 21496 15512
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 20901 15379 20959 15385
rect 21008 15388 21496 15416
rect 22296 15416 22324 15447
rect 22848 15416 22876 15524
rect 22925 15521 22937 15524
rect 22971 15552 22983 15555
rect 23198 15552 23204 15564
rect 22971 15524 23204 15552
rect 22971 15521 22983 15524
rect 22925 15515 22983 15521
rect 23198 15512 23204 15524
rect 23256 15512 23262 15564
rect 23676 15552 23704 15592
rect 23750 15580 23756 15632
rect 23808 15620 23814 15632
rect 24136 15629 24164 15660
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 24489 15691 24547 15697
rect 24489 15657 24501 15691
rect 24535 15688 24547 15691
rect 24670 15688 24676 15700
rect 24535 15660 24676 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 24854 15648 24860 15700
rect 24912 15688 24918 15700
rect 24949 15691 25007 15697
rect 24949 15688 24961 15691
rect 24912 15660 24961 15688
rect 24912 15648 24918 15660
rect 24949 15657 24961 15660
rect 24995 15657 25007 15691
rect 24949 15651 25007 15657
rect 26142 15648 26148 15700
rect 26200 15688 26206 15700
rect 26200 15660 27200 15688
rect 26200 15648 26206 15660
rect 24121 15623 24179 15629
rect 24121 15620 24133 15623
rect 23808 15592 24133 15620
rect 23808 15580 23814 15592
rect 24121 15589 24133 15592
rect 24167 15589 24179 15623
rect 24121 15583 24179 15589
rect 24210 15580 24216 15632
rect 24268 15620 24274 15632
rect 25225 15623 25283 15629
rect 25225 15620 25237 15623
rect 24268 15592 25084 15620
rect 24268 15580 24274 15592
rect 25056 15564 25084 15592
rect 25148 15592 25237 15620
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 23676 15524 23857 15552
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24394 15561 24400 15564
rect 24351 15555 24400 15561
rect 23992 15524 24037 15552
rect 23992 15512 23998 15524
rect 24351 15521 24363 15555
rect 24397 15521 24400 15555
rect 24351 15515 24400 15521
rect 24394 15512 24400 15515
rect 24452 15512 24458 15564
rect 25038 15512 25044 15564
rect 25096 15512 25102 15564
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 23952 15484 23980 15512
rect 25148 15484 25176 15592
rect 25225 15589 25237 15592
rect 25271 15589 25283 15623
rect 25225 15583 25283 15589
rect 25685 15623 25743 15629
rect 25685 15589 25697 15623
rect 25731 15620 25743 15623
rect 26418 15620 26424 15632
rect 25731 15592 26424 15620
rect 25731 15589 25743 15592
rect 25685 15583 25743 15589
rect 25410 15577 25468 15583
rect 26418 15580 26424 15592
rect 26476 15580 26482 15632
rect 25410 15543 25422 15577
rect 25456 15543 25468 15577
rect 25410 15537 25468 15543
rect 25777 15555 25835 15561
rect 25424 15524 25453 15537
rect 25424 15496 25452 15524
rect 25777 15521 25789 15555
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 25869 15555 25927 15561
rect 25869 15521 25881 15555
rect 25915 15521 25927 15555
rect 25869 15515 25927 15521
rect 26053 15555 26111 15561
rect 26053 15521 26065 15555
rect 26099 15521 26111 15555
rect 26053 15515 26111 15521
rect 25222 15484 25228 15496
rect 23532 15456 23980 15484
rect 24228 15456 25228 15484
rect 23532 15444 23538 15456
rect 24228 15428 24256 15456
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25406 15444 25412 15496
rect 25464 15444 25470 15496
rect 25682 15444 25688 15496
rect 25740 15444 25746 15496
rect 22296 15388 22876 15416
rect 19300 15320 19656 15348
rect 19300 15308 19306 15320
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 21008 15348 21036 15388
rect 24210 15376 24216 15428
rect 24268 15376 24274 15428
rect 24578 15376 24584 15428
rect 24636 15376 24642 15428
rect 24670 15376 24676 15428
rect 24728 15416 24734 15428
rect 25792 15416 25820 15515
rect 24728 15388 25820 15416
rect 24728 15376 24734 15388
rect 20128 15320 21036 15348
rect 22373 15351 22431 15357
rect 20128 15308 20134 15320
rect 22373 15317 22385 15351
rect 22419 15348 22431 15351
rect 22554 15348 22560 15360
rect 22419 15320 22560 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 22554 15308 22560 15320
rect 22612 15308 22618 15360
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 24596 15348 24624 15376
rect 23624 15320 24624 15348
rect 23624 15308 23630 15320
rect 25314 15308 25320 15360
rect 25372 15348 25378 15360
rect 25501 15351 25559 15357
rect 25501 15348 25513 15351
rect 25372 15320 25513 15348
rect 25372 15308 25378 15320
rect 25501 15317 25513 15320
rect 25547 15317 25559 15351
rect 25884 15348 25912 15515
rect 26068 15428 26096 15515
rect 26142 15512 26148 15564
rect 26200 15512 26206 15564
rect 26237 15555 26295 15561
rect 26237 15521 26249 15555
rect 26283 15552 26295 15555
rect 26605 15555 26663 15561
rect 26605 15552 26617 15555
rect 26283 15524 26617 15552
rect 26283 15521 26295 15524
rect 26237 15515 26295 15521
rect 26605 15521 26617 15524
rect 26651 15521 26663 15555
rect 26605 15515 26663 15521
rect 26786 15512 26792 15564
rect 26844 15512 26850 15564
rect 27172 15561 27200 15660
rect 27522 15648 27528 15700
rect 27580 15688 27586 15700
rect 27985 15691 28043 15697
rect 27985 15688 27997 15691
rect 27580 15660 27997 15688
rect 27580 15648 27586 15660
rect 27985 15657 27997 15660
rect 28031 15657 28043 15691
rect 27985 15651 28043 15657
rect 29546 15648 29552 15700
rect 29604 15688 29610 15700
rect 29917 15691 29975 15697
rect 29917 15688 29929 15691
rect 29604 15660 29929 15688
rect 29604 15648 29610 15660
rect 29917 15657 29929 15660
rect 29963 15657 29975 15691
rect 29917 15651 29975 15657
rect 27341 15623 27399 15629
rect 27341 15589 27353 15623
rect 27387 15620 27399 15623
rect 27617 15623 27675 15629
rect 27617 15620 27629 15623
rect 27387 15592 27629 15620
rect 27387 15589 27399 15592
rect 27341 15583 27399 15589
rect 27617 15589 27629 15592
rect 27663 15589 27675 15623
rect 27617 15583 27675 15589
rect 27706 15580 27712 15632
rect 27764 15580 27770 15632
rect 28169 15623 28227 15629
rect 28169 15589 28181 15623
rect 28215 15620 28227 15623
rect 29564 15620 29592 15648
rect 28215 15592 28672 15620
rect 28215 15589 28227 15592
rect 28169 15583 28227 15589
rect 28644 15564 28672 15592
rect 29288 15592 29592 15620
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15521 27215 15555
rect 27157 15515 27215 15521
rect 27430 15512 27436 15564
rect 27488 15512 27494 15564
rect 27522 15512 27528 15564
rect 27580 15552 27586 15564
rect 27801 15555 27859 15561
rect 27801 15552 27813 15555
rect 27580 15524 27813 15552
rect 27580 15512 27586 15524
rect 27801 15521 27813 15524
rect 27847 15521 27859 15555
rect 27801 15515 27859 15521
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28077 15555 28135 15561
rect 28077 15552 28089 15555
rect 28040 15524 28089 15552
rect 28040 15512 28046 15524
rect 28077 15521 28089 15524
rect 28123 15521 28135 15555
rect 28077 15515 28135 15521
rect 28258 15512 28264 15564
rect 28316 15552 28322 15564
rect 28353 15555 28411 15561
rect 28353 15552 28365 15555
rect 28316 15524 28365 15552
rect 28316 15512 28322 15524
rect 28353 15521 28365 15524
rect 28399 15521 28411 15555
rect 28353 15515 28411 15521
rect 28626 15512 28632 15564
rect 28684 15512 28690 15564
rect 29288 15561 29316 15592
rect 30374 15580 30380 15632
rect 30432 15580 30438 15632
rect 29273 15555 29331 15561
rect 29273 15521 29285 15555
rect 29319 15521 29331 15555
rect 29273 15515 29331 15521
rect 29362 15512 29368 15564
rect 29420 15512 29426 15564
rect 29457 15555 29515 15561
rect 29457 15521 29469 15555
rect 29503 15521 29515 15555
rect 29457 15515 29515 15521
rect 26160 15484 26188 15512
rect 26881 15487 26939 15493
rect 26881 15484 26893 15487
rect 26160 15456 26893 15484
rect 26881 15453 26893 15456
rect 26927 15453 26939 15487
rect 26881 15447 26939 15453
rect 26973 15487 27031 15493
rect 26973 15453 26985 15487
rect 27019 15484 27031 15487
rect 28997 15487 29055 15493
rect 28997 15484 29009 15487
rect 27019 15456 29009 15484
rect 27019 15453 27031 15456
rect 26973 15447 27031 15453
rect 28997 15453 29009 15456
rect 29043 15453 29055 15487
rect 29472 15484 29500 15515
rect 29638 15512 29644 15564
rect 29696 15512 29702 15564
rect 29730 15512 29736 15564
rect 29788 15552 29794 15564
rect 30101 15555 30159 15561
rect 30101 15552 30113 15555
rect 29788 15524 30113 15552
rect 29788 15512 29794 15524
rect 30101 15521 30113 15524
rect 30147 15521 30159 15555
rect 30101 15515 30159 15521
rect 30190 15512 30196 15564
rect 30248 15512 30254 15564
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15552 30343 15555
rect 30392 15552 30420 15580
rect 30558 15552 30564 15564
rect 30331 15524 30564 15552
rect 30331 15521 30343 15524
rect 30285 15515 30343 15521
rect 30558 15512 30564 15524
rect 30616 15512 30622 15564
rect 29822 15484 29828 15496
rect 29472 15456 29828 15484
rect 28997 15447 29055 15453
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 30374 15444 30380 15496
rect 30432 15444 30438 15496
rect 26050 15376 26056 15428
rect 26108 15376 26114 15428
rect 28534 15348 28540 15360
rect 25884 15320 28540 15348
rect 25501 15311 25559 15317
rect 28534 15308 28540 15320
rect 28592 15308 28598 15360
rect 552 15258 31648 15280
rect 552 15206 4285 15258
rect 4337 15206 4349 15258
rect 4401 15206 4413 15258
rect 4465 15206 4477 15258
rect 4529 15206 4541 15258
rect 4593 15206 12059 15258
rect 12111 15206 12123 15258
rect 12175 15206 12187 15258
rect 12239 15206 12251 15258
rect 12303 15206 12315 15258
rect 12367 15206 19833 15258
rect 19885 15206 19897 15258
rect 19949 15206 19961 15258
rect 20013 15206 20025 15258
rect 20077 15206 20089 15258
rect 20141 15206 27607 15258
rect 27659 15206 27671 15258
rect 27723 15206 27735 15258
rect 27787 15206 27799 15258
rect 27851 15206 27863 15258
rect 27915 15206 31648 15258
rect 552 15184 31648 15206
rect 3329 15147 3387 15153
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3418 15144 3424 15156
rect 3375 15116 3424 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3694 15104 3700 15156
rect 3752 15104 3758 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 5592 15116 6653 15144
rect 5592 15104 5598 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 8389 15147 8447 15153
rect 8389 15113 8401 15147
rect 8435 15144 8447 15147
rect 8846 15144 8852 15156
rect 8435 15116 8852 15144
rect 8435 15113 8447 15116
rect 8389 15107 8447 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 10226 15104 10232 15156
rect 10284 15104 10290 15156
rect 10428 15116 11836 15144
rect 3142 15076 3148 15088
rect 2608 15048 3148 15076
rect 750 14968 756 15020
rect 808 15008 814 15020
rect 2608 15008 2636 15048
rect 3142 15036 3148 15048
rect 3200 15036 3206 15088
rect 3712 15076 3740 15104
rect 3452 15048 3648 15076
rect 3712 15048 4568 15076
rect 808 14980 2636 15008
rect 808 14968 814 14980
rect 2682 14968 2688 15020
rect 2740 15008 2746 15020
rect 3452 15008 3480 15048
rect 2740 14980 3480 15008
rect 2740 14968 2746 14980
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 3620 15008 3648 15048
rect 4540 15017 4568 15048
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 10428 15076 10456 15116
rect 11808 15088 11836 15116
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 16117 15147 16175 15153
rect 11940 15116 12664 15144
rect 11940 15104 11946 15116
rect 9180 15048 10456 15076
rect 9180 15036 9186 15048
rect 11790 15036 11796 15088
rect 11848 15036 11854 15088
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 3620 14980 4261 15008
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 6822 14968 6828 15020
rect 6880 15008 6886 15020
rect 8570 15008 8576 15020
rect 6880 14980 8576 15008
rect 6880 14968 6886 14980
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 8849 15011 8907 15017
rect 8849 15008 8861 15011
rect 8680 14980 8861 15008
rect 845 14943 903 14949
rect 845 14909 857 14943
rect 891 14940 903 14943
rect 934 14940 940 14952
rect 891 14912 940 14940
rect 891 14909 903 14912
rect 845 14903 903 14909
rect 934 14900 940 14912
rect 992 14900 998 14952
rect 1210 14900 1216 14952
rect 1268 14900 1274 14952
rect 3528 14925 3556 14968
rect 3513 14919 3571 14925
rect 3513 14885 3525 14919
rect 3559 14885 3571 14919
rect 3602 14900 3608 14952
rect 3660 14940 3666 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 3660 14912 4169 14940
rect 3660 14900 3666 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 6914 14940 6920 14952
rect 5934 14912 6920 14940
rect 4157 14903 4215 14909
rect 6914 14900 6920 14912
rect 6972 14940 6978 14952
rect 7374 14940 7380 14952
rect 6972 14912 7380 14940
rect 6972 14900 6978 14912
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 8680 14940 8708 14980
rect 8849 14977 8861 14980
rect 8895 14977 8907 15011
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8849 14971 8907 14977
rect 8956 14980 9045 15008
rect 8956 14952 8984 14980
rect 9033 14977 9045 14980
rect 9079 14977 9091 15011
rect 9582 15008 9588 15020
rect 9033 14971 9091 14977
rect 9232 14980 9588 15008
rect 7984 14912 8708 14940
rect 7984 14900 7990 14912
rect 8754 14900 8760 14952
rect 8812 14900 8818 14952
rect 8938 14900 8944 14952
rect 8996 14900 9002 14952
rect 9232 14949 9260 14980
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 10008 14980 10333 15008
rect 10008 14968 10014 14980
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 10686 15008 10692 15020
rect 10643 14980 10692 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11606 15008 11612 15020
rect 11112 14980 11612 15008
rect 11112 14968 11118 14980
rect 11606 14968 11612 14980
rect 11664 15008 11670 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11664 14980 12081 15008
rect 11664 14968 11670 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12636 15008 12664 15116
rect 16117 15113 16129 15147
rect 16163 15144 16175 15147
rect 16206 15144 16212 15156
rect 16163 15116 16212 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15144 16727 15147
rect 16758 15144 16764 15156
rect 16715 15116 16764 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17586 15104 17592 15156
rect 17644 15144 17650 15156
rect 17644 15116 18276 15144
rect 17644 15104 17650 15116
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 13354 15076 13360 15088
rect 12860 15048 13360 15076
rect 12860 15036 12866 15048
rect 13354 15036 13360 15048
rect 13412 15076 13418 15088
rect 17034 15076 17040 15088
rect 13412 15048 17040 15076
rect 13412 15036 13418 15048
rect 17034 15036 17040 15048
rect 17092 15076 17098 15088
rect 17862 15076 17868 15088
rect 17092 15048 17868 15076
rect 17092 15036 17098 15048
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 18248 15076 18276 15116
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18472 15116 18797 15144
rect 18472 15104 18478 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 19518 15104 19524 15156
rect 19576 15104 19582 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20162 15144 20168 15156
rect 19935 15116 20168 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 19536 15076 19564 15104
rect 18248 15048 19564 15076
rect 19720 15076 19748 15107
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 22554 15144 22560 15156
rect 20272 15116 22560 15144
rect 19978 15076 19984 15088
rect 19720 15048 19984 15076
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 12636 14980 14841 15008
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9364 14912 9413 14940
rect 9364 14900 9370 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9490 14900 9496 14952
rect 9548 14900 9554 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2774 14872 2780 14884
rect 2280 14844 2780 14872
rect 2280 14832 2286 14844
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 3513 14879 3571 14885
rect 4798 14832 4804 14884
rect 4856 14832 4862 14884
rect 6104 14844 7144 14872
rect 2590 14764 2596 14816
rect 2648 14813 2654 14816
rect 2648 14807 2697 14813
rect 2648 14773 2651 14807
rect 2685 14773 2697 14807
rect 2648 14767 2697 14773
rect 2648 14764 2654 14767
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 3697 14807 3755 14813
rect 3697 14804 3709 14807
rect 3660 14776 3709 14804
rect 3660 14764 3666 14776
rect 3697 14773 3709 14776
rect 3743 14773 3755 14807
rect 3697 14767 3755 14773
rect 4062 14764 4068 14816
rect 4120 14764 4126 14816
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4614 14804 4620 14816
rect 4304 14776 4620 14804
rect 4304 14764 4310 14776
rect 4614 14764 4620 14776
rect 4672 14804 4678 14816
rect 6104 14804 6132 14844
rect 7116 14816 7144 14844
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 8113 14875 8171 14881
rect 8113 14872 8125 14875
rect 8076 14844 8125 14872
rect 8076 14832 8082 14844
rect 8113 14841 8125 14844
rect 8159 14872 8171 14875
rect 8478 14872 8484 14884
rect 8159 14844 8484 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 4672 14776 6132 14804
rect 4672 14764 4678 14776
rect 6270 14764 6276 14816
rect 6328 14764 6334 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 9030 14804 9036 14816
rect 7156 14776 9036 14804
rect 7156 14764 7162 14776
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9306 14764 9312 14816
rect 9364 14764 9370 14816
rect 9692 14804 9720 14903
rect 9766 14900 9772 14952
rect 9824 14900 9830 14952
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 12434 14900 12440 14952
rect 12492 14900 12498 14952
rect 12636 14940 12664 14980
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12636 14912 12817 14940
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 13740 14949 13768 14980
rect 14829 14977 14841 14980
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 20272 15008 20300 15116
rect 22554 15104 22560 15116
rect 22612 15144 22618 15156
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22612 15116 22661 15144
rect 22612 15104 22618 15116
rect 22649 15113 22661 15116
rect 22695 15144 22707 15147
rect 22738 15144 22744 15156
rect 22695 15116 22744 15144
rect 22695 15113 22707 15116
rect 22649 15107 22707 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 23014 15144 23020 15156
rect 22888 15116 23020 15144
rect 22888 15104 22894 15116
rect 23014 15104 23020 15116
rect 23072 15104 23078 15156
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 25593 15147 25651 15153
rect 23532 15116 25544 15144
rect 23532 15104 23538 15116
rect 20438 15036 20444 15088
rect 20496 15076 20502 15088
rect 22925 15079 22983 15085
rect 20496 15048 22232 15076
rect 20496 15036 20502 15048
rect 22204 15020 22232 15048
rect 22925 15045 22937 15079
rect 22971 15076 22983 15079
rect 25406 15076 25412 15088
rect 22971 15048 25412 15076
rect 22971 15045 22983 15048
rect 22925 15039 22983 15045
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 20898 15008 20904 15020
rect 15344 14980 20300 15008
rect 20364 14980 20904 15008
rect 15344 14968 15350 14980
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 13044 14912 13185 14940
rect 13044 14900 13050 14912
rect 13173 14909 13185 14912
rect 13219 14940 13231 14943
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13219 14912 13553 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 9784 14872 9812 14900
rect 10594 14872 10600 14884
rect 9784 14844 10600 14872
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 12452 14872 12480 14900
rect 14016 14872 14044 14903
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14332 14912 14565 14940
rect 14332 14900 14338 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 14553 14903 14611 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 14645 14903 14703 14909
rect 14752 14912 15485 14940
rect 10928 14844 11086 14872
rect 12452 14844 14044 14872
rect 10928 14832 10934 14844
rect 11882 14804 11888 14816
rect 9692 14776 11888 14804
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14660 14804 14688 14903
rect 14752 14816 14780 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 15488 14872 15516 14903
rect 15654 14900 15660 14952
rect 15712 14900 15718 14952
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 15804 14912 15853 14940
rect 15804 14900 15810 14912
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 16022 14900 16028 14952
rect 16080 14940 16086 14952
rect 16298 14940 16304 14952
rect 16080 14912 16304 14940
rect 16080 14900 16086 14912
rect 16298 14900 16304 14912
rect 16356 14940 16362 14952
rect 16393 14943 16451 14949
rect 16393 14940 16405 14943
rect 16356 14912 16405 14940
rect 16356 14900 16362 14912
rect 16393 14909 16405 14912
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17218 14940 17224 14952
rect 16816 14912 17224 14940
rect 16816 14900 16822 14912
rect 17218 14900 17224 14912
rect 17276 14940 17282 14952
rect 17276 14912 20116 14940
rect 17276 14900 17282 14912
rect 17402 14872 17408 14884
rect 15488 14844 17408 14872
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 19061 14875 19119 14881
rect 19061 14841 19073 14875
rect 19107 14841 19119 14875
rect 19061 14835 19119 14841
rect 13964 14776 14688 14804
rect 13964 14764 13970 14776
rect 14734 14764 14740 14816
rect 14792 14764 14798 14816
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 17218 14804 17224 14816
rect 15528 14776 17224 14804
rect 15528 14764 15534 14776
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 18046 14804 18052 14816
rect 17368 14776 18052 14804
rect 17368 14764 17374 14776
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 19076 14804 19104 14835
rect 19150 14832 19156 14884
rect 19208 14872 19214 14884
rect 19521 14875 19579 14881
rect 19521 14872 19533 14875
rect 19208 14844 19533 14872
rect 19208 14832 19214 14844
rect 19521 14841 19533 14844
rect 19567 14841 19579 14875
rect 19521 14835 19579 14841
rect 19610 14832 19616 14884
rect 19668 14872 19674 14884
rect 19668 14844 20024 14872
rect 19668 14832 19674 14844
rect 19996 14816 20024 14844
rect 19426 14804 19432 14816
rect 19076 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19731 14807 19789 14813
rect 19731 14773 19743 14807
rect 19777 14804 19789 14807
rect 19886 14804 19892 14816
rect 19777 14776 19892 14804
rect 19777 14773 19789 14776
rect 19731 14767 19789 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 19978 14764 19984 14816
rect 20036 14764 20042 14816
rect 20088 14804 20116 14912
rect 20162 14900 20168 14952
rect 20220 14900 20226 14952
rect 20364 14949 20392 14980
rect 20898 14968 20904 14980
rect 20956 15008 20962 15020
rect 21726 15008 21732 15020
rect 20956 14980 21732 15008
rect 20956 14968 20962 14980
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 22186 14968 22192 15020
rect 22244 14968 22250 15020
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 15008 22615 15011
rect 23750 15008 23756 15020
rect 22603 14980 23756 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 20487 14912 20944 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 20180 14872 20208 14900
rect 20622 14872 20628 14884
rect 20180 14844 20628 14872
rect 20622 14832 20628 14844
rect 20680 14832 20686 14884
rect 20916 14816 20944 14912
rect 20990 14900 20996 14952
rect 21048 14900 21054 14952
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21174 14940 21180 14952
rect 21131 14912 21180 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 21174 14900 21180 14912
rect 21232 14940 21238 14952
rect 21634 14940 21640 14952
rect 21232 14912 21640 14940
rect 21232 14900 21238 14912
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 22370 14900 22376 14952
rect 22428 14900 22434 14952
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14940 22707 14943
rect 22830 14940 22836 14952
rect 22695 14912 22836 14940
rect 22695 14909 22707 14912
rect 22649 14903 22707 14909
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23014 14900 23020 14952
rect 23072 14940 23078 14952
rect 23109 14943 23167 14949
rect 23109 14940 23121 14943
rect 23072 14912 23121 14940
rect 23072 14900 23078 14912
rect 23109 14909 23121 14912
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14909 23259 14943
rect 23201 14903 23259 14909
rect 21266 14832 21272 14884
rect 21324 14832 21330 14884
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 22922 14872 22928 14884
rect 22796 14844 22928 14872
rect 22796 14832 22802 14844
rect 22922 14832 22928 14844
rect 22980 14832 22986 14884
rect 23216 14872 23244 14903
rect 23290 14900 23296 14952
rect 23348 14900 23354 14952
rect 23492 14949 23520 14980
rect 23750 14968 23756 14980
rect 23808 14968 23814 15020
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23992 14980 24225 15008
rect 23992 14968 23998 14980
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 24302 14968 24308 15020
rect 24360 15008 24366 15020
rect 24765 15011 24823 15017
rect 24360 14980 24624 15008
rect 24360 14968 24366 14980
rect 23477 14943 23535 14949
rect 23477 14909 23489 14943
rect 23523 14940 23535 14943
rect 23523 14912 23557 14940
rect 23523 14909 23535 14912
rect 23477 14903 23535 14909
rect 24026 14900 24032 14952
rect 24084 14940 24090 14952
rect 24596 14949 24624 14980
rect 24765 14977 24777 15011
rect 24811 15008 24823 15011
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 24811 14980 25237 15008
rect 24811 14977 24823 14980
rect 24765 14971 24823 14977
rect 25225 14977 25237 14980
rect 25271 14977 25283 15011
rect 25225 14971 25283 14977
rect 24397 14943 24455 14949
rect 24397 14940 24409 14943
rect 24084 14912 24409 14940
rect 24084 14900 24090 14912
rect 24228 14884 24256 14912
rect 24397 14909 24409 14912
rect 24443 14909 24455 14943
rect 24397 14903 24455 14909
rect 24581 14943 24639 14949
rect 24581 14909 24593 14943
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 25130 14900 25136 14952
rect 25188 14900 25194 14952
rect 25314 14900 25320 14952
rect 25372 14900 25378 14952
rect 25424 14949 25452 15036
rect 25516 15008 25544 15116
rect 25593 15113 25605 15147
rect 25639 15144 25651 15147
rect 27522 15144 27528 15156
rect 25639 15116 27528 15144
rect 25639 15113 25651 15116
rect 25593 15107 25651 15113
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 28166 15104 28172 15156
rect 28224 15144 28230 15156
rect 28261 15147 28319 15153
rect 28261 15144 28273 15147
rect 28224 15116 28273 15144
rect 28224 15104 28230 15116
rect 28261 15113 28273 15116
rect 28307 15113 28319 15147
rect 28261 15107 28319 15113
rect 28445 15147 28503 15153
rect 28445 15113 28457 15147
rect 28491 15144 28503 15147
rect 29362 15144 29368 15156
rect 28491 15116 29368 15144
rect 28491 15113 28503 15116
rect 28445 15107 28503 15113
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 30190 15104 30196 15156
rect 30248 15104 30254 15156
rect 30834 15104 30840 15156
rect 30892 15104 30898 15156
rect 25682 15036 25688 15088
rect 25740 15076 25746 15088
rect 30208 15076 30236 15104
rect 25740 15048 30236 15076
rect 25740 15036 25746 15048
rect 27154 15008 27160 15020
rect 25516 14980 27160 15008
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14909 25467 14943
rect 25409 14903 25467 14909
rect 26602 14900 26608 14952
rect 26660 14900 26666 14952
rect 26804 14949 26832 14980
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 27982 15008 27988 15020
rect 27632 14980 27988 15008
rect 26789 14943 26847 14949
rect 26789 14909 26801 14943
rect 26835 14909 26847 14943
rect 26789 14903 26847 14909
rect 26878 14900 26884 14952
rect 26936 14900 26942 14952
rect 26970 14900 26976 14952
rect 27028 14940 27034 14952
rect 27632 14940 27660 14980
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 31110 15008 31116 15020
rect 30484 14980 31116 15008
rect 30484 14940 30512 14980
rect 31110 14968 31116 14980
rect 31168 14968 31174 15020
rect 27028 14912 27660 14940
rect 27724 14912 30512 14940
rect 27028 14900 27034 14912
rect 23385 14875 23443 14881
rect 23385 14872 23397 14875
rect 23216 14844 23397 14872
rect 23385 14841 23397 14844
rect 23431 14841 23443 14875
rect 23385 14835 23443 14841
rect 24210 14832 24216 14884
rect 24268 14832 24274 14884
rect 26620 14872 26648 14900
rect 27724 14872 27752 14912
rect 30558 14900 30564 14952
rect 30616 14900 30622 14952
rect 24412 14844 24992 14872
rect 26620 14844 27752 14872
rect 20346 14804 20352 14816
rect 20088 14776 20352 14804
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 20898 14764 20904 14816
rect 20956 14764 20962 14816
rect 21170 14807 21228 14813
rect 21170 14773 21182 14807
rect 21216 14804 21228 14807
rect 24412 14804 24440 14844
rect 21216 14776 24440 14804
rect 21216 14773 21228 14776
rect 21170 14767 21228 14773
rect 24486 14764 24492 14816
rect 24544 14764 24550 14816
rect 24964 14804 24992 14844
rect 28074 14832 28080 14884
rect 28132 14832 28138 14884
rect 30466 14872 30472 14884
rect 28184 14844 30472 14872
rect 26786 14804 26792 14816
rect 24964 14776 26792 14804
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 26878 14764 26884 14816
rect 26936 14804 26942 14816
rect 28184 14804 28212 14844
rect 30466 14832 30472 14844
rect 30524 14832 30530 14884
rect 26936 14776 28212 14804
rect 28287 14807 28345 14813
rect 26936 14764 26942 14776
rect 28287 14773 28299 14807
rect 28333 14804 28345 14807
rect 28442 14804 28448 14816
rect 28333 14776 28448 14804
rect 28333 14773 28345 14776
rect 28287 14767 28345 14773
rect 28442 14764 28448 14776
rect 28500 14764 28506 14816
rect 552 14714 31808 14736
rect 552 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 15946 14714
rect 15998 14662 16010 14714
rect 16062 14662 16074 14714
rect 16126 14662 16138 14714
rect 16190 14662 16202 14714
rect 16254 14662 23720 14714
rect 23772 14662 23784 14714
rect 23836 14662 23848 14714
rect 23900 14662 23912 14714
rect 23964 14662 23976 14714
rect 24028 14662 31494 14714
rect 31546 14662 31558 14714
rect 31610 14662 31622 14714
rect 31674 14662 31686 14714
rect 31738 14662 31750 14714
rect 31802 14662 31808 14714
rect 552 14640 31808 14662
rect 1210 14560 1216 14612
rect 1268 14600 1274 14612
rect 1397 14603 1455 14609
rect 1397 14600 1409 14603
rect 1268 14572 1409 14600
rect 1268 14560 1274 14572
rect 1397 14569 1409 14572
rect 1443 14569 1455 14603
rect 1397 14563 1455 14569
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14569 1731 14603
rect 1673 14563 1731 14569
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1688 14464 1716 14563
rect 2130 14560 2136 14612
rect 2188 14560 2194 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3970 14600 3976 14612
rect 3283 14572 3976 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4706 14560 4712 14612
rect 4764 14560 4770 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 4856 14572 5457 14600
rect 4856 14560 4862 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 6086 14600 6092 14612
rect 5684 14572 6092 14600
rect 5684 14560 5690 14572
rect 6086 14560 6092 14572
rect 6144 14600 6150 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 6144 14572 6285 14600
rect 6144 14560 6150 14572
rect 6273 14569 6285 14572
rect 6319 14569 6331 14603
rect 6273 14563 6331 14569
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7098 14600 7104 14612
rect 7055 14572 7104 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7926 14600 7932 14612
rect 7423 14572 7932 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8662 14560 8668 14612
rect 8720 14560 8726 14612
rect 9214 14600 9220 14612
rect 8772 14572 9220 14600
rect 2148 14532 2176 14560
rect 4724 14532 4752 14560
rect 2148 14504 2268 14532
rect 4462 14504 4752 14532
rect 1627 14436 1716 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1762 14424 1768 14476
rect 1820 14464 1826 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1820 14436 2053 14464
rect 1820 14424 1826 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2056 14328 2084 14427
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 2240 14405 2268 14504
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 7745 14535 7803 14541
rect 7745 14532 7757 14535
rect 7616 14504 7757 14532
rect 7616 14492 7622 14504
rect 7745 14501 7757 14504
rect 7791 14501 7803 14535
rect 7745 14495 7803 14501
rect 2590 14424 2596 14476
rect 2648 14464 2654 14476
rect 2869 14467 2927 14473
rect 2869 14464 2881 14467
rect 2648 14436 2881 14464
rect 2648 14424 2654 14436
rect 2869 14433 2881 14436
rect 2915 14433 2927 14467
rect 2869 14427 2927 14433
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14464 5227 14467
rect 5534 14464 5540 14476
rect 5215 14436 5540 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 2608 14328 2636 14424
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 2056 14300 2636 14328
rect 2700 14328 2728 14359
rect 2774 14356 2780 14408
rect 2832 14356 2838 14408
rect 2884 14396 2912 14427
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 6181 14467 6239 14473
rect 5675 14436 5856 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 4154 14396 4160 14408
rect 2884 14368 4160 14396
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4890 14356 4896 14408
rect 4948 14356 4954 14408
rect 5828 14337 5856 14436
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6270 14464 6276 14476
rect 6227 14436 6276 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6270 14424 6276 14436
rect 6328 14464 6334 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6328 14436 6929 14464
rect 6328 14424 6334 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14365 6883 14399
rect 6932 14396 6960 14427
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 7466 14464 7472 14476
rect 7156 14436 7472 14464
rect 7156 14424 7162 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 8386 14464 8392 14476
rect 7883 14436 8392 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 8478 14424 8484 14476
rect 8536 14424 8542 14476
rect 8772 14473 8800 14572
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 9306 14560 9312 14612
rect 9364 14560 9370 14612
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 9490 14600 9496 14612
rect 9447 14572 9496 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 10100 14572 10149 14600
rect 10100 14560 10106 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 10318 14560 10324 14612
rect 10376 14560 10382 14612
rect 13630 14600 13636 14612
rect 11440 14572 13636 14600
rect 9324 14532 9352 14560
rect 8956 14504 9352 14532
rect 8956 14473 8984 14504
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9640 14504 9873 14532
rect 9640 14492 9646 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 9861 14495 9919 14501
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 8905 14467 8984 14473
rect 8905 14433 8917 14467
rect 8951 14436 8984 14467
rect 8951 14433 8963 14436
rect 8905 14427 8963 14433
rect 9030 14424 9036 14476
rect 9088 14424 9094 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 9263 14467 9321 14473
rect 9263 14433 9275 14467
rect 9309 14464 9321 14467
rect 10042 14464 10048 14476
rect 9309 14436 10048 14464
rect 9309 14433 9321 14436
rect 9263 14427 9321 14433
rect 7282 14396 7288 14408
rect 6932 14368 7288 14396
rect 6825 14359 6883 14365
rect 5813 14331 5871 14337
rect 2700 14300 3924 14328
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 3510 14260 3516 14272
rect 3467 14232 3516 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 3896 14260 3924 14300
rect 5813 14297 5825 14331
rect 5859 14297 5871 14331
rect 5813 14291 5871 14297
rect 4522 14260 4528 14272
rect 3896 14232 4528 14260
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 6380 14260 6408 14359
rect 6840 14328 6868 14359
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7650 14356 7656 14408
rect 7708 14356 7714 14408
rect 8294 14356 8300 14408
rect 8352 14356 8358 14408
rect 8404 14396 8432 14424
rect 9140 14396 9168 14427
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10336 14464 10364 14560
rect 10100 14436 10364 14464
rect 10100 14424 10106 14436
rect 11146 14424 11152 14476
rect 11204 14424 11210 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 11440 14473 11468 14572
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 16209 14603 16267 14609
rect 15528 14572 15792 14600
rect 15528 14560 15534 14572
rect 11974 14532 11980 14544
rect 11624 14504 11980 14532
rect 11333 14467 11391 14473
rect 11333 14464 11345 14467
rect 11296 14436 11345 14464
rect 11296 14424 11302 14436
rect 11333 14433 11345 14436
rect 11379 14433 11391 14467
rect 11333 14427 11391 14433
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 11517 14467 11575 14473
rect 11517 14433 11529 14467
rect 11563 14464 11575 14467
rect 11624 14464 11652 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 12526 14492 12532 14544
rect 12584 14532 12590 14544
rect 14550 14532 14556 14544
rect 12584 14504 14556 14532
rect 12584 14492 12590 14504
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 14826 14532 14832 14544
rect 14752 14504 14832 14532
rect 11563 14436 11652 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 9766 14396 9772 14408
rect 8404 14368 9168 14396
rect 9232 14368 9772 14396
rect 7668 14328 7696 14356
rect 6840 14300 7696 14328
rect 8205 14331 8263 14337
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 9232 14328 9260 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 9916 14368 10273 14396
rect 9916 14356 9922 14368
rect 8251 14300 9260 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9493 14331 9551 14337
rect 9493 14328 9505 14331
rect 9456 14300 9505 14328
rect 9456 14288 9462 14300
rect 9493 14297 9505 14300
rect 9539 14297 9551 14331
rect 10134 14328 10140 14340
rect 9493 14291 9551 14297
rect 9876 14300 10140 14328
rect 7006 14260 7012 14272
rect 6380 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14260 7070 14272
rect 7466 14260 7472 14272
rect 7064 14232 7472 14260
rect 7064 14220 7070 14232
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 9122 14260 9128 14272
rect 8536 14232 9128 14260
rect 8536 14220 8542 14232
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9674 14260 9680 14272
rect 9272 14232 9680 14260
rect 9272 14220 9278 14232
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9876 14269 9904 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10245 14328 10273 14368
rect 10318 14356 10324 14408
rect 10376 14396 10382 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10376 14368 10701 14396
rect 10376 14356 10382 14368
rect 10689 14365 10701 14368
rect 10735 14396 10747 14399
rect 11054 14396 11060 14408
rect 10735 14368 11060 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11624 14328 11652 14436
rect 11698 14424 11704 14476
rect 11756 14424 11762 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 11992 14436 12173 14464
rect 11882 14356 11888 14408
rect 11940 14356 11946 14408
rect 11992 14340 12020 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 12802 14464 12808 14476
rect 12667 14436 12808 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14433 13047 14467
rect 12989 14427 13047 14433
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 13906 14464 13912 14476
rect 13587 14436 13912 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12176 14368 12449 14396
rect 10245 14300 11652 14328
rect 11974 14288 11980 14340
rect 12032 14288 12038 14340
rect 9861 14263 9919 14269
rect 9861 14229 9873 14263
rect 9907 14229 9919 14263
rect 9861 14223 9919 14229
rect 10045 14263 10103 14269
rect 10045 14229 10057 14263
rect 10091 14260 10103 14263
rect 10226 14260 10232 14272
rect 10091 14232 10232 14260
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 12176 14260 12204 14368
rect 12437 14365 12449 14368
rect 12483 14396 12495 14399
rect 13004 14396 13032 14427
rect 12483 14368 13032 14396
rect 13081 14399 13139 14405
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13446 14396 13452 14408
rect 13127 14368 13452 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 13556 14328 13584 14427
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 14642 14424 14648 14476
rect 14700 14424 14706 14476
rect 14752 14473 14780 14504
rect 14826 14492 14832 14504
rect 14884 14532 14890 14544
rect 15378 14532 15384 14544
rect 14884 14504 15384 14532
rect 14884 14492 14890 14504
rect 15378 14492 15384 14504
rect 15436 14532 15442 14544
rect 15764 14532 15792 14572
rect 16209 14569 16221 14603
rect 16255 14600 16267 14603
rect 16298 14600 16304 14612
rect 16255 14572 16304 14600
rect 16255 14569 16267 14572
rect 16209 14563 16267 14569
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 16485 14603 16543 14609
rect 16485 14569 16497 14603
rect 16531 14600 16543 14603
rect 16574 14600 16580 14612
rect 16531 14572 16580 14600
rect 16531 14569 16543 14572
rect 16485 14563 16543 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 16945 14603 17003 14609
rect 16945 14569 16957 14603
rect 16991 14600 17003 14603
rect 17218 14600 17224 14612
rect 16991 14572 17224 14600
rect 16991 14569 17003 14572
rect 16945 14563 17003 14569
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 17402 14560 17408 14612
rect 17460 14560 17466 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 18104 14572 18153 14600
rect 18104 14560 18110 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 18141 14563 18199 14569
rect 19334 14560 19340 14612
rect 19392 14560 19398 14612
rect 19429 14603 19487 14609
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 19518 14600 19524 14612
rect 19475 14572 19524 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 20990 14600 20996 14612
rect 19843 14572 20996 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 21324 14572 21465 14600
rect 21324 14560 21330 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 21453 14563 21511 14569
rect 21910 14560 21916 14612
rect 21968 14560 21974 14612
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 23845 14603 23903 14609
rect 23845 14600 23857 14603
rect 22428 14572 23857 14600
rect 22428 14560 22434 14572
rect 23845 14569 23857 14572
rect 23891 14569 23903 14603
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 23845 14563 23903 14569
rect 24136 14572 24593 14600
rect 17034 14532 17040 14544
rect 15436 14504 15607 14532
rect 15436 14492 15442 14504
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15470 14464 15476 14476
rect 15068 14436 15476 14464
rect 15068 14424 15074 14436
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15579 14473 15607 14504
rect 15764 14504 17040 14532
rect 15564 14467 15622 14473
rect 15564 14433 15576 14467
rect 15610 14433 15622 14467
rect 15564 14427 15622 14433
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 15764 14473 15792 14504
rect 16132 14473 16160 14504
rect 17034 14492 17040 14504
rect 17092 14492 17098 14544
rect 17420 14532 17448 14560
rect 17957 14535 18015 14541
rect 17144 14504 17356 14532
rect 17420 14504 17908 14532
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14433 16359 14467
rect 17144 14464 17172 14504
rect 16301 14427 16359 14433
rect 16592 14436 17172 14464
rect 17328 14464 17356 14504
rect 17880 14473 17908 14504
rect 17957 14501 17969 14535
rect 18003 14532 18015 14535
rect 18417 14535 18475 14541
rect 18417 14532 18429 14535
rect 18003 14504 18429 14532
rect 18003 14501 18015 14504
rect 17957 14495 18015 14501
rect 18417 14501 18429 14504
rect 18463 14532 18475 14535
rect 18463 14504 19472 14532
rect 18463 14501 18475 14504
rect 18417 14495 18475 14501
rect 19444 14476 19472 14504
rect 19978 14492 19984 14544
rect 20036 14532 20042 14544
rect 23474 14532 23480 14544
rect 20036 14504 23480 14532
rect 20036 14492 20042 14504
rect 23474 14492 23480 14504
rect 23532 14492 23538 14544
rect 17405 14467 17463 14473
rect 17405 14464 17417 14467
rect 17328 14436 17417 14464
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 12299 14300 13584 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 11664 14232 12204 14260
rect 11664 14220 11670 14232
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13740 14260 13768 14359
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14424 14368 15117 14396
rect 14424 14356 14430 14368
rect 15105 14365 15117 14368
rect 15151 14396 15163 14399
rect 15948 14396 15976 14427
rect 16316 14396 16344 14427
rect 16592 14408 16620 14436
rect 17405 14433 17417 14436
rect 17451 14433 17463 14467
rect 17405 14427 17463 14433
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 18046 14424 18052 14476
rect 18104 14424 18110 14476
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 18509 14467 18567 14473
rect 18509 14433 18521 14467
rect 18555 14433 18567 14467
rect 18509 14427 18567 14433
rect 16574 14396 16580 14408
rect 15151 14368 16580 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 15289 14331 15347 14337
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 16482 14328 16488 14340
rect 15335 14300 16488 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 13504 14232 13768 14260
rect 13504 14220 13510 14232
rect 14090 14220 14096 14272
rect 14148 14220 14154 14272
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 17052 14260 17080 14359
rect 17126 14356 17132 14408
rect 17184 14356 17190 14408
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 17236 14328 17264 14359
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 18230 14396 18236 14408
rect 17368 14368 18236 14396
rect 17368 14356 17374 14368
rect 18230 14356 18236 14368
rect 18288 14396 18294 14408
rect 18340 14396 18368 14427
rect 18414 14396 18420 14408
rect 18288 14368 18420 14396
rect 18288 14356 18294 14368
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 17144 14300 17264 14328
rect 17589 14331 17647 14337
rect 17144 14272 17172 14300
rect 17589 14297 17601 14331
rect 17635 14297 17647 14331
rect 17589 14291 17647 14297
rect 16448 14232 17080 14260
rect 16448 14220 16454 14232
rect 17126 14220 17132 14272
rect 17184 14220 17190 14272
rect 17604 14260 17632 14291
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18524 14328 18552 14427
rect 18598 14424 18604 14476
rect 18656 14473 18662 14476
rect 18656 14467 18705 14473
rect 18656 14433 18659 14467
rect 18693 14464 18705 14467
rect 19242 14464 19248 14476
rect 18693 14436 19248 14464
rect 18693 14433 18705 14436
rect 18656 14427 18705 14433
rect 18656 14424 18662 14427
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19426 14424 19432 14476
rect 19484 14424 19490 14476
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 19794 14464 19800 14476
rect 19567 14436 19800 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 20438 14464 20444 14476
rect 19896 14436 20444 14464
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 18966 14396 18972 14408
rect 18840 14368 18972 14396
rect 18840 14356 18846 14368
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 19058 14356 19064 14408
rect 19116 14356 19122 14408
rect 19153 14399 19211 14405
rect 19153 14365 19165 14399
rect 19199 14396 19211 14399
rect 19334 14396 19340 14408
rect 19199 14368 19340 14396
rect 19199 14365 19211 14368
rect 19153 14359 19211 14365
rect 19334 14356 19340 14368
rect 19392 14396 19398 14408
rect 19896 14396 19924 14436
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14464 20591 14467
rect 22922 14464 22928 14476
rect 20579 14436 22928 14464
rect 20579 14433 20591 14436
rect 20533 14427 20591 14433
rect 22922 14424 22928 14436
rect 22980 14464 22986 14476
rect 23382 14464 23388 14476
rect 22980 14436 23388 14464
rect 22980 14424 22986 14436
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 24136 14473 24164 14572
rect 24581 14569 24593 14572
rect 24627 14600 24639 14603
rect 24670 14600 24676 14612
rect 24627 14572 24676 14600
rect 24627 14569 24639 14572
rect 24581 14563 24639 14569
rect 24670 14560 24676 14572
rect 24728 14600 24734 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 24728 14572 25237 14600
rect 24728 14560 24734 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 26234 14600 26240 14612
rect 25225 14563 25283 14569
rect 25976 14572 26240 14600
rect 24228 14504 24808 14532
rect 24121 14467 24179 14473
rect 24121 14464 24133 14467
rect 23900 14436 24133 14464
rect 23900 14424 23906 14436
rect 24121 14433 24133 14436
rect 24167 14433 24179 14467
rect 24121 14427 24179 14433
rect 20162 14396 20168 14408
rect 19392 14368 19924 14396
rect 20088 14368 20168 14396
rect 19392 14356 19398 14368
rect 20088 14328 20116 14368
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 20404 14368 20637 14396
rect 20404 14356 20410 14368
rect 20625 14365 20637 14368
rect 20671 14396 20683 14399
rect 21358 14396 21364 14408
rect 20671 14368 21364 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 21542 14356 21548 14408
rect 21600 14396 21606 14408
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21600 14368 21649 14396
rect 21600 14356 21606 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 18012 14300 20116 14328
rect 18012 14288 18018 14300
rect 20438 14288 20444 14340
rect 20496 14328 20502 14340
rect 22020 14328 22048 14359
rect 22094 14356 22100 14408
rect 22152 14356 22158 14408
rect 23014 14356 23020 14408
rect 23072 14396 23078 14408
rect 23753 14399 23811 14405
rect 23753 14396 23765 14399
rect 23072 14368 23765 14396
rect 23072 14356 23078 14368
rect 23753 14365 23765 14368
rect 23799 14396 23811 14399
rect 24228 14396 24256 14504
rect 24780 14476 24808 14504
rect 24854 14492 24860 14544
rect 24912 14532 24918 14544
rect 24949 14535 25007 14541
rect 24949 14532 24961 14535
rect 24912 14504 24961 14532
rect 24912 14492 24918 14504
rect 24949 14501 24961 14504
rect 24995 14532 25007 14535
rect 25774 14532 25780 14544
rect 24995 14504 25780 14532
rect 24995 14501 25007 14504
rect 24949 14495 25007 14501
rect 25774 14492 25780 14504
rect 25832 14492 25838 14544
rect 24489 14467 24547 14473
rect 24489 14433 24501 14467
rect 24535 14433 24547 14467
rect 24489 14427 24547 14433
rect 23799 14368 24256 14396
rect 24305 14399 24363 14405
rect 23799 14365 23811 14368
rect 23753 14359 23811 14365
rect 24305 14365 24317 14399
rect 24351 14396 24363 14399
rect 24504 14396 24532 14427
rect 24762 14424 24768 14476
rect 24820 14424 24826 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 25148 14396 25176 14427
rect 25222 14424 25228 14476
rect 25280 14464 25286 14476
rect 25409 14467 25467 14473
rect 25409 14464 25421 14467
rect 25280 14436 25421 14464
rect 25280 14424 25286 14436
rect 25409 14433 25421 14436
rect 25455 14433 25467 14467
rect 25409 14427 25467 14433
rect 25866 14424 25872 14476
rect 25924 14424 25930 14476
rect 25976 14473 26004 14572
rect 26234 14560 26240 14572
rect 26292 14560 26298 14612
rect 26605 14603 26663 14609
rect 26605 14569 26617 14603
rect 26651 14600 26663 14603
rect 26694 14600 26700 14612
rect 26651 14572 26700 14600
rect 26651 14569 26663 14572
rect 26605 14563 26663 14569
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 27154 14560 27160 14612
rect 27212 14600 27218 14612
rect 28258 14600 28264 14612
rect 27212 14572 28264 14600
rect 27212 14560 27218 14572
rect 27430 14532 27436 14544
rect 26252 14504 27436 14532
rect 26252 14473 26280 14504
rect 27430 14492 27436 14504
rect 27488 14532 27494 14544
rect 27488 14504 27660 14532
rect 27488 14492 27494 14504
rect 25961 14467 26019 14473
rect 25961 14433 25973 14467
rect 26007 14433 26019 14467
rect 25961 14427 26019 14433
rect 26237 14467 26295 14473
rect 26237 14433 26249 14467
rect 26283 14433 26295 14467
rect 26237 14427 26295 14433
rect 25976 14396 26004 14427
rect 26602 14424 26608 14476
rect 26660 14424 26666 14476
rect 26786 14424 26792 14476
rect 26844 14424 26850 14476
rect 27632 14473 27660 14504
rect 27724 14473 27752 14572
rect 28258 14560 28264 14572
rect 28316 14560 28322 14612
rect 29822 14560 29828 14612
rect 29880 14600 29886 14612
rect 30009 14603 30067 14609
rect 30009 14600 30021 14603
rect 29880 14572 30021 14600
rect 29880 14560 29886 14572
rect 30009 14569 30021 14572
rect 30055 14569 30067 14603
rect 30009 14563 30067 14569
rect 30098 14560 30104 14612
rect 30156 14600 30162 14612
rect 30466 14600 30472 14612
rect 30156 14572 30472 14600
rect 30156 14560 30162 14572
rect 30466 14560 30472 14572
rect 30524 14600 30530 14612
rect 30926 14600 30932 14612
rect 30524 14572 30932 14600
rect 30524 14560 30530 14572
rect 30926 14560 30932 14572
rect 30984 14560 30990 14612
rect 31021 14603 31079 14609
rect 31021 14569 31033 14603
rect 31067 14600 31079 14603
rect 31110 14600 31116 14612
rect 31067 14572 31116 14600
rect 31067 14569 31079 14572
rect 31021 14563 31079 14569
rect 31110 14560 31116 14572
rect 31168 14560 31174 14612
rect 28276 14532 28304 14560
rect 30374 14532 30380 14544
rect 28276 14504 30380 14532
rect 27617 14467 27675 14473
rect 27617 14433 27629 14467
rect 27663 14433 27675 14467
rect 27617 14427 27675 14433
rect 27709 14467 27767 14473
rect 27709 14433 27721 14467
rect 27755 14433 27767 14467
rect 27709 14427 27767 14433
rect 27893 14467 27951 14473
rect 27893 14433 27905 14467
rect 27939 14433 27951 14467
rect 27893 14427 27951 14433
rect 27985 14467 28043 14473
rect 27985 14433 27997 14467
rect 28031 14464 28043 14467
rect 28534 14464 28540 14476
rect 28031 14436 28540 14464
rect 28031 14433 28043 14436
rect 27985 14427 28043 14433
rect 24351 14368 25176 14396
rect 25884 14368 26004 14396
rect 26053 14399 26111 14405
rect 24351 14365 24363 14368
rect 24305 14359 24363 14365
rect 22462 14328 22468 14340
rect 20496 14300 22468 14328
rect 20496 14288 20502 14300
rect 22462 14288 22468 14300
rect 22520 14328 22526 14340
rect 23934 14328 23940 14340
rect 22520 14300 23940 14328
rect 22520 14288 22526 14300
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 24026 14288 24032 14340
rect 24084 14328 24090 14340
rect 24320 14328 24348 14359
rect 25884 14340 25912 14368
rect 26053 14365 26065 14399
rect 26099 14396 26111 14399
rect 26620 14396 26648 14424
rect 26099 14368 26648 14396
rect 27065 14399 27123 14405
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 27065 14365 27077 14399
rect 27111 14365 27123 14399
rect 27908 14396 27936 14427
rect 28534 14424 28540 14436
rect 28592 14424 28598 14476
rect 28644 14473 28672 14504
rect 30374 14492 30380 14504
rect 30432 14532 30438 14544
rect 30745 14535 30803 14541
rect 30745 14532 30757 14535
rect 30432 14504 30757 14532
rect 30432 14492 30438 14504
rect 30745 14501 30757 14504
rect 30791 14501 30803 14535
rect 30745 14495 30803 14501
rect 28629 14467 28687 14473
rect 28629 14433 28641 14467
rect 28675 14433 28687 14467
rect 28629 14427 28687 14433
rect 28718 14424 28724 14476
rect 28776 14464 28782 14476
rect 28813 14467 28871 14473
rect 28813 14464 28825 14467
rect 28776 14436 28825 14464
rect 28776 14424 28782 14436
rect 28813 14433 28825 14436
rect 28859 14464 28871 14467
rect 29086 14464 29092 14476
rect 28859 14436 29092 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 29638 14424 29644 14476
rect 29696 14464 29702 14476
rect 29733 14467 29791 14473
rect 29733 14464 29745 14467
rect 29696 14436 29745 14464
rect 29696 14424 29702 14436
rect 29733 14433 29745 14436
rect 29779 14433 29791 14467
rect 29733 14427 29791 14433
rect 29917 14467 29975 14473
rect 29917 14433 29929 14467
rect 29963 14464 29975 14467
rect 30006 14464 30012 14476
rect 29963 14436 30012 14464
rect 29963 14433 29975 14436
rect 29917 14427 29975 14433
rect 30006 14424 30012 14436
rect 30064 14464 30070 14476
rect 30469 14467 30527 14473
rect 30469 14464 30481 14467
rect 30064 14436 30481 14464
rect 30064 14424 30070 14436
rect 30469 14433 30481 14436
rect 30515 14433 30527 14467
rect 30469 14427 30527 14433
rect 30834 14424 30840 14476
rect 30892 14424 30898 14476
rect 31018 14424 31024 14476
rect 31076 14424 31082 14476
rect 27908 14368 28028 14396
rect 27065 14359 27123 14365
rect 24084 14300 24348 14328
rect 24084 14288 24090 14300
rect 25866 14288 25872 14340
rect 25924 14288 25930 14340
rect 26237 14331 26295 14337
rect 26237 14297 26249 14331
rect 26283 14328 26295 14331
rect 27080 14328 27108 14359
rect 26283 14300 27108 14328
rect 26283 14297 26295 14300
rect 26237 14291 26295 14297
rect 28000 14272 28028 14368
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 30193 14399 30251 14405
rect 30193 14396 30205 14399
rect 30156 14368 30205 14396
rect 30156 14356 30162 14368
rect 30193 14365 30205 14368
rect 30239 14365 30251 14399
rect 30193 14359 30251 14365
rect 30285 14399 30343 14405
rect 30285 14365 30297 14399
rect 30331 14365 30343 14399
rect 30285 14359 30343 14365
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30852 14396 30880 14424
rect 30423 14368 30880 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 30300 14328 30328 14359
rect 31036 14328 31064 14424
rect 30300 14300 31064 14328
rect 30392 14272 30420 14300
rect 19150 14260 19156 14272
rect 17604 14232 19156 14260
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 20533 14263 20591 14269
rect 20533 14260 20545 14263
rect 19300 14232 20545 14260
rect 19300 14220 19306 14232
rect 20533 14229 20545 14232
rect 20579 14260 20591 14263
rect 20622 14260 20628 14272
rect 20579 14232 20628 14260
rect 20579 14229 20591 14232
rect 20533 14223 20591 14229
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21174 14260 21180 14272
rect 20947 14232 21180 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 23198 14260 23204 14272
rect 22888 14232 23204 14260
rect 22888 14220 22894 14232
rect 23198 14220 23204 14232
rect 23256 14260 23262 14272
rect 24854 14260 24860 14272
rect 23256 14232 24860 14260
rect 23256 14220 23262 14232
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 25409 14263 25467 14269
rect 25409 14229 25421 14263
rect 25455 14260 25467 14263
rect 26878 14260 26884 14272
rect 25455 14232 26884 14260
rect 25455 14229 25467 14232
rect 25409 14223 25467 14229
rect 26878 14220 26884 14232
rect 26936 14220 26942 14272
rect 26973 14263 27031 14269
rect 26973 14229 26985 14263
rect 27019 14260 27031 14263
rect 27433 14263 27491 14269
rect 27433 14260 27445 14263
rect 27019 14232 27445 14260
rect 27019 14229 27031 14232
rect 26973 14223 27031 14229
rect 27433 14229 27445 14232
rect 27479 14229 27491 14263
rect 27433 14223 27491 14229
rect 27982 14220 27988 14272
rect 28040 14220 28046 14272
rect 29822 14220 29828 14272
rect 29880 14220 29886 14272
rect 30374 14220 30380 14272
rect 30432 14220 30438 14272
rect 552 14170 31648 14192
rect 552 14118 4285 14170
rect 4337 14118 4349 14170
rect 4401 14118 4413 14170
rect 4465 14118 4477 14170
rect 4529 14118 4541 14170
rect 4593 14118 12059 14170
rect 12111 14118 12123 14170
rect 12175 14118 12187 14170
rect 12239 14118 12251 14170
rect 12303 14118 12315 14170
rect 12367 14118 19833 14170
rect 19885 14118 19897 14170
rect 19949 14118 19961 14170
rect 20013 14118 20025 14170
rect 20077 14118 20089 14170
rect 20141 14118 27607 14170
rect 27659 14118 27671 14170
rect 27723 14118 27735 14170
rect 27787 14118 27799 14170
rect 27851 14118 27863 14170
rect 27915 14118 31648 14170
rect 552 14096 31648 14118
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3283 14059 3341 14065
rect 3283 14056 3295 14059
rect 2832 14028 3295 14056
rect 2832 14016 2838 14028
rect 3283 14025 3295 14028
rect 3329 14056 3341 14059
rect 3418 14056 3424 14068
rect 3329 14028 3424 14056
rect 3329 14025 3341 14028
rect 3283 14019 3341 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 4154 14056 4160 14068
rect 3568 14028 4160 14056
rect 3568 14016 3574 14028
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4890 14016 4896 14068
rect 4948 14056 4954 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 4948 14028 5181 14056
rect 4948 14016 4954 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 10413 14059 10471 14065
rect 5408 14028 10180 14056
rect 5408 14016 5414 14028
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13957 3111 13991
rect 3053 13951 3111 13957
rect 3068 13920 3096 13951
rect 8294 13948 8300 14000
rect 8352 13988 8358 14000
rect 9490 13988 9496 14000
rect 8352 13960 9496 13988
rect 8352 13948 8358 13960
rect 9490 13948 9496 13960
rect 9548 13988 9554 14000
rect 9858 13988 9864 14000
rect 9548 13960 9864 13988
rect 9548 13948 9554 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 4709 13923 4767 13929
rect 4709 13920 4721 13923
rect 3068 13892 4721 13920
rect 4709 13889 4721 13892
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5534 13920 5540 13932
rect 5123 13892 5540 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5534 13880 5540 13892
rect 5592 13920 5598 13932
rect 6362 13920 6368 13932
rect 5592 13892 6368 13920
rect 5592 13880 5598 13892
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 7524 13892 8033 13920
rect 7524 13880 7530 13892
rect 8021 13889 8033 13892
rect 8067 13889 8079 13923
rect 8938 13920 8944 13932
rect 8021 13883 8079 13889
rect 8404 13892 8944 13920
rect 845 13855 903 13861
rect 845 13821 857 13855
rect 891 13852 903 13855
rect 934 13852 940 13864
rect 891 13824 940 13852
rect 891 13821 903 13824
rect 845 13815 903 13821
rect 934 13812 940 13824
rect 992 13812 998 13864
rect 1210 13812 1216 13864
rect 1268 13812 1274 13864
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 5224 13824 5365 13852
rect 5224 13812 5230 13824
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 2222 13744 2228 13796
rect 2280 13744 2286 13796
rect 4370 13756 4476 13784
rect 2639 13719 2697 13725
rect 2639 13685 2651 13719
rect 2685 13716 2697 13719
rect 2774 13716 2780 13728
rect 2685 13688 2780 13716
rect 2685 13685 2697 13688
rect 2639 13679 2697 13685
rect 2774 13676 2780 13688
rect 2832 13716 2838 13728
rect 3878 13716 3884 13728
rect 2832 13688 3884 13716
rect 2832 13676 2838 13688
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 4448 13716 4476 13756
rect 5810 13744 5816 13796
rect 5868 13744 5874 13796
rect 7837 13787 7895 13793
rect 7300 13756 7604 13784
rect 4706 13716 4712 13728
rect 4448 13688 4712 13716
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 7300 13725 7328 13756
rect 7576 13728 7604 13756
rect 7837 13753 7849 13787
rect 7883 13753 7895 13787
rect 8036 13784 8064 13883
rect 8404 13861 8432 13892
rect 8938 13880 8944 13892
rect 8996 13920 9002 13932
rect 8996 13892 9628 13920
rect 8996 13880 9002 13892
rect 9600 13864 9628 13892
rect 9674 13880 9680 13932
rect 9732 13880 9738 13932
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8757 13855 8815 13861
rect 8757 13852 8769 13855
rect 8628 13824 8769 13852
rect 8628 13812 8634 13824
rect 8757 13821 8769 13824
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9398 13852 9404 13864
rect 9263 13824 9404 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 9582 13812 9588 13864
rect 9640 13812 9646 13864
rect 9692 13852 9720 13880
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9692 13824 9781 13852
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 9862 13855 9920 13861
rect 9862 13821 9874 13855
rect 9908 13846 9920 13855
rect 9950 13846 9956 13864
rect 9908 13821 9956 13846
rect 9862 13818 9956 13821
rect 9862 13815 9920 13818
rect 9950 13812 9956 13818
rect 10008 13812 10014 13864
rect 10152 13861 10180 14028
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 11146 14056 11152 14068
rect 10459 14028 11152 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11504 14059 11562 14065
rect 11504 14025 11516 14059
rect 11550 14056 11562 14059
rect 11882 14056 11888 14068
rect 11550 14028 11888 14056
rect 11550 14025 11562 14028
rect 11504 14019 11562 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 13446 14056 13452 14068
rect 12032 14028 13452 14056
rect 12032 14016 12038 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13817 14059 13875 14065
rect 13817 14025 13829 14059
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 14001 14059 14059 14065
rect 14001 14025 14013 14059
rect 14047 14056 14059 14059
rect 14182 14056 14188 14068
rect 14047 14028 14188 14056
rect 14047 14025 14059 14028
rect 14001 14019 14059 14025
rect 13832 13988 13860 14019
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14700 14028 14749 14056
rect 14700 14016 14706 14028
rect 14737 14025 14749 14028
rect 14783 14056 14795 14059
rect 15654 14056 15660 14068
rect 14783 14028 15660 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 17586 14056 17592 14068
rect 16724 14028 17592 14056
rect 16724 14016 16730 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 19334 14056 19340 14068
rect 17828 14028 19340 14056
rect 17828 14016 17834 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 20346 14056 20352 14068
rect 19843 14028 20352 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 20438 14016 20444 14068
rect 20496 14016 20502 14068
rect 20622 14016 20628 14068
rect 20680 14016 20686 14068
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 20772 14028 20821 14056
rect 20772 14016 20778 14028
rect 20809 14025 20821 14028
rect 20855 14025 20867 14059
rect 20809 14019 20867 14025
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 22649 14059 22707 14065
rect 22649 14056 22661 14059
rect 21784 14028 22661 14056
rect 21784 14016 21790 14028
rect 22649 14025 22661 14028
rect 22695 14025 22707 14059
rect 22649 14019 22707 14025
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23109 14059 23167 14065
rect 23109 14056 23121 14059
rect 22796 14028 23121 14056
rect 22796 14016 22802 14028
rect 23109 14025 23121 14028
rect 23155 14056 23167 14059
rect 23842 14056 23848 14068
rect 23155 14028 23848 14056
rect 23155 14025 23167 14028
rect 23109 14019 23167 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 24394 14016 24400 14068
rect 24452 14016 24458 14068
rect 24596 14028 25912 14056
rect 24596 14000 24624 14028
rect 13832 13960 14228 13988
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13920 11299 13923
rect 11514 13920 11520 13932
rect 11287 13892 11520 13920
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 13044 13892 13277 13920
rect 13044 13880 13050 13892
rect 13265 13889 13277 13892
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 14200 13864 14228 13960
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 21542 13988 21548 14000
rect 17920 13960 21548 13988
rect 17920 13948 17926 13960
rect 21542 13948 21548 13960
rect 21600 13988 21606 14000
rect 24486 13988 24492 14000
rect 21600 13960 24492 13988
rect 21600 13948 21606 13960
rect 24486 13948 24492 13960
rect 24544 13948 24550 14000
rect 24578 13948 24584 14000
rect 24636 13948 24642 14000
rect 24854 13948 24860 14000
rect 24912 13988 24918 14000
rect 24912 13960 25544 13988
rect 24912 13948 24918 13960
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15378 13920 15384 13932
rect 14875 13892 15384 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15378 13880 15384 13892
rect 15436 13920 15442 13932
rect 15436 13892 17080 13920
rect 15436 13880 15442 13892
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 10275 13855 10333 13861
rect 10275 13821 10287 13855
rect 10321 13852 10333 13855
rect 10410 13852 10416 13864
rect 10321 13824 10416 13852
rect 10321 13821 10333 13824
rect 10275 13815 10333 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10778 13852 10784 13864
rect 10735 13824 10784 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 8665 13787 8723 13793
rect 8665 13784 8677 13787
rect 8036 13756 8677 13784
rect 7837 13747 7895 13753
rect 8665 13753 8677 13756
rect 8711 13753 8723 13787
rect 9140 13784 9168 13812
rect 9309 13787 9367 13793
rect 9309 13784 9321 13787
rect 9140 13756 9321 13784
rect 8665 13747 8723 13753
rect 9309 13753 9321 13756
rect 9355 13753 9367 13787
rect 9309 13747 9367 13753
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 10045 13787 10103 13793
rect 10045 13784 10057 13787
rect 9723 13756 10057 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 10045 13753 10057 13756
rect 10091 13753 10103 13787
rect 10980 13784 11008 13815
rect 13170 13812 13176 13864
rect 13228 13852 13234 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13228 13824 13553 13852
rect 13228 13812 13234 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 13725 13855 13783 13861
rect 13725 13821 13737 13855
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13852 13875 13855
rect 13998 13852 14004 13864
rect 13863 13824 14004 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 11974 13784 11980 13796
rect 10045 13747 10103 13753
rect 10428 13756 11008 13784
rect 11072 13756 11980 13784
rect 7285 13719 7343 13725
rect 7285 13685 7297 13719
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 7374 13676 7380 13728
rect 7432 13676 7438 13728
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 7745 13719 7803 13725
rect 7745 13716 7757 13719
rect 7616 13688 7757 13716
rect 7616 13676 7622 13688
rect 7745 13685 7757 13688
rect 7791 13685 7803 13719
rect 7852 13716 7880 13747
rect 10428 13728 10456 13756
rect 7926 13716 7932 13728
rect 7852 13688 7932 13716
rect 7745 13679 7803 13685
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 10318 13716 10324 13728
rect 9180 13688 10324 13716
rect 9180 13676 9186 13688
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10410 13676 10416 13728
rect 10468 13676 10474 13728
rect 10502 13676 10508 13728
rect 10560 13676 10566 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10836 13688 10885 13716
rect 10836 13676 10842 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11072 13716 11100 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 11020 13688 11100 13716
rect 11020 13676 11026 13688
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 13740 13716 13768 13815
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 14367 13855 14425 13861
rect 14367 13821 14379 13855
rect 14413 13852 14425 13855
rect 15010 13852 15016 13864
rect 14413 13824 15016 13852
rect 14413 13821 14425 13824
rect 14367 13815 14425 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15654 13812 15660 13864
rect 15712 13812 15718 13864
rect 16942 13812 16948 13864
rect 17000 13812 17006 13864
rect 17052 13861 17080 13892
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 17184 13892 17969 13920
rect 17184 13880 17190 13892
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 22002 13920 22008 13932
rect 19024 13892 22008 13920
rect 19024 13880 19030 13892
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 25516 13920 25544 13960
rect 25884 13920 25912 14028
rect 27430 14016 27436 14068
rect 27488 14016 27494 14068
rect 30558 14016 30564 14068
rect 30616 14016 30622 14068
rect 27985 13923 28043 13929
rect 27985 13920 27997 13923
rect 22112 13892 24256 13920
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 15194 13784 15200 13796
rect 14516 13756 15200 13784
rect 14516 13744 14522 13756
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 15672 13784 15700 13812
rect 17604 13784 17632 13815
rect 17678 13812 17684 13864
rect 17736 13852 17742 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17736 13824 17785 13852
rect 17736 13812 17742 13824
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 18230 13812 18236 13864
rect 18288 13812 18294 13864
rect 19334 13812 19340 13864
rect 19392 13812 19398 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19484 13824 19533 13852
rect 19484 13812 19490 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 21634 13852 21640 13864
rect 19521 13815 19579 13821
rect 20916 13824 21640 13852
rect 15528 13756 17632 13784
rect 15528 13744 15534 13756
rect 13814 13716 13820 13728
rect 11296 13688 13820 13716
rect 11296 13676 11302 13688
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 14148 13688 14197 13716
rect 14148 13676 14154 13688
rect 14185 13685 14197 13688
rect 14231 13685 14243 13719
rect 14185 13679 14243 13685
rect 14366 13676 14372 13728
rect 14424 13676 14430 13728
rect 15654 13676 15660 13728
rect 15712 13676 15718 13728
rect 17604 13716 17632 13756
rect 20162 13744 20168 13796
rect 20220 13744 20226 13796
rect 20793 13787 20851 13793
rect 20793 13753 20805 13787
rect 20839 13784 20851 13787
rect 20916 13784 20944 13824
rect 21634 13812 21640 13824
rect 21692 13852 21698 13864
rect 22112 13861 22140 13892
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 21692 13824 22109 13852
rect 21692 13812 21698 13824
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 22517 13855 22575 13861
rect 22517 13821 22529 13855
rect 22563 13852 22575 13855
rect 22646 13852 22652 13864
rect 22563 13824 22652 13852
rect 22563 13821 22575 13824
rect 22517 13815 22575 13821
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 22833 13855 22891 13861
rect 22833 13821 22845 13855
rect 22879 13852 22891 13855
rect 22922 13852 22928 13864
rect 22879 13824 22928 13852
rect 22879 13821 22891 13824
rect 22833 13815 22891 13821
rect 22922 13812 22928 13824
rect 22980 13812 22986 13864
rect 23032 13824 23428 13852
rect 20839 13756 20944 13784
rect 20839 13753 20851 13756
rect 20793 13747 20851 13753
rect 20990 13744 20996 13796
rect 21048 13744 21054 13796
rect 21542 13744 21548 13796
rect 21600 13784 21606 13796
rect 22281 13787 22339 13793
rect 22281 13784 22293 13787
rect 21600 13756 22293 13784
rect 21600 13744 21606 13756
rect 22281 13753 22293 13756
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 22373 13787 22431 13793
rect 22373 13753 22385 13787
rect 22419 13784 22431 13787
rect 22738 13784 22744 13796
rect 22419 13756 22744 13784
rect 22419 13753 22431 13756
rect 22373 13747 22431 13753
rect 18506 13716 18512 13728
rect 17604 13688 18512 13716
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 20180 13716 20208 13744
rect 20898 13716 20904 13728
rect 20180 13688 20904 13716
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 22296 13716 22324 13747
rect 22738 13744 22744 13756
rect 22796 13744 22802 13796
rect 23032 13716 23060 13824
rect 23198 13744 23204 13796
rect 23256 13784 23262 13796
rect 23293 13787 23351 13793
rect 23293 13784 23305 13787
rect 23256 13756 23305 13784
rect 23256 13744 23262 13756
rect 23293 13753 23305 13756
rect 23339 13753 23351 13787
rect 23400 13784 23428 13824
rect 23842 13812 23848 13864
rect 23900 13812 23906 13864
rect 24228 13861 24256 13892
rect 24596 13892 25452 13920
rect 25516 13892 25820 13920
rect 25884 13892 27997 13920
rect 24596 13861 24624 13892
rect 25424 13864 25452 13892
rect 24213 13855 24271 13861
rect 24213 13821 24225 13855
rect 24259 13852 24271 13855
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24259 13824 24593 13852
rect 24259 13821 24271 13824
rect 24213 13815 24271 13821
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 24762 13812 24768 13864
rect 24820 13852 24826 13864
rect 24857 13855 24915 13861
rect 24857 13852 24869 13855
rect 24820 13824 24869 13852
rect 24820 13812 24826 13824
rect 24857 13821 24869 13824
rect 24903 13821 24915 13855
rect 24857 13815 24915 13821
rect 25406 13812 25412 13864
rect 25464 13812 25470 13864
rect 25792 13861 25820 13892
rect 27985 13889 27997 13892
rect 28031 13920 28043 13923
rect 28258 13920 28264 13932
rect 28031 13892 28264 13920
rect 28031 13889 28043 13892
rect 27985 13883 28043 13889
rect 28258 13880 28264 13892
rect 28316 13920 28322 13932
rect 28626 13920 28632 13932
rect 28316 13892 28632 13920
rect 28316 13880 28322 13892
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 30576 13920 30604 14016
rect 28966 13892 30604 13920
rect 25593 13855 25651 13861
rect 25593 13852 25605 13855
rect 25516 13824 25605 13852
rect 24121 13787 24179 13793
rect 24121 13784 24133 13787
rect 23400 13756 24133 13784
rect 23293 13747 23351 13753
rect 24121 13753 24133 13756
rect 24167 13753 24179 13787
rect 24121 13747 24179 13753
rect 22296 13688 23060 13716
rect 23109 13719 23167 13725
rect 23109 13685 23121 13719
rect 23155 13716 23167 13719
rect 23566 13716 23572 13728
rect 23155 13688 23572 13716
rect 23155 13685 23167 13688
rect 23109 13679 23167 13685
rect 23566 13676 23572 13688
rect 23624 13716 23630 13728
rect 24026 13716 24032 13728
rect 23624 13688 24032 13716
rect 23624 13676 23630 13688
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24136 13716 24164 13747
rect 24394 13744 24400 13796
rect 24452 13784 24458 13796
rect 25041 13787 25099 13793
rect 25041 13784 25053 13787
rect 24452 13756 25053 13784
rect 24452 13744 24458 13756
rect 25041 13753 25053 13756
rect 25087 13784 25099 13787
rect 25222 13784 25228 13796
rect 25087 13756 25228 13784
rect 25087 13753 25099 13756
rect 25041 13747 25099 13753
rect 25222 13744 25228 13756
rect 25280 13744 25286 13796
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 24136 13688 24685 13716
rect 24673 13685 24685 13688
rect 24719 13716 24731 13719
rect 24854 13716 24860 13728
rect 24719 13688 24860 13716
rect 24719 13685 24731 13688
rect 24673 13679 24731 13685
rect 24854 13676 24860 13688
rect 24912 13716 24918 13728
rect 25516 13716 25544 13824
rect 25593 13821 25605 13824
rect 25639 13821 25651 13855
rect 25593 13815 25651 13821
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13852 25835 13855
rect 28966 13852 28994 13892
rect 25823 13824 28994 13852
rect 25823 13821 25835 13824
rect 25777 13815 25835 13821
rect 30190 13812 30196 13864
rect 30248 13812 30254 13864
rect 30374 13812 30380 13864
rect 30432 13852 30438 13864
rect 30469 13855 30527 13861
rect 30469 13852 30481 13855
rect 30432 13824 30481 13852
rect 30432 13812 30438 13824
rect 30469 13821 30481 13824
rect 30515 13821 30527 13855
rect 30469 13815 30527 13821
rect 26510 13744 26516 13796
rect 26568 13744 26574 13796
rect 26694 13744 26700 13796
rect 26752 13784 26758 13796
rect 27801 13787 27859 13793
rect 27801 13784 27813 13787
rect 26752 13756 27813 13784
rect 26752 13744 26758 13756
rect 27801 13753 27813 13756
rect 27847 13784 27859 13787
rect 28350 13784 28356 13796
rect 27847 13756 28356 13784
rect 27847 13753 27859 13756
rect 27801 13747 27859 13753
rect 28350 13744 28356 13756
rect 28408 13744 28414 13796
rect 24912 13688 25544 13716
rect 26528 13716 26556 13744
rect 27062 13716 27068 13728
rect 26528 13688 27068 13716
rect 24912 13676 24918 13688
rect 27062 13676 27068 13688
rect 27120 13716 27126 13728
rect 27893 13719 27951 13725
rect 27893 13716 27905 13719
rect 27120 13688 27905 13716
rect 27120 13676 27126 13688
rect 27893 13685 27905 13688
rect 27939 13685 27951 13719
rect 27893 13679 27951 13685
rect 552 13626 31808 13648
rect 552 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 15946 13626
rect 15998 13574 16010 13626
rect 16062 13574 16074 13626
rect 16126 13574 16138 13626
rect 16190 13574 16202 13626
rect 16254 13574 23720 13626
rect 23772 13574 23784 13626
rect 23836 13574 23848 13626
rect 23900 13574 23912 13626
rect 23964 13574 23976 13626
rect 24028 13574 31494 13626
rect 31546 13574 31558 13626
rect 31610 13574 31622 13626
rect 31674 13574 31686 13626
rect 31738 13574 31750 13626
rect 31802 13574 31808 13626
rect 552 13552 31808 13574
rect 1210 13472 1216 13524
rect 1268 13472 1274 13524
rect 1857 13515 1915 13521
rect 1857 13481 1869 13515
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1872 13376 1900 13475
rect 2240 13444 2268 13475
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2924 13484 3065 13512
rect 2924 13472 2930 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 3418 13472 3424 13524
rect 3476 13472 3482 13524
rect 5534 13512 5540 13524
rect 3896 13484 5540 13512
rect 2774 13444 2780 13456
rect 2240 13416 2780 13444
rect 2774 13404 2780 13416
rect 2832 13404 2838 13456
rect 3068 13416 3556 13444
rect 1443 13348 1900 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 2188 13348 2329 13376
rect 2188 13336 2194 13348
rect 2317 13345 2329 13348
rect 2363 13376 2375 13379
rect 2958 13376 2964 13388
rect 2363 13348 2964 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2958 13336 2964 13348
rect 3016 13376 3022 13388
rect 3068 13376 3096 13416
rect 3528 13385 3556 13416
rect 3896 13385 3924 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5868 13484 6009 13512
rect 5868 13472 5874 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 8386 13512 8392 13524
rect 5997 13475 6055 13481
rect 6085 13484 8392 13512
rect 4706 13404 4712 13456
rect 4764 13404 4770 13456
rect 3016 13348 3096 13376
rect 3513 13379 3571 13385
rect 3016 13336 3022 13348
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 3881 13379 3939 13385
rect 3881 13345 3893 13379
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2682 13308 2688 13320
rect 2547 13280 2688 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3694 13268 3700 13320
rect 3752 13268 3758 13320
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 3896 13240 3924 13339
rect 4154 13268 4160 13320
rect 4212 13268 4218 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6085 13308 6113 13484
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 9293 13515 9351 13521
rect 9293 13481 9305 13515
rect 9339 13512 9351 13515
rect 9766 13512 9772 13524
rect 9339 13484 9772 13512
rect 9339 13481 9351 13484
rect 9293 13475 9351 13481
rect 9766 13472 9772 13484
rect 9824 13512 9830 13524
rect 10410 13512 10416 13524
rect 9824 13484 10416 13512
rect 9824 13472 9830 13484
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10686 13472 10692 13524
rect 10744 13472 10750 13524
rect 11517 13515 11575 13521
rect 11517 13481 11529 13515
rect 11563 13512 11575 13515
rect 12342 13512 12348 13524
rect 11563 13484 12348 13512
rect 11563 13481 11575 13484
rect 11517 13475 11575 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 18966 13512 18972 13524
rect 15764 13484 18552 13512
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 8665 13447 8723 13453
rect 6972 13416 7314 13444
rect 6972 13404 6978 13416
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 8754 13444 8760 13456
rect 8711 13416 8760 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 8849 13447 8907 13453
rect 8849 13413 8861 13447
rect 8895 13444 8907 13447
rect 9122 13444 9128 13456
rect 8895 13416 9128 13444
rect 8895 13413 8907 13416
rect 8849 13407 8907 13413
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 9490 13404 9496 13456
rect 9548 13404 9554 13456
rect 9861 13447 9919 13453
rect 9861 13413 9873 13447
rect 9907 13444 9919 13447
rect 10502 13444 10508 13456
rect 9907 13416 10508 13444
rect 9907 13413 9919 13416
rect 9861 13407 9919 13413
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 10704 13444 10732 13472
rect 12066 13444 12072 13456
rect 10617 13416 10732 13444
rect 11348 13416 12072 13444
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 5684 13280 6113 13308
rect 5684 13268 5690 13280
rect 992 13212 3924 13240
rect 992 13200 998 13212
rect 6196 13172 6224 13339
rect 6270 13336 6276 13388
rect 6328 13336 6334 13388
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6420 13348 6561 13376
rect 6420 13336 6426 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6472 13280 6837 13308
rect 6472 13249 6500 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13209 6515 13243
rect 8404 13240 8432 13339
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 9030 13336 9036 13388
rect 9088 13336 9094 13388
rect 9582 13336 9588 13388
rect 9640 13336 9646 13388
rect 9723 13379 9781 13385
rect 9723 13345 9735 13379
rect 9769 13345 9781 13379
rect 9723 13339 9781 13345
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8527 13280 9635 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8662 13240 8668 13252
rect 8404 13212 8668 13240
rect 6457 13203 6515 13209
rect 8662 13200 8668 13212
rect 8720 13240 8726 13252
rect 9030 13240 9036 13252
rect 8720 13212 9036 13240
rect 8720 13200 8726 13212
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 9125 13243 9183 13249
rect 9125 13209 9137 13243
rect 9171 13240 9183 13243
rect 9214 13240 9220 13252
rect 9171 13212 9220 13240
rect 9171 13209 9183 13212
rect 9125 13203 9183 13209
rect 7374 13172 7380 13184
rect 6196 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8478 13172 8484 13184
rect 8352 13144 8484 13172
rect 8352 13132 8358 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 9140 13172 9168 13203
rect 9214 13200 9220 13212
rect 9272 13200 9278 13252
rect 9607 13240 9635 13280
rect 9738 13240 9766 13339
rect 9968 13308 9996 13339
rect 10042 13336 10048 13388
rect 10100 13385 10106 13388
rect 10100 13376 10108 13385
rect 10100 13348 10145 13376
rect 10100 13339 10108 13348
rect 10100 13336 10106 13339
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10284 13348 10425 13376
rect 10284 13336 10290 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 10134 13308 10140 13320
rect 9968 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10617 13240 10645 13416
rect 11348 13388 11376 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 12308 13416 12466 13444
rect 12308 13404 12314 13416
rect 13446 13404 13452 13456
rect 13504 13444 13510 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13504 13416 13737 13444
rect 13504 13404 13510 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 15764 13444 15792 13484
rect 15620 13416 15792 13444
rect 16669 13447 16727 13453
rect 15620 13404 15626 13416
rect 16669 13413 16681 13447
rect 16715 13444 16727 13447
rect 16850 13444 16856 13456
rect 16715 13416 16856 13444
rect 16715 13413 16727 13416
rect 16669 13407 16727 13413
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 17034 13404 17040 13456
rect 17092 13453 17098 13456
rect 17092 13447 17141 13453
rect 17092 13413 17095 13447
rect 17129 13413 17141 13447
rect 18046 13444 18052 13456
rect 17092 13407 17141 13413
rect 17328 13416 18052 13444
rect 17092 13404 17098 13407
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10744 13348 11069 13376
rect 10744 13336 10750 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 11238 13336 11244 13388
rect 11296 13336 11302 13388
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 13596 13348 13860 13376
rect 13596 13336 13602 13348
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 11572 13280 11713 13308
rect 11572 13268 11578 13280
rect 11701 13277 11713 13280
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 9607 13212 9766 13240
rect 10153 13212 11560 13240
rect 8628 13144 9168 13172
rect 9309 13175 9367 13181
rect 8628 13132 8634 13144
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 10153 13172 10181 13212
rect 11532 13184 11560 13212
rect 9355 13144 10181 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 10226 13132 10232 13184
rect 10284 13132 10290 13184
rect 10502 13132 10508 13184
rect 10560 13132 10566 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11422 13172 11428 13184
rect 11379 13144 11428 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11514 13132 11520 13184
rect 11572 13132 11578 13184
rect 11716 13172 11744 13271
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 13832 13308 13860 13348
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14424 13348 14657 13376
rect 14424 13336 14430 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 15010 13336 15016 13388
rect 15068 13336 15074 13388
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 15197 13379 15255 13385
rect 15197 13376 15209 13379
rect 15160 13348 15209 13376
rect 15160 13336 15166 13348
rect 15197 13345 15209 13348
rect 15243 13376 15255 13379
rect 15378 13376 15384 13388
rect 15243 13348 15384 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15470 13336 15476 13388
rect 15528 13336 15534 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15896 13348 16313 13376
rect 15896 13336 15902 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 16206 13308 16212 13320
rect 12124 13280 13124 13308
rect 13832 13280 16212 13308
rect 12124 13268 12130 13280
rect 12986 13200 12992 13252
rect 13044 13200 13050 13252
rect 13096 13240 13124 13280
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16408 13308 16436 13339
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 17328 13385 17356 13416
rect 18046 13404 18052 13416
rect 18104 13444 18110 13456
rect 18104 13416 18184 13444
rect 18104 13404 18110 13416
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16632 13348 16957 13376
rect 16632 13336 16638 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17221 13379 17279 13385
rect 17221 13345 17233 13379
rect 17267 13345 17279 13379
rect 17221 13339 17279 13345
rect 17313 13379 17371 13385
rect 17313 13345 17325 13379
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 16408 13280 16712 13308
rect 16684 13252 16712 13280
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 13998 13240 14004 13252
rect 13096 13212 14004 13240
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 15105 13243 15163 13249
rect 15105 13240 15117 13243
rect 14976 13212 15117 13240
rect 14976 13200 14982 13212
rect 15105 13209 15117 13212
rect 15151 13209 15163 13243
rect 15105 13203 15163 13209
rect 15746 13200 15752 13252
rect 15804 13240 15810 13252
rect 15804 13212 16620 13240
rect 15804 13200 15810 13212
rect 11974 13172 11980 13184
rect 11716 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 13004 13172 13032 13200
rect 16117 13175 16175 13181
rect 16117 13172 16129 13175
rect 13004 13144 16129 13172
rect 16117 13141 16129 13144
rect 16163 13141 16175 13175
rect 16592 13172 16620 13212
rect 16666 13200 16672 13252
rect 16724 13200 16730 13252
rect 17236 13240 17264 13339
rect 17402 13336 17408 13388
rect 17460 13336 17466 13388
rect 17954 13376 17960 13388
rect 17512 13348 17960 13376
rect 17512 13240 17540 13348
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 18156 13385 18184 13416
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 18233 13379 18291 13385
rect 18233 13345 18245 13379
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18325 13379 18383 13385
rect 18325 13345 18337 13379
rect 18371 13376 18383 13379
rect 18524 13376 18552 13484
rect 18708 13484 18972 13512
rect 18708 13453 18736 13484
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 20530 13512 20536 13524
rect 19720 13484 20536 13512
rect 18693 13447 18751 13453
rect 18693 13413 18705 13447
rect 18739 13413 18751 13447
rect 19720 13444 19748 13484
rect 20530 13472 20536 13484
rect 20588 13512 20594 13524
rect 21174 13512 21180 13524
rect 20588 13484 21180 13512
rect 20588 13472 20594 13484
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 21634 13472 21640 13524
rect 21692 13472 21698 13524
rect 21818 13472 21824 13524
rect 21876 13472 21882 13524
rect 22186 13472 22192 13524
rect 22244 13472 22250 13524
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 24213 13515 24271 13521
rect 23891 13484 24164 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 20806 13444 20812 13456
rect 18693 13407 18751 13413
rect 18892 13416 19748 13444
rect 18371 13348 18552 13376
rect 18371 13345 18383 13348
rect 18325 13339 18383 13345
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 18156 13308 18184 13339
rect 17696 13280 18184 13308
rect 17236 13212 17540 13240
rect 17696 13172 17724 13280
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 18248 13240 18276 13339
rect 18892 13308 18920 13416
rect 19337 13379 19395 13385
rect 19337 13376 19349 13379
rect 18340 13280 18920 13308
rect 18984 13348 19349 13376
rect 18340 13252 18368 13280
rect 18012 13212 18276 13240
rect 18012 13200 18018 13212
rect 16592 13144 17724 13172
rect 17773 13175 17831 13181
rect 16117 13135 16175 13141
rect 17773 13141 17785 13175
rect 17819 13172 17831 13175
rect 17862 13172 17868 13184
rect 17819 13144 17868 13172
rect 17819 13141 17831 13144
rect 17773 13135 17831 13141
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 18248 13172 18276 13212
rect 18322 13200 18328 13252
rect 18380 13200 18386 13252
rect 18506 13200 18512 13252
rect 18564 13200 18570 13252
rect 18984 13172 19012 13348
rect 19337 13345 19349 13348
rect 19383 13376 19395 13379
rect 19610 13376 19616 13388
rect 19383 13348 19616 13376
rect 19383 13345 19395 13348
rect 19337 13339 19395 13345
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 19720 13385 19748 13416
rect 19904 13416 20812 13444
rect 19904 13385 19932 13416
rect 20806 13404 20812 13416
rect 20864 13444 20870 13456
rect 20864 13416 21404 13444
rect 20864 13404 20870 13416
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 19242 13268 19248 13320
rect 19300 13268 19306 13320
rect 19996 13240 20024 13339
rect 20254 13336 20260 13388
rect 20312 13336 20318 13388
rect 20438 13336 20444 13388
rect 20496 13376 20502 13388
rect 20496 13348 20576 13376
rect 20496 13336 20502 13348
rect 19076 13212 20024 13240
rect 20073 13243 20131 13249
rect 19076 13184 19104 13212
rect 20073 13209 20085 13243
rect 20119 13240 20131 13243
rect 20162 13240 20168 13252
rect 20119 13212 20168 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 20162 13200 20168 13212
rect 20220 13200 20226 13252
rect 18248 13144 19012 13172
rect 19058 13132 19064 13184
rect 19116 13132 19122 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 20272 13172 20300 13336
rect 20548 13317 20576 13348
rect 20714 13336 20720 13388
rect 20772 13336 20778 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21376 13385 21404 13416
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 21232 13348 21281 13376
rect 21232 13336 21238 13348
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 21269 13339 21327 13345
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 21542 13336 21548 13388
rect 21600 13336 21606 13388
rect 21652 13385 21680 13472
rect 22646 13404 22652 13456
rect 22704 13444 22710 13456
rect 24136 13444 24164 13484
rect 24213 13481 24225 13515
rect 24259 13512 24271 13515
rect 24946 13512 24952 13524
rect 24259 13484 24952 13512
rect 24259 13481 24271 13484
rect 24213 13475 24271 13481
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 25038 13472 25044 13524
rect 25096 13512 25102 13524
rect 25774 13512 25780 13524
rect 25096 13484 25780 13512
rect 25096 13472 25102 13484
rect 25774 13472 25780 13484
rect 25832 13472 25838 13524
rect 25866 13472 25872 13524
rect 25924 13472 25930 13524
rect 27065 13515 27123 13521
rect 26068 13484 27016 13512
rect 24302 13444 24308 13456
rect 22704 13416 23612 13444
rect 24136 13416 24308 13444
rect 22704 13404 22710 13416
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13345 21695 13379
rect 21637 13339 21695 13345
rect 22094 13336 22100 13388
rect 22152 13336 22158 13388
rect 22738 13336 22744 13388
rect 22796 13336 22802 13388
rect 22940 13385 22968 13416
rect 23584 13388 23612 13416
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 26068 13444 26096 13484
rect 26789 13447 26847 13453
rect 26789 13444 26801 13447
rect 25608 13416 26096 13444
rect 26160 13416 26801 13444
rect 24029 13389 24087 13395
rect 24029 13388 24041 13389
rect 24075 13388 24087 13389
rect 25608 13388 25636 13416
rect 22925 13379 22983 13385
rect 22925 13345 22937 13379
rect 22971 13345 22983 13379
rect 22925 13339 22983 13345
rect 23109 13345 23167 13351
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13277 20591 13311
rect 20732 13308 20760 13336
rect 21560 13308 21588 13336
rect 23109 13311 23121 13345
rect 23155 13311 23167 13345
rect 23566 13336 23572 13388
rect 23624 13336 23630 13388
rect 23658 13336 23664 13388
rect 23716 13336 23722 13388
rect 24026 13336 24032 13388
rect 24084 13386 24090 13388
rect 24084 13358 24119 13386
rect 24084 13336 24090 13358
rect 24210 13336 24216 13388
rect 24268 13336 24274 13388
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 24765 13379 24823 13385
rect 24765 13376 24777 13379
rect 24728 13348 24777 13376
rect 24728 13336 24734 13348
rect 24765 13345 24777 13348
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 23109 13308 23167 13311
rect 23198 13308 23204 13320
rect 20732 13280 21588 13308
rect 22066 13280 23204 13308
rect 20533 13271 20591 13277
rect 22066 13240 22094 13280
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 24394 13268 24400 13320
rect 24452 13308 24458 13320
rect 25056 13308 25084 13339
rect 25590 13336 25596 13388
rect 25648 13336 25654 13388
rect 26160 13385 26188 13416
rect 26789 13413 26801 13416
rect 26835 13413 26847 13447
rect 26988 13444 27016 13484
rect 27065 13481 27077 13515
rect 27111 13512 27123 13515
rect 27111 13484 28580 13512
rect 27111 13481 27123 13484
rect 27065 13475 27123 13481
rect 26988 13416 27660 13444
rect 26789 13407 26847 13413
rect 26145 13379 26203 13385
rect 26145 13376 26157 13379
rect 25792 13348 26157 13376
rect 24452 13280 25084 13308
rect 24452 13268 24458 13280
rect 21468 13212 22094 13240
rect 21468 13184 21496 13212
rect 23290 13200 23296 13252
rect 23348 13200 23354 13252
rect 25792 13184 25820 13348
rect 26145 13345 26157 13348
rect 26191 13345 26203 13379
rect 26145 13339 26203 13345
rect 26418 13336 26424 13388
rect 26476 13336 26482 13388
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 26326 13268 26332 13320
rect 26384 13308 26390 13320
rect 26528 13308 26556 13339
rect 26694 13336 26700 13388
rect 26752 13336 26758 13388
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 26927 13348 27016 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 26988 13320 27016 13348
rect 27430 13336 27436 13388
rect 27488 13376 27494 13388
rect 27525 13379 27583 13385
rect 27525 13376 27537 13379
rect 27488 13348 27537 13376
rect 27488 13336 27494 13348
rect 27525 13345 27537 13348
rect 27571 13345 27583 13379
rect 27632 13376 27660 13416
rect 27706 13404 27712 13456
rect 27764 13444 27770 13456
rect 28074 13444 28080 13456
rect 27764 13416 28080 13444
rect 27764 13404 27770 13416
rect 28074 13404 28080 13416
rect 28132 13404 28138 13456
rect 28350 13404 28356 13456
rect 28408 13404 28414 13456
rect 27893 13379 27951 13385
rect 27893 13376 27905 13379
rect 27632 13348 27905 13376
rect 27525 13339 27583 13345
rect 27893 13345 27905 13348
rect 27939 13345 27951 13379
rect 27893 13339 27951 13345
rect 27985 13379 28043 13385
rect 27985 13345 27997 13379
rect 28031 13376 28043 13379
rect 28368 13376 28396 13404
rect 28552 13385 28580 13484
rect 30466 13472 30472 13524
rect 30524 13472 30530 13524
rect 30834 13472 30840 13524
rect 30892 13472 30898 13524
rect 31018 13472 31024 13524
rect 31076 13472 31082 13524
rect 30484 13444 30512 13472
rect 30852 13444 30880 13472
rect 30484 13416 30696 13444
rect 28031 13348 28396 13376
rect 28537 13379 28595 13385
rect 28031 13345 28043 13348
rect 27985 13339 28043 13345
rect 28537 13345 28549 13379
rect 28583 13345 28595 13379
rect 28537 13339 28595 13345
rect 28997 13379 29055 13385
rect 28997 13345 29009 13379
rect 29043 13345 29055 13379
rect 28997 13339 29055 13345
rect 26384 13280 26556 13308
rect 26384 13268 26390 13280
rect 26970 13268 26976 13320
rect 27028 13268 27034 13320
rect 27062 13268 27068 13320
rect 27120 13308 27126 13320
rect 27706 13308 27712 13320
rect 27120 13280 27712 13308
rect 27120 13268 27126 13280
rect 27706 13268 27712 13280
rect 27764 13268 27770 13320
rect 27801 13311 27859 13317
rect 27801 13277 27813 13311
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 27246 13200 27252 13252
rect 27304 13240 27310 13252
rect 27816 13240 27844 13271
rect 27304 13212 27844 13240
rect 27304 13200 27310 13212
rect 19484 13144 20300 13172
rect 19484 13132 19490 13144
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 20990 13172 20996 13184
rect 20404 13144 20996 13172
rect 20404 13132 20410 13144
rect 20990 13132 20996 13144
rect 21048 13172 21054 13184
rect 21450 13172 21456 13184
rect 21048 13144 21456 13172
rect 21048 13132 21054 13144
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 21910 13172 21916 13184
rect 21600 13144 21916 13172
rect 21600 13132 21606 13144
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 24302 13132 24308 13184
rect 24360 13172 24366 13184
rect 24949 13175 25007 13181
rect 24949 13172 24961 13175
rect 24360 13144 24961 13172
rect 24360 13132 24366 13144
rect 24949 13141 24961 13144
rect 24995 13141 25007 13175
rect 24949 13135 25007 13141
rect 25774 13132 25780 13184
rect 25832 13132 25838 13184
rect 27908 13172 27936 13339
rect 28169 13311 28227 13317
rect 28169 13277 28181 13311
rect 28215 13308 28227 13311
rect 29012 13308 29040 13339
rect 29086 13336 29092 13388
rect 29144 13376 29150 13388
rect 29457 13379 29515 13385
rect 29457 13376 29469 13379
rect 29144 13348 29469 13376
rect 29144 13336 29150 13348
rect 29457 13345 29469 13348
rect 29503 13345 29515 13379
rect 29457 13339 29515 13345
rect 29733 13379 29791 13385
rect 29733 13345 29745 13379
rect 29779 13376 29791 13379
rect 29822 13376 29828 13388
rect 29779 13348 29828 13376
rect 29779 13345 29791 13348
rect 29733 13339 29791 13345
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 30668 13385 30696 13416
rect 30760 13416 30880 13444
rect 30760 13385 30788 13416
rect 31036 13385 31064 13472
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30469 13379 30527 13385
rect 30469 13376 30481 13379
rect 30055 13348 30481 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30469 13345 30481 13348
rect 30515 13345 30527 13379
rect 30469 13339 30527 13345
rect 30653 13379 30711 13385
rect 30653 13345 30665 13379
rect 30699 13345 30711 13379
rect 30653 13339 30711 13345
rect 30745 13379 30803 13385
rect 30745 13345 30757 13379
rect 30791 13345 30803 13379
rect 30929 13379 30987 13385
rect 30929 13376 30941 13379
rect 30745 13339 30803 13345
rect 30852 13348 30941 13376
rect 28215 13280 29040 13308
rect 28215 13277 28227 13280
rect 28169 13271 28227 13277
rect 28626 13200 28632 13252
rect 28684 13200 28690 13252
rect 29454 13172 29460 13184
rect 27908 13144 29460 13172
rect 29454 13132 29460 13144
rect 29512 13172 29518 13184
rect 30852 13172 30880 13348
rect 30929 13345 30941 13348
rect 30975 13345 30987 13379
rect 30929 13339 30987 13345
rect 31021 13379 31079 13385
rect 31021 13345 31033 13379
rect 31067 13345 31079 13379
rect 31021 13339 31079 13345
rect 29512 13144 30880 13172
rect 29512 13132 29518 13144
rect 552 13082 31648 13104
rect 552 13030 4285 13082
rect 4337 13030 4349 13082
rect 4401 13030 4413 13082
rect 4465 13030 4477 13082
rect 4529 13030 4541 13082
rect 4593 13030 12059 13082
rect 12111 13030 12123 13082
rect 12175 13030 12187 13082
rect 12239 13030 12251 13082
rect 12303 13030 12315 13082
rect 12367 13030 19833 13082
rect 19885 13030 19897 13082
rect 19949 13030 19961 13082
rect 20013 13030 20025 13082
rect 20077 13030 20089 13082
rect 20141 13030 27607 13082
rect 27659 13030 27671 13082
rect 27723 13030 27735 13082
rect 27787 13030 27799 13082
rect 27851 13030 27863 13082
rect 27915 13030 31648 13082
rect 552 13008 31648 13030
rect 3697 12971 3755 12977
rect 3697 12937 3709 12971
rect 3743 12968 3755 12971
rect 4154 12968 4160 12980
rect 3743 12940 4160 12968
rect 3743 12937 3755 12940
rect 3697 12931 3755 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6328 12940 7205 12968
rect 6328 12928 6334 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7926 12968 7932 12980
rect 7708 12940 7932 12968
rect 7708 12928 7714 12940
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9490 12968 9496 12980
rect 9272 12940 9496 12968
rect 9272 12928 9278 12940
rect 9490 12928 9496 12940
rect 9548 12968 9554 12980
rect 9548 12940 10456 12968
rect 9548 12928 9554 12940
rect 10428 12912 10456 12940
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11422 12968 11428 12980
rect 11020 12940 11428 12968
rect 11020 12928 11026 12940
rect 11422 12928 11428 12940
rect 11480 12968 11486 12980
rect 11480 12940 12664 12968
rect 11480 12928 11486 12940
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 5442 12900 5448 12912
rect 2832 12872 5448 12900
rect 2832 12860 2838 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 9582 12900 9588 12912
rect 6932 12872 8340 12900
rect 6932 12844 6960 12872
rect 934 12792 940 12844
rect 992 12832 998 12844
rect 1029 12835 1087 12841
rect 1029 12832 1041 12835
rect 992 12804 1041 12832
rect 992 12792 998 12804
rect 1029 12801 1041 12804
rect 1075 12801 1087 12835
rect 1029 12795 1087 12801
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3200 12804 4384 12832
rect 3200 12792 3206 12804
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2372 12736 2438 12764
rect 2372 12724 2378 12736
rect 3418 12724 3424 12776
rect 3476 12724 3482 12776
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 3602 12764 3608 12776
rect 3559 12736 3608 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12733 3847 12767
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3789 12727 3847 12733
rect 3896 12736 4077 12764
rect 1302 12656 1308 12708
rect 1360 12656 1366 12708
rect 3436 12696 3464 12724
rect 3804 12696 3832 12727
rect 3896 12708 3924 12736
rect 4065 12733 4077 12736
rect 4111 12733 4123 12767
rect 4065 12727 4123 12733
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12764 4215 12767
rect 4246 12764 4252 12776
rect 4203 12736 4252 12764
rect 4203 12733 4215 12736
rect 4157 12727 4215 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4356 12764 4384 12804
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7650 12792 7656 12844
rect 7708 12792 7714 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7800 12804 7849 12832
rect 7800 12792 7806 12804
rect 7837 12801 7849 12804
rect 7883 12832 7895 12835
rect 8110 12832 8116 12844
rect 7883 12804 8116 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8312 12832 8340 12872
rect 9324 12872 9588 12900
rect 9033 12835 9091 12841
rect 8312 12804 8524 12832
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4356 12736 4721 12764
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5626 12764 5632 12776
rect 4847 12736 5632 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 3436 12668 3832 12696
rect 3878 12656 3884 12708
rect 3936 12656 3942 12708
rect 3970 12656 3976 12708
rect 4028 12656 4034 12708
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 4816 12696 4844 12727
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 8496 12764 8524 12804
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9122 12832 9128 12844
rect 9079 12804 9128 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 8846 12764 8852 12776
rect 5736 12736 8432 12764
rect 8496 12736 8852 12764
rect 4580 12668 4844 12696
rect 4580 12656 4586 12668
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 4948 12668 5396 12696
rect 4948 12656 4954 12668
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4341 12631 4399 12637
rect 4341 12628 4353 12631
rect 4212 12600 4353 12628
rect 4212 12588 4218 12600
rect 4341 12597 4353 12600
rect 4387 12597 4399 12631
rect 4341 12591 4399 12597
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 5368 12628 5396 12668
rect 5442 12656 5448 12708
rect 5500 12696 5506 12708
rect 5736 12696 5764 12736
rect 7009 12699 7067 12705
rect 7009 12696 7021 12699
rect 5500 12668 5764 12696
rect 5920 12668 7021 12696
rect 5500 12656 5506 12668
rect 5920 12628 5948 12668
rect 7009 12665 7021 12668
rect 7055 12696 7067 12699
rect 7098 12696 7104 12708
rect 7055 12668 7104 12696
rect 7055 12665 7067 12668
rect 7009 12659 7067 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 8294 12696 8300 12708
rect 7852 12668 8300 12696
rect 5368 12600 5948 12628
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6733 12631 6791 12637
rect 6733 12628 6745 12631
rect 6604 12600 6745 12628
rect 6604 12588 6610 12600
rect 6733 12597 6745 12600
rect 6779 12597 6791 12631
rect 6733 12591 6791 12597
rect 7561 12631 7619 12637
rect 7561 12597 7573 12631
rect 7607 12628 7619 12631
rect 7852 12628 7880 12668
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 8404 12696 8432 12736
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 9324 12773 9352 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 9953 12903 10011 12909
rect 9953 12869 9965 12903
rect 9999 12900 10011 12903
rect 9999 12872 10277 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9600 12804 10057 12832
rect 9490 12773 9496 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9457 12767 9496 12773
rect 9457 12733 9469 12767
rect 9457 12727 9496 12733
rect 9490 12724 9496 12727
rect 9548 12724 9554 12776
rect 9600 12773 9628 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10249 12832 10277 12872
rect 10410 12860 10416 12912
rect 10468 12900 10474 12912
rect 10778 12900 10784 12912
rect 10468 12872 10784 12900
rect 10468 12860 10474 12872
rect 10778 12860 10784 12872
rect 10836 12900 10842 12912
rect 10836 12872 10916 12900
rect 10836 12860 10842 12872
rect 10888 12841 10916 12872
rect 10873 12835 10931 12841
rect 10249 12804 10548 12832
rect 10045 12795 10103 12801
rect 10520 12773 10548 12804
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11146 12832 11152 12844
rect 10919 12804 11152 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11974 12832 11980 12844
rect 11379 12804 11980 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12636 12832 12664 12940
rect 15102 12928 15108 12980
rect 15160 12928 15166 12980
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 16390 12968 16396 12980
rect 15252 12940 16396 12968
rect 15252 12928 15258 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17497 12971 17555 12977
rect 17497 12968 17509 12971
rect 16816 12940 17509 12968
rect 16816 12928 16822 12940
rect 17497 12937 17509 12940
rect 17543 12968 17555 12971
rect 17543 12940 17632 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 13078 12860 13084 12912
rect 13136 12900 13142 12912
rect 13136 12872 14504 12900
rect 13136 12860 13142 12872
rect 14476 12841 14504 12872
rect 14461 12835 14519 12841
rect 12636 12804 14228 12832
rect 14200 12776 14228 12804
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12832 14979 12835
rect 15120 12832 15148 12928
rect 15657 12903 15715 12909
rect 15657 12869 15669 12903
rect 15703 12900 15715 12903
rect 15746 12900 15752 12912
rect 15703 12872 15752 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 14967 12804 15148 12832
rect 17604 12832 17632 12940
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 18322 12968 18328 12980
rect 17828 12940 18328 12968
rect 17828 12928 17834 12940
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 18414 12928 18420 12980
rect 18472 12928 18478 12980
rect 19242 12968 19248 12980
rect 18892 12940 19248 12968
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 17604 12804 18153 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18892 12832 18920 12940
rect 19242 12928 19248 12940
rect 19300 12968 19306 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 19300 12940 19625 12968
rect 19300 12928 19306 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 20220 12940 20453 12968
rect 20220 12928 20226 12940
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20441 12931 20499 12937
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 19337 12903 19395 12909
rect 19337 12900 19349 12903
rect 19208 12872 19349 12900
rect 19208 12860 19214 12872
rect 19337 12869 19349 12872
rect 19383 12869 19395 12903
rect 19337 12863 19395 12869
rect 19518 12860 19524 12912
rect 19576 12900 19582 12912
rect 20070 12900 20076 12912
rect 19576 12872 20076 12900
rect 19576 12860 19582 12872
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 18141 12795 18199 12801
rect 18248 12804 18920 12832
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12733 9643 12767
rect 9585 12727 9643 12733
rect 9815 12767 9873 12773
rect 9815 12733 9827 12767
rect 9861 12764 9873 12767
rect 10505 12767 10563 12773
rect 9861 12736 10088 12764
rect 9861 12733 9873 12736
rect 9815 12727 9873 12733
rect 10060 12708 10088 12736
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 10652 12736 10701 12764
rect 10652 12724 10658 12736
rect 10689 12733 10701 12736
rect 10735 12733 10747 12767
rect 10689 12727 10747 12733
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 8404 12668 9689 12696
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 10318 12696 10324 12708
rect 10275 12668 10324 12696
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 10413 12699 10471 12705
rect 10413 12665 10425 12699
rect 10459 12665 10471 12699
rect 10704 12696 10732 12727
rect 10778 12724 10784 12776
rect 10836 12724 10842 12776
rect 11057 12767 11115 12773
rect 11057 12733 11069 12767
rect 11103 12764 11115 12767
rect 11103 12736 11192 12764
rect 11103 12733 11115 12736
rect 11057 12727 11115 12733
rect 10704 12668 11100 12696
rect 10413 12659 10471 12665
rect 7607 12600 7880 12628
rect 7607 12597 7619 12600
rect 7561 12591 7619 12597
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 7984 12600 8401 12628
rect 7984 12588 7990 12600
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 8389 12591 8447 12597
rect 8754 12588 8760 12640
rect 8812 12588 8818 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9306 12628 9312 12640
rect 9088 12600 9312 12628
rect 9088 12588 9094 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10428 12628 10456 12659
rect 11072 12640 11100 12668
rect 10008 12600 10456 12628
rect 10008 12588 10014 12600
rect 11054 12588 11060 12640
rect 11112 12588 11118 12640
rect 11164 12628 11192 12736
rect 13998 12724 14004 12776
rect 14056 12724 14062 12776
rect 14182 12724 14188 12776
rect 14240 12724 14246 12776
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 11609 12699 11667 12705
rect 11609 12696 11621 12699
rect 11287 12668 11621 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 11609 12665 11621 12668
rect 11655 12665 11667 12699
rect 11609 12659 11667 12665
rect 11698 12656 11704 12708
rect 11756 12656 11762 12708
rect 12342 12656 12348 12708
rect 12400 12656 12406 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 14292 12696 14320 12727
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15252 12736 15761 12764
rect 15252 12724 15258 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 15749 12727 15807 12733
rect 18046 12724 18052 12776
rect 18104 12764 18110 12776
rect 18248 12764 18276 12804
rect 18892 12773 18920 12804
rect 18104 12736 18276 12764
rect 18325 12767 18383 12773
rect 18104 12724 18110 12736
rect 18325 12733 18337 12767
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12733 19027 12767
rect 18969 12727 19027 12733
rect 19095 12767 19153 12773
rect 19095 12733 19107 12767
rect 19141 12764 19153 12767
rect 20180 12764 20208 12928
rect 20456 12900 20484 12931
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 20588 12940 20761 12968
rect 20588 12928 20594 12940
rect 20456 12872 20668 12900
rect 20346 12792 20352 12844
rect 20404 12792 20410 12844
rect 20640 12776 20668 12872
rect 20733 12832 20761 12940
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 20864 12940 21097 12968
rect 20864 12928 20870 12940
rect 21085 12937 21097 12940
rect 21131 12968 21143 12971
rect 21266 12968 21272 12980
rect 21131 12940 21272 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 21453 12971 21511 12977
rect 21453 12937 21465 12971
rect 21499 12968 21511 12971
rect 22094 12968 22100 12980
rect 21499 12940 22100 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 23293 12971 23351 12977
rect 23293 12968 23305 12971
rect 22796 12940 23305 12968
rect 22796 12928 22802 12940
rect 23293 12937 23305 12940
rect 23339 12937 23351 12971
rect 23293 12931 23351 12937
rect 23477 12971 23535 12977
rect 23477 12937 23489 12971
rect 23523 12968 23535 12971
rect 23658 12968 23664 12980
rect 23523 12940 23664 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 23658 12928 23664 12940
rect 23716 12928 23722 12980
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24578 12968 24584 12980
rect 24535 12940 24584 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 24949 12971 25007 12977
rect 24949 12968 24961 12971
rect 24912 12940 24961 12968
rect 24912 12928 24918 12940
rect 24949 12937 24961 12940
rect 24995 12968 25007 12971
rect 25038 12968 25044 12980
rect 24995 12940 25044 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 25133 12971 25191 12977
rect 25133 12937 25145 12971
rect 25179 12968 25191 12971
rect 25590 12968 25596 12980
rect 25179 12940 25596 12968
rect 25179 12937 25191 12940
rect 25133 12931 25191 12937
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 25774 12928 25780 12980
rect 25832 12928 25838 12980
rect 25866 12928 25872 12980
rect 25924 12968 25930 12980
rect 25924 12940 27282 12968
rect 25924 12928 25930 12940
rect 20898 12860 20904 12912
rect 20956 12900 20962 12912
rect 20993 12903 21051 12909
rect 20993 12900 21005 12903
rect 20956 12872 21005 12900
rect 20956 12860 20962 12872
rect 20993 12869 21005 12872
rect 21039 12869 21051 12903
rect 20993 12863 21051 12869
rect 21729 12903 21787 12909
rect 21729 12869 21741 12903
rect 21775 12900 21787 12903
rect 21775 12872 27200 12900
rect 21775 12869 21787 12872
rect 21729 12863 21787 12869
rect 20733 12804 21772 12832
rect 19141 12736 20208 12764
rect 20441 12767 20499 12773
rect 19141 12733 19153 12736
rect 19095 12727 19153 12733
rect 20441 12733 20453 12767
rect 20487 12764 20499 12767
rect 20533 12767 20591 12773
rect 20533 12764 20545 12767
rect 20487 12736 20545 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20533 12733 20545 12736
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 14458 12696 14464 12708
rect 13872 12668 14464 12696
rect 13872 12656 13878 12668
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 14918 12656 14924 12708
rect 14976 12696 14982 12708
rect 15105 12699 15163 12705
rect 15105 12696 15117 12699
rect 14976 12668 15117 12696
rect 14976 12656 14982 12668
rect 15105 12665 15117 12668
rect 15151 12665 15163 12699
rect 15105 12659 15163 12665
rect 15470 12656 15476 12708
rect 15528 12656 15534 12708
rect 16025 12699 16083 12705
rect 16025 12665 16037 12699
rect 16071 12665 16083 12699
rect 17310 12696 17316 12708
rect 17250 12668 17316 12696
rect 16025 12659 16083 12665
rect 11716 12628 11744 12656
rect 11164 12600 11744 12628
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 15194 12628 15200 12640
rect 14332 12600 15200 12628
rect 14332 12588 14338 12600
rect 15194 12588 15200 12600
rect 15252 12628 15258 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15252 12600 15301 12628
rect 15252 12588 15258 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 15289 12591 15347 12597
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 15838 12628 15844 12640
rect 15427 12600 15844 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 16040 12628 16068 12659
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17862 12656 17868 12708
rect 17920 12696 17926 12708
rect 18340 12696 18368 12727
rect 17920 12668 18368 12696
rect 17920 12656 17926 12668
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 18524 12696 18552 12727
rect 18472 12668 18552 12696
rect 18472 12656 18478 12668
rect 16758 12628 16764 12640
rect 16040 12600 16764 12628
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 17586 12588 17592 12640
rect 17644 12588 17650 12640
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18708 12628 18736 12727
rect 18984 12696 19012 12727
rect 18984 12668 19104 12696
rect 19076 12640 19104 12668
rect 19426 12656 19432 12708
rect 19484 12656 19490 12708
rect 20456 12696 20484 12727
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20680 12736 20729 12764
rect 20680 12724 20686 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20806 12724 20812 12776
rect 20864 12724 20870 12776
rect 21100 12773 21128 12804
rect 21085 12767 21143 12773
rect 21085 12733 21097 12767
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 19536 12668 20484 12696
rect 18012 12600 18736 12628
rect 18012 12588 18018 12600
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19536 12628 19564 12668
rect 20898 12656 20904 12708
rect 20956 12696 20962 12708
rect 21192 12696 21220 12727
rect 21266 12724 21272 12776
rect 21324 12764 21330 12776
rect 21744 12773 21772 12804
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 22922 12832 22928 12844
rect 22060 12804 22928 12832
rect 22060 12792 22066 12804
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 24118 12832 24124 12844
rect 23032 12804 24124 12832
rect 21545 12767 21603 12773
rect 21545 12764 21557 12767
rect 21324 12736 21557 12764
rect 21324 12724 21330 12736
rect 21545 12733 21557 12736
rect 21591 12733 21603 12767
rect 21545 12727 21603 12733
rect 21729 12767 21787 12773
rect 21729 12733 21741 12767
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 23032 12764 23060 12804
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24213 12835 24271 12841
rect 24213 12801 24225 12835
rect 24259 12832 24271 12835
rect 25130 12832 25136 12844
rect 24259 12804 25136 12832
rect 24259 12801 24271 12804
rect 24213 12795 24271 12801
rect 25130 12792 25136 12804
rect 25188 12832 25194 12844
rect 25188 12804 25636 12832
rect 25188 12792 25194 12804
rect 24673 12767 24731 12773
rect 22520 12736 23060 12764
rect 23124 12736 24532 12764
rect 22520 12724 22526 12736
rect 23124 12705 23152 12736
rect 22649 12699 22707 12705
rect 22649 12696 22661 12699
rect 20956 12668 22661 12696
rect 20956 12656 20962 12668
rect 22649 12665 22661 12668
rect 22695 12696 22707 12699
rect 23109 12699 23167 12705
rect 23109 12696 23121 12699
rect 22695 12668 23121 12696
rect 22695 12665 22707 12668
rect 22649 12659 22707 12665
rect 23109 12665 23121 12668
rect 23155 12665 23167 12699
rect 23109 12659 23167 12665
rect 23198 12656 23204 12708
rect 23256 12696 23262 12708
rect 23937 12699 23995 12705
rect 23937 12696 23949 12699
rect 23256 12668 23949 12696
rect 23256 12656 23262 12668
rect 23937 12665 23949 12668
rect 23983 12665 23995 12699
rect 23937 12659 23995 12665
rect 19116 12600 19564 12628
rect 19116 12588 19122 12600
rect 19610 12588 19616 12640
rect 19668 12588 19674 12640
rect 19797 12631 19855 12637
rect 19797 12597 19809 12631
rect 19843 12628 19855 12631
rect 21542 12628 21548 12640
rect 19843 12600 21548 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21692 12600 22109 12628
rect 21692 12588 21698 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22097 12591 22155 12597
rect 23319 12631 23377 12637
rect 23319 12597 23331 12631
rect 23365 12628 23377 12631
rect 23566 12628 23572 12640
rect 23365 12600 23572 12628
rect 23365 12597 23377 12600
rect 23319 12591 23377 12597
rect 23566 12588 23572 12600
rect 23624 12628 23630 12640
rect 24394 12628 24400 12640
rect 23624 12600 24400 12628
rect 23624 12588 23630 12600
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 24504 12628 24532 12736
rect 24673 12733 24685 12767
rect 24719 12764 24731 12767
rect 24854 12764 24860 12776
rect 24719 12736 24860 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 24964 12736 25329 12764
rect 24762 12656 24768 12708
rect 24820 12656 24826 12708
rect 24670 12628 24676 12640
rect 24504 12600 24676 12628
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 24964 12637 24992 12736
rect 25317 12733 25329 12736
rect 25363 12764 25375 12767
rect 25406 12764 25412 12776
rect 25363 12736 25412 12764
rect 25363 12733 25375 12736
rect 25317 12727 25375 12733
rect 25406 12724 25412 12736
rect 25464 12724 25470 12776
rect 25608 12773 25636 12804
rect 25593 12767 25651 12773
rect 25593 12733 25605 12767
rect 25639 12733 25651 12767
rect 25593 12727 25651 12733
rect 26697 12767 26755 12773
rect 26697 12733 26709 12767
rect 26743 12764 26755 12767
rect 27062 12764 27068 12776
rect 26743 12736 27068 12764
rect 26743 12733 26755 12736
rect 26697 12727 26755 12733
rect 27062 12724 27068 12736
rect 27120 12724 27126 12776
rect 27172 12764 27200 12872
rect 27254 12832 27282 12940
rect 27338 12928 27344 12980
rect 27396 12968 27402 12980
rect 27433 12971 27491 12977
rect 27433 12968 27445 12971
rect 27396 12940 27445 12968
rect 27396 12928 27402 12940
rect 27433 12937 27445 12940
rect 27479 12937 27491 12971
rect 27433 12931 27491 12937
rect 27709 12971 27767 12977
rect 27709 12937 27721 12971
rect 27755 12968 27767 12971
rect 27982 12968 27988 12980
rect 27755 12940 27988 12968
rect 27755 12937 27767 12940
rect 27709 12931 27767 12937
rect 27982 12928 27988 12940
rect 28040 12928 28046 12980
rect 29822 12928 29828 12980
rect 29880 12968 29886 12980
rect 29917 12971 29975 12977
rect 29917 12968 29929 12971
rect 29880 12940 29929 12968
rect 29880 12928 29886 12940
rect 29917 12937 29929 12940
rect 29963 12937 29975 12971
rect 29917 12931 29975 12937
rect 30282 12928 30288 12980
rect 30340 12928 30346 12980
rect 30650 12928 30656 12980
rect 30708 12928 30714 12980
rect 28166 12900 28172 12912
rect 27540 12872 28172 12900
rect 27540 12844 27568 12872
rect 28166 12860 28172 12872
rect 28224 12860 28230 12912
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 27254 12804 27353 12832
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27522 12792 27528 12844
rect 27580 12792 27586 12844
rect 30668 12832 30696 12928
rect 27632 12804 30696 12832
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 27172 12736 27261 12764
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 25038 12656 25044 12708
rect 25096 12696 25102 12708
rect 25096 12668 25452 12696
rect 25096 12656 25102 12668
rect 25424 12637 25452 12668
rect 26326 12656 26332 12708
rect 26384 12656 26390 12708
rect 26878 12656 26884 12708
rect 26936 12656 26942 12708
rect 27264 12696 27292 12727
rect 27430 12724 27436 12776
rect 27488 12764 27494 12776
rect 27632 12764 27660 12804
rect 27488 12736 27660 12764
rect 27985 12767 28043 12773
rect 27488 12724 27494 12736
rect 27985 12733 27997 12767
rect 28031 12764 28043 12767
rect 28258 12764 28264 12776
rect 28031 12736 28264 12764
rect 28031 12733 28043 12736
rect 27985 12727 28043 12733
rect 28258 12724 28264 12736
rect 28316 12724 28322 12776
rect 29932 12773 29960 12804
rect 29917 12767 29975 12773
rect 29917 12733 29929 12767
rect 29963 12733 29975 12767
rect 29917 12727 29975 12733
rect 30009 12767 30067 12773
rect 30009 12733 30021 12767
rect 30055 12733 30067 12767
rect 30009 12727 30067 12733
rect 27709 12699 27767 12705
rect 27709 12696 27721 12699
rect 27264 12668 27721 12696
rect 27709 12665 27721 12668
rect 27755 12665 27767 12699
rect 30024 12696 30052 12727
rect 30374 12724 30380 12776
rect 30432 12724 30438 12776
rect 27709 12659 27767 12665
rect 27816 12668 30052 12696
rect 24949 12631 25007 12637
rect 24949 12597 24961 12631
rect 24995 12597 25007 12631
rect 24949 12591 25007 12597
rect 25409 12631 25467 12637
rect 25409 12597 25421 12631
rect 25455 12597 25467 12631
rect 25409 12591 25467 12597
rect 26970 12588 26976 12640
rect 27028 12628 27034 12640
rect 27816 12628 27844 12668
rect 27028 12600 27844 12628
rect 27893 12631 27951 12637
rect 27028 12588 27034 12600
rect 27893 12597 27905 12631
rect 27939 12628 27951 12631
rect 30392 12628 30420 12724
rect 27939 12600 30420 12628
rect 27939 12597 27951 12600
rect 27893 12591 27951 12597
rect 552 12538 31808 12560
rect 552 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 15946 12538
rect 15998 12486 16010 12538
rect 16062 12486 16074 12538
rect 16126 12486 16138 12538
rect 16190 12486 16202 12538
rect 16254 12486 23720 12538
rect 23772 12486 23784 12538
rect 23836 12486 23848 12538
rect 23900 12486 23912 12538
rect 23964 12486 23976 12538
rect 24028 12486 31494 12538
rect 31546 12486 31558 12538
rect 31610 12486 31622 12538
rect 31674 12486 31686 12538
rect 31738 12486 31750 12538
rect 31802 12486 31808 12538
rect 552 12464 31808 12486
rect 1302 12384 1308 12436
rect 1360 12424 1366 12436
rect 1489 12427 1547 12433
rect 1489 12424 1501 12427
rect 1360 12396 1501 12424
rect 1360 12384 1366 12396
rect 1489 12393 1501 12396
rect 1535 12393 1547 12427
rect 2774 12424 2780 12436
rect 1489 12387 1547 12393
rect 2746 12384 2780 12424
rect 2832 12384 2838 12436
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 3936 12396 4813 12424
rect 3936 12384 3942 12396
rect 4801 12393 4813 12396
rect 4847 12424 4859 12427
rect 5350 12424 5356 12436
rect 4847 12396 5356 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6641 12427 6699 12433
rect 6641 12424 6653 12427
rect 6328 12396 6653 12424
rect 6328 12384 6334 12396
rect 6641 12393 6653 12396
rect 6687 12393 6699 12427
rect 6641 12387 6699 12393
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 8812 12396 9229 12424
rect 8812 12384 8818 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9674 12424 9680 12436
rect 9456 12396 9680 12424
rect 9456 12384 9462 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9877 12396 10180 12424
rect 2409 12359 2467 12365
rect 2409 12325 2421 12359
rect 2455 12356 2467 12359
rect 2746 12356 2774 12384
rect 2455 12328 2774 12356
rect 2455 12325 2467 12328
rect 2409 12319 2467 12325
rect 3970 12316 3976 12368
rect 4028 12316 4034 12368
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4522 12356 4528 12368
rect 4120 12328 4528 12356
rect 4120 12316 4126 12328
rect 4522 12316 4528 12328
rect 4580 12316 4586 12368
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 6362 12356 6368 12368
rect 4672 12328 6368 12356
rect 4672 12316 4678 12328
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 8478 12316 8484 12368
rect 8536 12316 8542 12368
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 9180 12328 9536 12356
rect 9180 12316 9186 12328
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 1719 12260 2084 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 2056 12161 2084 12260
rect 3786 12248 3792 12300
rect 3844 12248 3850 12300
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4246 12288 4252 12300
rect 4203 12260 4252 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 4246 12248 4252 12260
rect 4304 12288 4310 12300
rect 5074 12288 5080 12300
rect 4304 12260 5080 12288
rect 4304 12248 4310 12260
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6549 12291 6607 12297
rect 6135 12260 6224 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 2498 12180 2504 12232
rect 2556 12180 2562 12232
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 4614 12180 4620 12232
rect 4672 12180 4678 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 2041 12155 2099 12161
rect 2041 12121 2053 12155
rect 2087 12121 2099 12155
rect 2700 12152 2728 12180
rect 6196 12161 6224 12260
rect 6549 12257 6561 12291
rect 6595 12288 6607 12291
rect 7374 12288 7380 12300
rect 6595 12260 7380 12288
rect 6595 12257 6607 12260
rect 6549 12251 6607 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 6871 12192 6960 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 6181 12155 6239 12161
rect 2700 12124 6132 12152
rect 2041 12115 2099 12121
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 3326 12084 3332 12096
rect 2188 12056 3332 12084
rect 2188 12044 2194 12056
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4614 12084 4620 12096
rect 4387 12056 4620 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5350 12084 5356 12096
rect 5215 12056 5356 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 5994 12084 6000 12096
rect 5951 12056 6000 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6104 12084 6132 12124
rect 6181 12121 6193 12155
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 6932 12084 6960 12192
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 9140 12084 9168 12316
rect 9306 12248 9312 12300
rect 9364 12248 9370 12300
rect 9398 12248 9404 12300
rect 9456 12248 9462 12300
rect 9508 12288 9536 12328
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 9877 12356 9905 12396
rect 9640 12328 9905 12356
rect 9640 12316 9646 12328
rect 9950 12316 9956 12368
rect 10008 12316 10014 12368
rect 9766 12288 9772 12300
rect 9508 12260 9772 12288
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12257 9919 12291
rect 9968 12288 9996 12316
rect 10152 12297 10180 12396
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 10284 12396 10640 12424
rect 10284 12384 10290 12396
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12325 10563 12359
rect 10612 12356 10640 12396
rect 11882 12384 11888 12436
rect 11940 12384 11946 12436
rect 14277 12427 14335 12433
rect 14277 12393 14289 12427
rect 14323 12424 14335 12427
rect 14642 12424 14648 12436
rect 14323 12396 14648 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15528 12396 16160 12424
rect 15528 12384 15534 12396
rect 13446 12356 13452 12368
rect 10612 12328 11192 12356
rect 10505 12319 10563 12325
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9968 12260 10057 12288
rect 9861 12251 9919 12257
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 10230 12291 10288 12297
rect 10230 12257 10242 12291
rect 10276 12257 10288 12291
rect 10230 12251 10288 12257
rect 9324 12220 9352 12248
rect 9876 12220 9904 12251
rect 9324 12192 9904 12220
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 10245 12220 10273 12251
rect 10410 12248 10416 12300
rect 10468 12248 10474 12300
rect 10520 12232 10548 12319
rect 11164 12297 11192 12328
rect 11440 12328 13452 12356
rect 11440 12297 11468 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 15565 12359 15623 12365
rect 15565 12356 15577 12359
rect 15068 12328 15577 12356
rect 15068 12316 15074 12328
rect 15565 12325 15577 12328
rect 15611 12325 15623 12359
rect 15565 12319 15623 12325
rect 15746 12316 15752 12368
rect 15804 12365 15810 12368
rect 16132 12365 16160 12396
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16264 12396 16405 12424
rect 16264 12384 16270 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 15804 12359 15839 12365
rect 15827 12356 15839 12359
rect 16117 12359 16175 12365
rect 15827 12328 16068 12356
rect 15827 12325 15839 12328
rect 15804 12319 15839 12325
rect 15804 12316 15810 12319
rect 10602 12291 10660 12297
rect 10602 12257 10614 12291
rect 10648 12257 10660 12291
rect 10602 12251 10660 12257
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 9999 12192 10273 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 10042 12152 10048 12164
rect 9784 12124 10048 12152
rect 6104 12056 9168 12084
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 9784 12084 9812 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10617 12152 10645 12251
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11348 12220 11376 12251
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11756 12260 13584 12288
rect 11756 12248 11762 12260
rect 11790 12220 11796 12232
rect 11112 12192 11796 12220
rect 11112 12180 11118 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 11940 12192 12173 12220
rect 11940 12180 11946 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 10192 12124 10645 12152
rect 10192 12112 10198 12124
rect 10686 12112 10692 12164
rect 10744 12152 10750 12164
rect 11146 12152 11152 12164
rect 10744 12124 11152 12152
rect 10744 12112 10750 12124
rect 11146 12112 11152 12124
rect 11204 12152 11210 12164
rect 13556 12152 13584 12260
rect 13630 12248 13636 12300
rect 13688 12248 13694 12300
rect 13814 12297 13820 12300
rect 13780 12291 13820 12297
rect 13780 12257 13792 12291
rect 13780 12251 13820 12257
rect 13814 12248 13820 12251
rect 13872 12248 13878 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 14148 12260 14657 12288
rect 14148 12248 14154 12260
rect 14645 12257 14657 12260
rect 14691 12288 14703 12291
rect 15286 12288 15292 12300
rect 14691 12260 15292 12288
rect 14691 12257 14703 12260
rect 14645 12251 14703 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15381 12291 15439 12297
rect 15381 12257 15393 12291
rect 15427 12288 15439 12291
rect 15930 12288 15936 12300
rect 15427 12260 15936 12288
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 16040 12288 16068 12328
rect 16117 12325 16129 12359
rect 16163 12325 16175 12359
rect 16408 12356 16436 12387
rect 16758 12384 16764 12436
rect 16816 12384 16822 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 18138 12424 18144 12436
rect 17000 12396 18144 12424
rect 17000 12384 17006 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18325 12427 18383 12433
rect 18325 12424 18337 12427
rect 18288 12396 18337 12424
rect 18288 12384 18294 12396
rect 18325 12393 18337 12396
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18564 12396 18828 12424
rect 18564 12384 18570 12396
rect 16669 12359 16727 12365
rect 16408 12328 16620 12356
rect 16117 12319 16175 12325
rect 16206 12288 16212 12300
rect 16040 12260 16212 12288
rect 16206 12248 16212 12260
rect 16264 12297 16270 12300
rect 16264 12291 16319 12297
rect 16264 12257 16273 12291
rect 16307 12257 16319 12291
rect 16264 12251 16319 12257
rect 16264 12248 16270 12251
rect 16390 12248 16396 12300
rect 16448 12288 16454 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16448 12260 16497 12288
rect 16448 12248 16454 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16592 12288 16620 12328
rect 16669 12325 16681 12359
rect 16715 12356 16727 12359
rect 17034 12356 17040 12368
rect 16715 12328 17040 12356
rect 16715 12325 16727 12328
rect 16669 12319 16727 12325
rect 17034 12316 17040 12328
rect 17092 12316 17098 12368
rect 18156 12356 18184 12384
rect 18693 12359 18751 12365
rect 18693 12356 18705 12359
rect 17144 12328 17908 12356
rect 18156 12328 18705 12356
rect 16850 12288 16856 12300
rect 16592 12260 16856 12288
rect 16485 12251 16543 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 17144 12297 17172 12328
rect 17880 12300 17908 12328
rect 18693 12325 18705 12328
rect 18739 12325 18751 12359
rect 18800 12356 18828 12396
rect 19058 12384 19064 12436
rect 19116 12384 19122 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19208 12396 20116 12424
rect 19208 12384 19214 12396
rect 18800 12328 19840 12356
rect 18693 12319 18751 12325
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 16960 12220 16988 12251
rect 14056 12192 15194 12220
rect 14056 12180 14062 12192
rect 11204 12124 13124 12152
rect 13556 12124 14688 12152
rect 11204 12112 11210 12124
rect 13096 12096 13124 12124
rect 9723 12056 9812 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10778 12044 10784 12096
rect 10836 12044 10842 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12584 12056 12817 12084
rect 12584 12044 12590 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13538 12044 13544 12096
rect 13596 12044 13602 12096
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14182 12084 14188 12096
rect 13955 12056 14188 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14660 12084 14688 12124
rect 14734 12112 14740 12164
rect 14792 12112 14798 12164
rect 15166 12152 15194 12192
rect 15948 12192 16988 12220
rect 17236 12220 17264 12251
rect 17402 12248 17408 12300
rect 17460 12248 17466 12300
rect 17862 12248 17868 12300
rect 17920 12248 17926 12300
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 18049 12291 18107 12297
rect 18049 12288 18061 12291
rect 18012 12260 18061 12288
rect 18012 12248 18018 12260
rect 18049 12257 18061 12260
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 17678 12220 17684 12232
rect 17236 12192 17684 12220
rect 15948 12161 15976 12192
rect 17678 12180 17684 12192
rect 17736 12220 17742 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17736 12192 17785 12220
rect 17736 12180 17742 12192
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 18064 12220 18092 12251
rect 18230 12248 18236 12300
rect 18288 12248 18294 12300
rect 18414 12248 18420 12300
rect 18472 12248 18478 12300
rect 18432 12220 18460 12248
rect 18598 12220 18604 12232
rect 18064 12192 18604 12220
rect 17773 12183 17831 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 18708 12220 18736 12319
rect 18782 12248 18788 12300
rect 18840 12248 18846 12300
rect 18874 12248 18880 12300
rect 18932 12248 18938 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19076 12260 19625 12288
rect 18966 12220 18972 12232
rect 18708 12192 18972 12220
rect 18966 12180 18972 12192
rect 19024 12220 19030 12232
rect 19076 12220 19104 12260
rect 19613 12257 19625 12260
rect 19659 12257 19671 12291
rect 19613 12251 19671 12257
rect 19024 12192 19104 12220
rect 19024 12180 19030 12192
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19208 12192 19441 12220
rect 19208 12180 19214 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 19812 12220 19840 12328
rect 20088 12297 20116 12396
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20990 12424 20996 12436
rect 20220 12396 20996 12424
rect 20220 12384 20226 12396
rect 20990 12384 20996 12396
rect 21048 12424 21054 12436
rect 21910 12424 21916 12436
rect 21048 12396 21916 12424
rect 21048 12384 21054 12396
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 22097 12427 22155 12433
rect 22097 12393 22109 12427
rect 22143 12424 22155 12427
rect 22278 12424 22284 12436
rect 22143 12396 22284 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 22572 12396 23796 12424
rect 20180 12356 20208 12384
rect 20533 12359 20591 12365
rect 20180 12328 20392 12356
rect 20073 12291 20131 12297
rect 20073 12257 20085 12291
rect 20119 12257 20131 12291
rect 20073 12251 20131 12257
rect 20162 12248 20168 12300
rect 20220 12248 20226 12300
rect 20364 12297 20392 12328
rect 20533 12325 20545 12359
rect 20579 12356 20591 12359
rect 20622 12356 20628 12368
rect 20579 12328 20628 12356
rect 20579 12325 20591 12328
rect 20533 12319 20591 12325
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 22186 12356 22192 12368
rect 21836 12328 22192 12356
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 20456 12260 21036 12288
rect 20456 12220 20484 12260
rect 19812 12192 20484 12220
rect 19705 12183 19763 12189
rect 15933 12155 15991 12161
rect 15166 12124 15884 12152
rect 15746 12084 15752 12096
rect 14660 12056 15752 12084
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 15856 12084 15884 12124
rect 15933 12121 15945 12155
rect 15979 12121 15991 12155
rect 15933 12115 15991 12121
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 16390 12152 16396 12164
rect 16172 12124 16396 12152
rect 16172 12112 16178 12124
rect 16390 12112 16396 12124
rect 16448 12152 16454 12164
rect 16850 12152 16856 12164
rect 16448 12124 16856 12152
rect 16448 12112 16454 12124
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 17512 12124 18000 12152
rect 17512 12084 17540 12124
rect 15856 12056 17540 12084
rect 17586 12044 17592 12096
rect 17644 12044 17650 12096
rect 17972 12084 18000 12124
rect 18046 12112 18052 12164
rect 18104 12152 18110 12164
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 18104 12124 18521 12152
rect 18104 12112 18110 12124
rect 18509 12121 18521 12124
rect 18555 12152 18567 12155
rect 18690 12152 18696 12164
rect 18555 12124 18696 12152
rect 18555 12121 18567 12124
rect 18509 12115 18567 12121
rect 18690 12112 18696 12124
rect 18748 12152 18754 12164
rect 19536 12152 19564 12183
rect 18748 12124 19564 12152
rect 19720 12152 19748 12183
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 20898 12220 20904 12232
rect 20588 12192 20904 12220
rect 20588 12180 20594 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21008 12220 21036 12260
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 21836 12297 21864 12328
rect 22186 12316 22192 12328
rect 22244 12316 22250 12368
rect 21361 12291 21419 12297
rect 21361 12257 21373 12291
rect 21407 12257 21419 12291
rect 21361 12251 21419 12257
rect 21821 12291 21879 12297
rect 21821 12257 21833 12291
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 21376 12220 21404 12251
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12288 22339 12291
rect 22572 12288 22600 12396
rect 23768 12356 23796 12396
rect 24118 12384 24124 12436
rect 24176 12384 24182 12436
rect 24394 12384 24400 12436
rect 24452 12384 24458 12436
rect 25133 12427 25191 12433
rect 25133 12424 25145 12427
rect 24504 12396 25145 12424
rect 24136 12356 24164 12384
rect 24504 12356 24532 12396
rect 25133 12393 25145 12396
rect 25179 12424 25191 12427
rect 25567 12427 25625 12433
rect 25567 12424 25579 12427
rect 25179 12396 25579 12424
rect 25179 12393 25191 12396
rect 25133 12387 25191 12393
rect 25567 12393 25579 12396
rect 25613 12393 25625 12427
rect 25567 12387 25625 12393
rect 27246 12384 27252 12436
rect 27304 12384 27310 12436
rect 25222 12356 25228 12368
rect 23768 12328 23888 12356
rect 24136 12328 24532 12356
rect 24596 12328 25228 12356
rect 22327 12260 22600 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22646 12248 22652 12300
rect 22704 12288 22710 12300
rect 22741 12291 22799 12297
rect 22741 12288 22753 12291
rect 22704 12260 22753 12288
rect 22704 12248 22710 12260
rect 22741 12257 22753 12260
rect 22787 12288 22799 12291
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 22787 12260 23581 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 23569 12257 23581 12260
rect 23615 12257 23627 12291
rect 23750 12288 23756 12300
rect 23569 12251 23627 12257
rect 23676 12260 23756 12288
rect 21008 12192 21404 12220
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 22465 12223 22523 12229
rect 22465 12220 22477 12223
rect 21784 12192 22477 12220
rect 21784 12180 21790 12192
rect 22465 12189 22477 12192
rect 22511 12220 22523 12223
rect 22511 12192 23060 12220
rect 22511 12189 22523 12192
rect 22465 12183 22523 12189
rect 20162 12152 20168 12164
rect 19720 12124 20168 12152
rect 18748 12112 18754 12124
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 20254 12112 20260 12164
rect 20312 12112 20318 12164
rect 20622 12112 20628 12164
rect 20680 12152 20686 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20680 12124 21005 12152
rect 20680 12112 20686 12124
rect 20993 12121 21005 12124
rect 21039 12152 21051 12155
rect 21082 12152 21088 12164
rect 21039 12124 21088 12152
rect 21039 12121 21051 12124
rect 20993 12115 21051 12121
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 22005 12155 22063 12161
rect 22005 12121 22017 12155
rect 22051 12152 22063 12155
rect 22554 12152 22560 12164
rect 22051 12124 22560 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 22554 12112 22560 12124
rect 22612 12112 22618 12164
rect 23032 12152 23060 12192
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 23676 12152 23704 12260
rect 23750 12248 23756 12260
rect 23808 12248 23814 12300
rect 23860 12297 23888 12328
rect 23845 12291 23903 12297
rect 23845 12257 23857 12291
rect 23891 12288 23903 12291
rect 24026 12288 24032 12300
rect 23891 12260 24032 12288
rect 23891 12257 23903 12260
rect 23845 12251 23903 12257
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 24486 12248 24492 12300
rect 24544 12248 24550 12300
rect 24596 12297 24624 12328
rect 25222 12316 25228 12328
rect 25280 12356 25286 12368
rect 25317 12359 25375 12365
rect 25317 12356 25329 12359
rect 25280 12328 25329 12356
rect 25280 12316 25286 12328
rect 25317 12325 25329 12328
rect 25363 12325 25375 12359
rect 25317 12319 25375 12325
rect 25682 12316 25688 12368
rect 25740 12356 25746 12368
rect 25777 12359 25835 12365
rect 25777 12356 25789 12359
rect 25740 12328 25789 12356
rect 25740 12316 25746 12328
rect 25777 12325 25789 12328
rect 25823 12325 25835 12359
rect 25777 12319 25835 12325
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 27264 12288 27292 12384
rect 24903 12260 27292 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 24118 12220 24124 12232
rect 23768 12192 24124 12220
rect 23768 12164 23796 12192
rect 24118 12180 24124 12192
rect 24176 12180 24182 12232
rect 24210 12180 24216 12232
rect 24268 12180 24274 12232
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 26418 12220 26424 12232
rect 24811 12192 26424 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 27525 12223 27583 12229
rect 27525 12220 27537 12223
rect 26936 12192 27537 12220
rect 26936 12180 26942 12192
rect 27525 12189 27537 12192
rect 27571 12189 27583 12223
rect 27525 12183 27583 12189
rect 22756 12124 22968 12152
rect 23032 12124 23704 12152
rect 19794 12084 19800 12096
rect 17972 12056 19800 12084
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 21726 12084 21732 12096
rect 19935 12056 21732 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 22094 12084 22100 12096
rect 21867 12056 22100 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22278 12044 22284 12096
rect 22336 12084 22342 12096
rect 22756 12084 22784 12124
rect 22336 12056 22784 12084
rect 22336 12044 22342 12056
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 22940 12084 22968 12124
rect 23750 12112 23756 12164
rect 23808 12112 23814 12164
rect 24029 12155 24087 12161
rect 24029 12121 24041 12155
rect 24075 12152 24087 12155
rect 24228 12152 24256 12180
rect 24075 12124 24256 12152
rect 24075 12121 24087 12124
rect 24029 12115 24087 12121
rect 23566 12084 23572 12096
rect 22940 12056 23572 12084
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 24228 12084 24256 12124
rect 25038 12112 25044 12164
rect 25096 12152 25102 12164
rect 25409 12155 25467 12161
rect 25409 12152 25421 12155
rect 25096 12124 25421 12152
rect 25096 12112 25102 12124
rect 25409 12121 25421 12124
rect 25455 12121 25467 12155
rect 25409 12115 25467 12121
rect 25133 12087 25191 12093
rect 25133 12084 25145 12087
rect 24228 12056 25145 12084
rect 25133 12053 25145 12056
rect 25179 12084 25191 12087
rect 25593 12087 25651 12093
rect 25593 12084 25605 12087
rect 25179 12056 25605 12084
rect 25179 12053 25191 12056
rect 25133 12047 25191 12053
rect 25593 12053 25605 12056
rect 25639 12053 25651 12087
rect 25593 12047 25651 12053
rect 26970 12044 26976 12096
rect 27028 12044 27034 12096
rect 552 11994 31648 12016
rect 552 11942 4285 11994
rect 4337 11942 4349 11994
rect 4401 11942 4413 11994
rect 4465 11942 4477 11994
rect 4529 11942 4541 11994
rect 4593 11942 12059 11994
rect 12111 11942 12123 11994
rect 12175 11942 12187 11994
rect 12239 11942 12251 11994
rect 12303 11942 12315 11994
rect 12367 11942 19833 11994
rect 19885 11942 19897 11994
rect 19949 11942 19961 11994
rect 20013 11942 20025 11994
rect 20077 11942 20089 11994
rect 20141 11942 27607 11994
rect 27659 11942 27671 11994
rect 27723 11942 27735 11994
rect 27787 11942 27799 11994
rect 27851 11942 27863 11994
rect 27915 11942 31648 11994
rect 552 11920 31648 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3418 11880 3424 11892
rect 3016 11852 3424 11880
rect 3016 11840 3022 11852
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 4522 11880 4528 11892
rect 3660 11852 4528 11880
rect 3660 11840 3666 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 5031 11883 5089 11889
rect 5031 11880 5043 11883
rect 4856 11852 5043 11880
rect 4856 11840 4862 11852
rect 5031 11849 5043 11852
rect 5077 11849 5089 11883
rect 5031 11843 5089 11849
rect 7742 11840 7748 11892
rect 7800 11840 7806 11892
rect 9122 11840 9128 11892
rect 9180 11840 9186 11892
rect 9490 11840 9496 11892
rect 9548 11840 9554 11892
rect 9600 11852 10640 11880
rect 3053 11815 3111 11821
rect 3053 11781 3065 11815
rect 3099 11781 3111 11815
rect 3053 11775 3111 11781
rect 842 11636 848 11688
rect 900 11636 906 11688
rect 2866 11636 2872 11688
rect 2924 11636 2930 11688
rect 3068 11676 3096 11775
rect 4430 11772 4436 11824
rect 4488 11812 4494 11824
rect 4816 11812 4844 11840
rect 4488 11784 4844 11812
rect 4488 11772 4494 11784
rect 7374 11772 7380 11824
rect 7432 11812 7438 11824
rect 7469 11815 7527 11821
rect 7469 11812 7481 11815
rect 7432 11784 7481 11812
rect 7432 11772 7438 11784
rect 7469 11781 7481 11784
rect 7515 11812 7527 11815
rect 9600 11812 9628 11852
rect 10612 11824 10640 11852
rect 10778 11840 10784 11892
rect 10836 11840 10842 11892
rect 10962 11840 10968 11892
rect 11020 11840 11026 11892
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11606 11880 11612 11892
rect 11379 11852 11612 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 11940 11852 12265 11880
rect 11940 11840 11946 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 13044 11852 13369 11880
rect 13044 11840 13050 11852
rect 13357 11849 13369 11852
rect 13403 11849 13415 11883
rect 14918 11880 14924 11892
rect 13357 11843 13415 11849
rect 13464 11852 14924 11880
rect 7515 11784 9628 11812
rect 7515 11781 7527 11784
rect 7469 11775 7527 11781
rect 10134 11772 10140 11824
rect 10192 11772 10198 11824
rect 10505 11815 10563 11821
rect 10505 11781 10517 11815
rect 10551 11781 10563 11815
rect 10505 11775 10563 11781
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3510 11744 3516 11756
rect 3283 11716 3516 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3510 11704 3516 11716
rect 3568 11744 3574 11756
rect 3568 11716 5764 11744
rect 3568 11704 3574 11716
rect 5736 11685 5764 11716
rect 5994 11704 6000 11756
rect 6052 11704 6058 11756
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 6420 11716 8493 11744
rect 6420 11704 6426 11716
rect 8481 11713 8493 11716
rect 8527 11744 8539 11747
rect 9030 11744 9036 11756
rect 8527 11716 9036 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9140 11716 9904 11744
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 3068 11648 3617 11676
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 1118 11568 1124 11620
rect 1176 11568 1182 11620
rect 1762 11568 1768 11620
rect 1820 11568 1826 11620
rect 2958 11568 2964 11620
rect 3016 11568 3022 11620
rect 5736 11608 5764 11639
rect 7926 11636 7932 11688
rect 7984 11636 7990 11688
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8846 11676 8852 11688
rect 8067 11648 8852 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 3896 11580 4002 11608
rect 5736 11580 5856 11608
rect 2590 11500 2596 11552
rect 2648 11500 2654 11552
rect 2976 11540 3004 11568
rect 3896 11540 3924 11580
rect 5828 11552 5856 11580
rect 6546 11568 6552 11620
rect 6604 11568 6610 11620
rect 8665 11611 8723 11617
rect 8665 11608 8677 11611
rect 7576 11580 8677 11608
rect 4890 11540 4896 11552
rect 2976 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5810 11500 5816 11552
rect 5868 11500 5874 11552
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 7576 11540 7604 11580
rect 8665 11577 8677 11580
rect 8711 11577 8723 11611
rect 8665 11571 8723 11577
rect 8754 11568 8760 11620
rect 8812 11608 8818 11620
rect 9140 11608 9168 11716
rect 9876 11688 9904 11716
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 8812 11580 9168 11608
rect 9232 11608 9260 11639
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 9364 11648 9505 11676
rect 9364 11636 9370 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 9582 11636 9588 11688
rect 9640 11636 9646 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 9692 11608 9720 11639
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10152 11676 10180 11772
rect 10520 11744 10548 11775
rect 10594 11772 10600 11824
rect 10652 11772 10658 11824
rect 10796 11812 10824 11840
rect 13078 11812 13084 11824
rect 10796 11784 11560 11812
rect 11057 11747 11115 11753
rect 10428 11716 10548 11744
rect 10796 11716 11008 11744
rect 9999 11648 10180 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10226 11636 10232 11688
rect 10284 11636 10290 11688
rect 10428 11685 10456 11716
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10686 11676 10692 11688
rect 10551 11648 10692 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 10796 11685 10824 11716
rect 10980 11688 11008 11716
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11238 11744 11244 11756
rect 11103 11716 11244 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10870 11636 10876 11688
rect 10928 11636 10934 11688
rect 10962 11636 10968 11688
rect 11020 11636 11026 11688
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11330 11676 11336 11688
rect 11195 11648 11336 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11532 11685 11560 11784
rect 11900 11784 12940 11812
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 11900 11744 11928 11784
rect 12912 11756 12940 11784
rect 13004 11784 13084 11812
rect 12710 11744 12716 11756
rect 11848 11716 11928 11744
rect 12084 11716 12716 11744
rect 11848 11704 11854 11716
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 11882 11636 11888 11688
rect 11940 11636 11946 11688
rect 12084 11685 12112 11716
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 12894 11704 12900 11756
rect 12952 11704 12958 11756
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 9232 11580 9444 11608
rect 9692 11580 10333 11608
rect 8812 11568 8818 11580
rect 6880 11512 7604 11540
rect 8205 11543 8263 11549
rect 6880 11500 6886 11512
rect 8205 11509 8217 11543
rect 8251 11540 8263 11543
rect 9030 11540 9036 11552
rect 8251 11512 9036 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9272 11512 9321 11540
rect 9272 11500 9278 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9416 11540 9444 11580
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 12636 11608 12664 11639
rect 10321 11571 10379 11577
rect 10612 11580 12664 11608
rect 12731 11608 12759 11704
rect 12802 11636 12808 11688
rect 12860 11636 12866 11688
rect 13004 11685 13032 11784
rect 13078 11772 13084 11784
rect 13136 11812 13142 11824
rect 13464 11812 13492 11852
rect 14918 11840 14924 11852
rect 14976 11880 14982 11892
rect 15289 11883 15347 11889
rect 15289 11880 15301 11883
rect 14976 11852 15301 11880
rect 14976 11840 14982 11852
rect 15289 11849 15301 11852
rect 15335 11849 15347 11883
rect 15289 11843 15347 11849
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 15562 11880 15568 11892
rect 15519 11852 15568 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 17589 11883 17647 11889
rect 15672 11852 17540 11880
rect 13136 11784 13492 11812
rect 13136 11772 13142 11784
rect 13538 11772 13544 11824
rect 13596 11772 13602 11824
rect 13556 11744 13584 11772
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13556 11716 13829 11744
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 15672 11744 15700 11852
rect 16206 11772 16212 11824
rect 16264 11812 16270 11824
rect 16761 11815 16819 11821
rect 16761 11812 16773 11815
rect 16264 11784 16773 11812
rect 16264 11772 16270 11784
rect 16761 11781 16773 11784
rect 16807 11812 16819 11815
rect 17512 11812 17540 11852
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 17770 11880 17776 11892
rect 17635 11852 17776 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 17862 11840 17868 11892
rect 17920 11840 17926 11892
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18325 11883 18383 11889
rect 18325 11880 18337 11883
rect 18196 11852 18337 11880
rect 18196 11840 18202 11852
rect 18325 11849 18337 11852
rect 18371 11849 18383 11883
rect 20254 11880 20260 11892
rect 18325 11843 18383 11849
rect 18432 11852 20260 11880
rect 18432 11812 18460 11852
rect 20254 11840 20260 11852
rect 20312 11880 20318 11892
rect 21177 11883 21235 11889
rect 20312 11852 21036 11880
rect 20312 11840 20318 11852
rect 20162 11812 20168 11824
rect 16807 11784 17448 11812
rect 17512 11784 18460 11812
rect 18800 11784 20168 11812
rect 16807 11781 16819 11784
rect 16761 11775 16819 11781
rect 14240 11716 15700 11744
rect 14240 11704 14246 11716
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13188 11608 13216 11639
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 16114 11676 16120 11688
rect 15344 11648 16120 11676
rect 15344 11636 15350 11648
rect 12731 11580 13216 11608
rect 9950 11540 9956 11552
rect 9416 11512 9956 11540
rect 9309 11503 9367 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10612 11540 10640 11580
rect 10183 11512 10640 11540
rect 10689 11543 10747 11549
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10689 11509 10701 11543
rect 10735 11540 10747 11543
rect 11514 11540 11520 11552
rect 10735 11512 11520 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 13188 11540 13216 11580
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 15562 11608 15568 11620
rect 13872 11580 14306 11608
rect 15120 11580 15568 11608
rect 13872 11568 13878 11580
rect 15120 11540 15148 11580
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 15764 11617 15792 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16224 11676 16252 11772
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16666 11744 16672 11756
rect 16531 11716 16672 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17420 11744 17448 11784
rect 18800 11756 18828 11784
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 20438 11772 20444 11824
rect 20496 11772 20502 11824
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 20714 11812 20720 11824
rect 20579 11784 20720 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 20806 11772 20812 11824
rect 20864 11772 20870 11824
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 21008 11812 21036 11852
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21358 11880 21364 11892
rect 21223 11852 21364 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 22554 11840 22560 11892
rect 22612 11880 22618 11892
rect 23474 11880 23480 11892
rect 22612 11852 23480 11880
rect 22612 11840 22618 11852
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 23937 11883 23995 11889
rect 23937 11880 23949 11883
rect 23624 11852 23949 11880
rect 23624 11840 23630 11852
rect 23937 11849 23949 11852
rect 23983 11849 23995 11883
rect 23937 11843 23995 11849
rect 24026 11840 24032 11892
rect 24084 11880 24090 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 24084 11852 24593 11880
rect 24084 11840 24090 11852
rect 24581 11849 24593 11852
rect 24627 11849 24639 11883
rect 24581 11843 24639 11849
rect 26743 11883 26801 11889
rect 26743 11849 26755 11883
rect 26789 11880 26801 11883
rect 26878 11880 26884 11892
rect 26789 11852 26884 11880
rect 26789 11849 26801 11852
rect 26743 11843 26801 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 26970 11840 26976 11892
rect 27028 11840 27034 11892
rect 22278 11812 22284 11824
rect 20947 11784 22284 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 22278 11772 22284 11784
rect 22336 11772 22342 11824
rect 18046 11744 18052 11756
rect 16908 11716 17356 11744
rect 17420 11716 18052 11744
rect 16908 11704 16914 11716
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 16224 11648 16313 11676
rect 16301 11645 16313 11648
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16577 11679 16635 11685
rect 16577 11645 16589 11679
rect 16623 11676 16635 11679
rect 16758 11676 16764 11688
rect 16623 11648 16764 11676
rect 16623 11645 16635 11648
rect 16577 11639 16635 11645
rect 15749 11611 15807 11617
rect 15749 11577 15761 11611
rect 15795 11577 15807 11611
rect 15749 11571 15807 11577
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16592 11608 16620 11639
rect 16758 11636 16764 11648
rect 16816 11676 16822 11688
rect 17328 11685 17356 11716
rect 17788 11685 17816 11716
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18432 11716 18705 11744
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16816 11648 17049 11676
rect 16816 11636 16822 11648
rect 17037 11645 17049 11648
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11676 17371 11679
rect 17773 11679 17831 11685
rect 17359 11648 17724 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 16071 11580 16620 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16850 11568 16856 11620
rect 16908 11608 16914 11620
rect 17696 11608 17724 11648
rect 17773 11645 17785 11679
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18322 11676 18328 11688
rect 18003 11648 18328 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18432 11608 18460 11716
rect 18693 11713 18705 11716
rect 18739 11744 18751 11747
rect 18782 11744 18788 11756
rect 18739 11716 18788 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 18892 11716 19104 11744
rect 18892 11688 18920 11716
rect 18506 11636 18512 11688
rect 18564 11636 18570 11688
rect 18874 11636 18880 11688
rect 18932 11636 18938 11688
rect 19076 11685 19104 11716
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19889 11747 19947 11753
rect 19576 11716 19656 11744
rect 19576 11704 19582 11716
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11676 19119 11679
rect 19628 11676 19656 11716
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 20456 11744 20484 11772
rect 19935 11716 20484 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19107 11648 19564 11676
rect 19628 11648 19993 11676
rect 19107 11645 19119 11648
rect 19061 11639 19119 11645
rect 16908 11580 17448 11608
rect 17696 11580 18460 11608
rect 16908 11568 16914 11580
rect 13188 11512 15148 11540
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15436 11512 15669 11540
rect 15436 11500 15442 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 15657 11503 15715 11509
rect 15838 11500 15844 11552
rect 15896 11500 15902 11552
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 15988 11512 16129 11540
rect 15988 11500 15994 11512
rect 16117 11509 16129 11512
rect 16163 11540 16175 11543
rect 16482 11540 16488 11552
rect 16163 11512 16488 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17420 11549 17448 11580
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 18984 11608 19012 11639
rect 18748 11580 19012 11608
rect 18748 11568 18754 11580
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17000 11512 17233 11540
rect 17000 11500 17006 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 18414 11540 18420 11552
rect 17451 11512 18420 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18984 11540 19012 11580
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19429 11611 19487 11617
rect 19429 11608 19441 11611
rect 19392 11580 19441 11608
rect 19392 11568 19398 11580
rect 19429 11577 19441 11580
rect 19475 11577 19487 11611
rect 19536 11608 19564 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20346 11636 20352 11688
rect 20404 11636 20410 11688
rect 20438 11636 20444 11688
rect 20496 11676 20502 11688
rect 20824 11685 20852 11772
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 24949 11747 25007 11753
rect 22244 11716 24532 11744
rect 22244 11704 22250 11716
rect 20990 11685 20996 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20496 11648 20729 11676
rect 20496 11636 20502 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 20981 11679 20996 11685
rect 20981 11645 20993 11679
rect 20981 11639 20996 11645
rect 20990 11636 20996 11639
rect 21048 11636 21054 11688
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21140 11648 21373 11676
rect 21140 11636 21146 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 21450 11636 21456 11688
rect 21508 11676 21514 11688
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 21508 11648 21833 11676
rect 21508 11636 21514 11648
rect 21821 11645 21833 11648
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 22278 11636 22284 11688
rect 22336 11636 22342 11688
rect 24504 11685 24532 11716
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 26988 11744 27016 11840
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 24995 11716 26832 11744
rect 26988 11716 27169 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 26804 11688 26832 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11645 22707 11679
rect 22649 11639 22707 11645
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11645 23259 11679
rect 23201 11639 23259 11645
rect 24489 11679 24547 11685
rect 24489 11645 24501 11679
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 21008 11608 21036 11636
rect 22664 11608 22692 11639
rect 19536 11580 20300 11608
rect 21008 11580 22692 11608
rect 23216 11608 23244 11639
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25317 11679 25375 11685
rect 25317 11676 25329 11679
rect 24912 11648 25329 11676
rect 24912 11636 24918 11648
rect 25317 11645 25329 11648
rect 25363 11645 25375 11679
rect 25317 11639 25375 11645
rect 26786 11636 26792 11688
rect 26844 11676 26850 11688
rect 26881 11679 26939 11685
rect 26881 11676 26893 11679
rect 26844 11648 26893 11676
rect 26844 11636 26850 11648
rect 26881 11645 26893 11648
rect 26927 11645 26939 11679
rect 26881 11639 26939 11645
rect 23290 11608 23296 11620
rect 23216 11580 23296 11608
rect 19429 11571 19487 11577
rect 20272 11549 20300 11580
rect 23290 11568 23296 11580
rect 23348 11568 23354 11620
rect 24213 11611 24271 11617
rect 24213 11577 24225 11611
rect 24259 11608 24271 11611
rect 24302 11608 24308 11620
rect 24259 11580 24308 11608
rect 24259 11577 24271 11580
rect 24213 11571 24271 11577
rect 24302 11568 24308 11580
rect 24360 11568 24366 11620
rect 26326 11568 26332 11620
rect 26384 11608 26390 11620
rect 26384 11580 27646 11608
rect 26384 11568 26390 11580
rect 27540 11552 27568 11580
rect 20165 11543 20223 11549
rect 20165 11540 20177 11543
rect 18984 11512 20177 11540
rect 20165 11509 20177 11512
rect 20211 11509 20223 11543
rect 20165 11503 20223 11509
rect 20257 11543 20315 11549
rect 20257 11509 20269 11543
rect 20303 11509 20315 11543
rect 20257 11503 20315 11509
rect 20898 11500 20904 11552
rect 20956 11540 20962 11552
rect 23382 11540 23388 11552
rect 20956 11512 23388 11540
rect 20956 11500 20962 11512
rect 23382 11500 23388 11512
rect 23440 11540 23446 11552
rect 24762 11540 24768 11552
rect 23440 11512 24768 11540
rect 23440 11500 23446 11512
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 27522 11500 27528 11552
rect 27580 11500 27586 11552
rect 28626 11500 28632 11552
rect 28684 11500 28690 11552
rect 552 11450 31808 11472
rect 552 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 15946 11450
rect 15998 11398 16010 11450
rect 16062 11398 16074 11450
rect 16126 11398 16138 11450
rect 16190 11398 16202 11450
rect 16254 11398 23720 11450
rect 23772 11398 23784 11450
rect 23836 11398 23848 11450
rect 23900 11398 23912 11450
rect 23964 11398 23976 11450
rect 24028 11398 31494 11450
rect 31546 11398 31558 11450
rect 31610 11398 31622 11450
rect 31674 11398 31686 11450
rect 31738 11398 31750 11450
rect 31802 11398 31808 11450
rect 552 11376 31808 11398
rect 1118 11296 1124 11348
rect 1176 11336 1182 11348
rect 1213 11339 1271 11345
rect 1213 11336 1225 11339
rect 1176 11308 1225 11336
rect 1176 11296 1182 11308
rect 1213 11305 1225 11308
rect 1259 11305 1271 11339
rect 1213 11299 1271 11305
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 2924 11308 3249 11336
rect 2924 11296 2930 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 4430 11336 4436 11348
rect 3237 11299 3295 11305
rect 3620 11308 4436 11336
rect 3620 11277 3648 11308
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 4672 11308 4752 11336
rect 4672 11296 4678 11308
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11237 3663 11271
rect 3605 11231 3663 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1443 11172 1716 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1688 11073 1716 11172
rect 2038 11160 2044 11212
rect 2096 11160 2102 11212
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11200 2191 11203
rect 2501 11203 2559 11209
rect 2501 11200 2513 11203
rect 2179 11172 2513 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 2501 11169 2513 11172
rect 2547 11169 2559 11203
rect 2501 11163 2559 11169
rect 2590 11160 2596 11212
rect 2648 11160 2654 11212
rect 4724 11200 4752 11308
rect 5092 11308 5396 11336
rect 5092 11277 5120 11308
rect 5368 11280 5396 11308
rect 8133 11308 9444 11336
rect 5077 11271 5135 11277
rect 5077 11237 5089 11271
rect 5123 11237 5135 11271
rect 5077 11231 5135 11237
rect 5166 11228 5172 11280
rect 5224 11228 5230 11280
rect 5350 11228 5356 11280
rect 5408 11228 5414 11280
rect 6546 11268 6552 11280
rect 5644 11240 6552 11268
rect 5644 11212 5672 11240
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 8133 11268 8161 11308
rect 7484 11240 8161 11268
rect 8849 11271 8907 11277
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4724 11172 4813 11200
rect 4801 11169 4813 11172
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 5266 11203 5324 11209
rect 5266 11200 5278 11203
rect 4948 11172 4993 11200
rect 5046 11172 5278 11200
rect 4948 11160 4954 11172
rect 2314 11092 2320 11144
rect 2372 11092 2378 11144
rect 2608 11132 2636 11160
rect 3053 11135 3111 11141
rect 3053 11132 3065 11135
rect 2608 11104 3065 11132
rect 3053 11101 3065 11104
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 1673 11067 1731 11073
rect 1673 11033 1685 11067
rect 1719 11033 1731 11067
rect 3068 11064 3096 11095
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3697 11135 3755 11141
rect 3697 11132 3709 11135
rect 3476 11104 3709 11132
rect 3476 11092 3482 11104
rect 3697 11101 3709 11104
rect 3743 11101 3755 11135
rect 3697 11095 3755 11101
rect 3878 11092 3884 11144
rect 3936 11092 3942 11144
rect 4890 11064 4896 11076
rect 3068 11036 4896 11064
rect 1673 11027 1731 11033
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 5046 10996 5074 11172
rect 5266 11169 5278 11172
rect 5312 11169 5324 11203
rect 5266 11163 5324 11169
rect 5626 11160 5632 11212
rect 5684 11160 5690 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 7484 11132 7512 11240
rect 7650 11160 7656 11212
rect 7708 11160 7714 11212
rect 7834 11209 7840 11212
rect 7801 11203 7840 11209
rect 7801 11169 7813 11203
rect 7801 11163 7840 11169
rect 7834 11160 7840 11163
rect 7892 11160 7898 11212
rect 7926 11160 7932 11212
rect 7984 11160 7990 11212
rect 8133 11209 8161 11240
rect 8619 11237 8677 11243
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8118 11203 8176 11209
rect 8118 11169 8130 11203
rect 8164 11169 8176 11203
rect 8619 11203 8631 11237
rect 8665 11203 8677 11237
rect 8849 11237 8861 11271
rect 8895 11268 8907 11271
rect 9309 11271 9367 11277
rect 9309 11268 9321 11271
rect 8895 11240 9321 11268
rect 8895 11237 8907 11240
rect 8849 11231 8907 11237
rect 9309 11237 9321 11240
rect 9355 11237 9367 11271
rect 9416 11268 9444 11308
rect 9490 11296 9496 11348
rect 9548 11296 9554 11348
rect 12986 11336 12992 11348
rect 9693 11308 10548 11336
rect 9693 11268 9721 11308
rect 9950 11268 9956 11280
rect 9416 11240 9721 11268
rect 9784 11240 9956 11268
rect 9309 11231 9367 11237
rect 8619 11200 8677 11203
rect 8938 11200 8944 11212
rect 8619 11197 8944 11200
rect 8644 11172 8944 11197
rect 8118 11163 8176 11169
rect 8036 11132 8064 11163
rect 8938 11160 8944 11172
rect 8996 11200 9002 11212
rect 9122 11200 9128 11212
rect 8996 11172 9128 11200
rect 8996 11160 9002 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 9324 11200 9352 11231
rect 9582 11200 9588 11212
rect 9324 11172 9588 11200
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 9784 11209 9812 11240
rect 9950 11228 9956 11240
rect 10008 11268 10014 11280
rect 10321 11271 10379 11277
rect 10321 11268 10333 11271
rect 10008 11240 10333 11268
rect 10008 11228 10014 11240
rect 10321 11237 10333 11240
rect 10367 11237 10379 11271
rect 10321 11231 10379 11237
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 6236 11104 7512 11132
rect 7576 11104 8064 11132
rect 6236 11092 6242 11104
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 5810 11064 5816 11076
rect 5491 11036 5816 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7374 11064 7380 11076
rect 7248 11036 7380 11064
rect 7248 11024 7254 11036
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 4028 10968 5074 10996
rect 4028 10956 4034 10968
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 6070 10999 6128 11005
rect 6070 10996 6082 10999
rect 5592 10968 6082 10996
rect 5592 10956 5598 10968
rect 6070 10965 6082 10968
rect 6116 10965 6128 10999
rect 6070 10959 6128 10965
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 7576 11005 7604 11104
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9916 11104 9965 11132
rect 9916 11092 9922 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 8481 11067 8539 11073
rect 8481 11033 8493 11067
rect 8527 11064 8539 11067
rect 8570 11064 8576 11076
rect 8527 11036 8576 11064
rect 8527 11033 8539 11036
rect 8481 11027 8539 11033
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 8938 11024 8944 11076
rect 8996 11024 9002 11076
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 9585 11067 9643 11073
rect 9585 11064 9597 11067
rect 9272 11036 9597 11064
rect 9272 11024 9278 11036
rect 9585 11033 9597 11036
rect 9631 11033 9643 11067
rect 9585 11027 9643 11033
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10060 11064 10088 11163
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10520 11209 10548 11308
rect 10796 11308 12992 11336
rect 10413 11203 10471 11209
rect 10192 11172 10237 11200
rect 10192 11160 10198 11172
rect 10413 11169 10425 11203
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10510 11203 10568 11209
rect 10510 11169 10522 11203
rect 10556 11200 10568 11203
rect 10686 11200 10692 11212
rect 10556 11172 10692 11200
rect 10556 11169 10568 11172
rect 10510 11163 10568 11169
rect 10428 11132 10456 11163
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10796 11132 10824 11308
rect 12986 11296 12992 11308
rect 13044 11336 13050 11348
rect 13262 11336 13268 11348
rect 13044 11308 13268 11336
rect 13044 11296 13050 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 10965 11271 11023 11277
rect 10965 11237 10977 11271
rect 11011 11268 11023 11271
rect 11054 11268 11060 11280
rect 11011 11240 11060 11268
rect 11011 11237 11023 11240
rect 10965 11231 11023 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11238 11228 11244 11280
rect 11296 11228 11302 11280
rect 11330 11228 11336 11280
rect 11388 11228 11394 11280
rect 11882 11268 11888 11280
rect 11449 11240 11888 11268
rect 11449 11212 11477 11240
rect 11882 11228 11888 11240
rect 11940 11268 11946 11280
rect 12158 11268 12164 11280
rect 11940 11240 12164 11268
rect 11940 11228 11946 11240
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12526 11268 12532 11280
rect 12299 11240 12532 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12710 11228 12716 11280
rect 12768 11228 12774 11280
rect 13740 11268 13768 11299
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 15470 11336 15476 11348
rect 14016 11308 15476 11336
rect 14016 11268 14044 11308
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 15620 11308 17724 11336
rect 15620 11296 15626 11308
rect 14090 11277 14096 11280
rect 13740 11240 14044 11268
rect 14077 11271 14096 11277
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11198 11207 11203
rect 11422 11200 11428 11212
rect 11256 11198 11428 11200
rect 11195 11172 11428 11198
rect 11195 11170 11284 11172
rect 11195 11169 11207 11170
rect 11149 11163 11207 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11698 11160 11704 11212
rect 11756 11160 11762 11212
rect 10428 11104 10824 11132
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11330 11132 11336 11144
rect 11020 11104 11336 11132
rect 11020 11092 11026 11104
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 13740 11132 13768 11240
rect 14077 11237 14089 11271
rect 14077 11231 14096 11237
rect 14090 11228 14096 11231
rect 14148 11228 14154 11280
rect 14274 11228 14280 11280
rect 14332 11228 14338 11280
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11200 14795 11203
rect 14826 11200 14832 11212
rect 14783 11172 14832 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 12308 11104 13768 11132
rect 12308 11092 12314 11104
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 9732 11036 10088 11064
rect 9732 11024 9738 11036
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 10652 11036 10701 11064
rect 10652 11024 10658 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 11992 11064 12020 11092
rect 14660 11076 14688 11163
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15562 11160 15568 11212
rect 15620 11160 15626 11212
rect 16316 11209 16344 11308
rect 17696 11280 17724 11308
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 17828 11308 18460 11336
rect 17828 11296 17834 11308
rect 16574 11228 16580 11280
rect 16632 11268 16638 11280
rect 17313 11271 17371 11277
rect 17313 11268 17325 11271
rect 16632 11240 16804 11268
rect 16632 11228 16638 11240
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 16448 11172 16497 11200
rect 16448 11160 16454 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 14976 11104 15485 11132
rect 14976 11092 14982 11104
rect 11664 11036 12020 11064
rect 11664 11024 11670 11036
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 6880 10968 7573 10996
rect 6880 10956 6886 10968
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 7561 10959 7619 10965
rect 7834 10956 7840 11008
rect 7892 10996 7898 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 7892 10968 8309 10996
rect 7892 10956 7898 10968
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 8297 10959 8355 10965
rect 8665 10999 8723 11005
rect 8665 10965 8677 10999
rect 8711 10996 8723 10999
rect 8956 10996 8984 11024
rect 8711 10968 8984 10996
rect 8711 10965 8723 10968
rect 8665 10959 8723 10965
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9180 10968 9321 10996
rect 9180 10956 9186 10968
rect 9309 10965 9321 10968
rect 9355 10996 9367 10999
rect 10778 10996 10784 11008
rect 9355 10968 10784 10996
rect 9355 10965 9367 10968
rect 9309 10959 9367 10965
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11882 10956 11888 11008
rect 11940 10956 11946 11008
rect 11992 10996 12020 11036
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 14642 11064 14648 11076
rect 13320 11036 14648 11064
rect 13320 11024 13326 11036
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15105 11067 15163 11073
rect 15105 11064 15117 11067
rect 15068 11036 15117 11064
rect 15068 11024 15074 11036
rect 15105 11033 15117 11036
rect 15151 11033 15163 11067
rect 15105 11027 15163 11033
rect 15194 11024 15200 11076
rect 15252 11024 15258 11076
rect 15396 11064 15424 11104
rect 15473 11101 15485 11104
rect 15519 11101 15531 11135
rect 15580 11132 15608 11160
rect 16408 11132 16436 11160
rect 15580 11104 16436 11132
rect 15473 11095 15531 11101
rect 16574 11092 16580 11144
rect 16632 11092 16638 11144
rect 15396 11036 15976 11064
rect 13538 10996 13544 11008
rect 11992 10968 13544 10996
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 14093 10999 14151 11005
rect 14093 10965 14105 10999
rect 14139 10996 14151 10999
rect 15838 10996 15844 11008
rect 14139 10968 15844 10996
rect 14139 10965 14151 10968
rect 14093 10959 14151 10965
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 15948 10996 15976 11036
rect 16114 11024 16120 11076
rect 16172 11024 16178 11076
rect 16684 11064 16712 11163
rect 16776 11132 16804 11240
rect 16868 11240 17325 11268
rect 16868 11209 16896 11240
rect 17313 11237 17325 11240
rect 17359 11237 17371 11271
rect 17313 11231 17371 11237
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 18432 11268 18460 11308
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 18564 11308 19717 11336
rect 18564 11296 18570 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20530 11336 20536 11348
rect 20395 11308 20536 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 21450 11336 21456 11348
rect 20864 11308 21456 11336
rect 20864 11296 20870 11308
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 29730 11296 29736 11348
rect 29788 11296 29794 11348
rect 19794 11268 19800 11280
rect 17736 11240 17908 11268
rect 18432 11240 19800 11268
rect 17736 11228 17742 11240
rect 16853 11203 16911 11209
rect 16853 11169 16865 11203
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 16942 11160 16948 11212
rect 17000 11160 17006 11212
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17144 11132 17172 11163
rect 17770 11160 17776 11212
rect 17828 11160 17834 11212
rect 17880 11209 17908 11240
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 19889 11271 19947 11277
rect 19889 11237 19901 11271
rect 19935 11268 19947 11271
rect 20898 11268 20904 11280
rect 19935 11240 20904 11268
rect 19935 11237 19947 11240
rect 19889 11231 19947 11237
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 21416 11240 22048 11268
rect 21416 11228 21422 11240
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11200 18015 11203
rect 18230 11200 18236 11212
rect 18003 11172 18236 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 18340 11172 18521 11200
rect 17218 11132 17224 11144
rect 16776 11104 17224 11132
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17126 11064 17132 11076
rect 16684 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 17696 11064 17724 11095
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18340 11132 18368 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18966 11160 18972 11212
rect 19024 11160 19030 11212
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 19306 11172 20085 11200
rect 18104 11104 18368 11132
rect 18104 11092 18110 11104
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 19306 11132 19334 11172
rect 20073 11169 20085 11172
rect 20119 11200 20131 11203
rect 20346 11200 20352 11212
rect 20119 11172 20352 11200
rect 20119 11169 20131 11172
rect 20073 11163 20131 11169
rect 20346 11160 20352 11172
rect 20404 11160 20410 11212
rect 20622 11160 20628 11212
rect 20680 11160 20686 11212
rect 21468 11209 21496 11240
rect 21085 11206 21143 11209
rect 21008 11203 21143 11206
rect 21008 11200 21097 11203
rect 20732 11178 21097 11200
rect 20732 11172 21036 11178
rect 18800 11104 19334 11132
rect 19613 11135 19671 11141
rect 18233 11067 18291 11073
rect 18233 11064 18245 11067
rect 17696 11036 18245 11064
rect 18233 11033 18245 11036
rect 18279 11033 18291 11067
rect 18233 11027 18291 11033
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18800 11064 18828 11104
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 19702 11132 19708 11144
rect 19659 11104 19708 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 20732 11132 20760 11172
rect 21085 11169 21097 11178
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11169 21511 11203
rect 21453 11163 21511 11169
rect 21545 11203 21603 11209
rect 21545 11169 21557 11203
rect 21591 11200 21603 11203
rect 21910 11200 21916 11212
rect 21591 11172 21916 11200
rect 21591 11169 21603 11172
rect 21545 11163 21603 11169
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22020 11200 22048 11240
rect 24670 11228 24676 11280
rect 24728 11268 24734 11280
rect 26326 11268 26332 11280
rect 24728 11240 26332 11268
rect 24728 11228 24734 11240
rect 26326 11228 26332 11240
rect 26384 11228 26390 11280
rect 26602 11228 26608 11280
rect 26660 11228 26666 11280
rect 29748 11268 29776 11296
rect 27080 11240 28488 11268
rect 29748 11240 30052 11268
rect 27080 11212 27108 11240
rect 26789 11203 26847 11209
rect 22020 11172 23428 11200
rect 20588 11104 20760 11132
rect 20809 11135 20867 11141
rect 20588 11092 20594 11104
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 22094 11132 22100 11144
rect 20855 11104 22100 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 22066 11092 22100 11104
rect 22152 11092 22158 11144
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23400 11141 23428 11172
rect 26789 11169 26801 11203
rect 26835 11169 26847 11203
rect 26789 11163 26847 11169
rect 23109 11135 23167 11141
rect 23109 11132 23121 11135
rect 23072 11104 23121 11132
rect 23072 11092 23078 11104
rect 23109 11101 23121 11104
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 24118 11092 24124 11144
rect 24176 11092 24182 11144
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 20901 11067 20959 11073
rect 18380 11036 18828 11064
rect 19352 11036 20852 11064
rect 18380 11024 18386 11036
rect 19352 11008 19380 11036
rect 18046 10996 18052 11008
rect 15948 10968 18052 10996
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18141 10999 18199 11005
rect 18141 10965 18153 10999
rect 18187 10996 18199 10999
rect 19150 10996 19156 11008
rect 18187 10968 19156 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 19334 10956 19340 11008
rect 19392 10956 19398 11008
rect 20438 10956 20444 11008
rect 20496 10996 20502 11008
rect 20714 10996 20720 11008
rect 20496 10968 20720 10996
rect 20496 10956 20502 10968
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 20824 10996 20852 11036
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 21726 11064 21732 11076
rect 20947 11036 21732 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 21726 11024 21732 11036
rect 21784 11064 21790 11076
rect 22066 11064 22094 11092
rect 24136 11064 24164 11092
rect 21784 11036 21956 11064
rect 22066 11036 24164 11064
rect 25424 11064 25452 11095
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 26804 11132 26832 11163
rect 26878 11160 26884 11212
rect 26936 11200 26942 11212
rect 26936 11172 27016 11200
rect 26936 11160 26942 11172
rect 26988 11132 27016 11172
rect 27062 11160 27068 11212
rect 27120 11160 27126 11212
rect 28460 11209 28488 11240
rect 27433 11203 27491 11209
rect 27433 11169 27445 11203
rect 27479 11169 27491 11203
rect 27433 11163 27491 11169
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11200 28503 11203
rect 28626 11200 28632 11212
rect 28491 11172 28632 11200
rect 28491 11169 28503 11172
rect 28445 11163 28503 11169
rect 27448 11132 27476 11163
rect 28626 11160 28632 11172
rect 28684 11200 28690 11212
rect 28905 11203 28963 11209
rect 28905 11200 28917 11203
rect 28684 11172 28917 11200
rect 28684 11160 28690 11172
rect 28905 11169 28917 11172
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 29914 11160 29920 11212
rect 29972 11160 29978 11212
rect 30024 11209 30052 11240
rect 30009 11203 30067 11209
rect 30009 11169 30021 11203
rect 30055 11169 30067 11203
rect 30009 11163 30067 11169
rect 26660 11104 26924 11132
rect 26988 11104 27476 11132
rect 27617 11135 27675 11141
rect 26660 11092 26666 11104
rect 26786 11064 26792 11076
rect 25424 11036 26792 11064
rect 21784 11024 21790 11036
rect 21361 10999 21419 11005
rect 21361 10996 21373 10999
rect 20824 10968 21373 10996
rect 21361 10965 21373 10968
rect 21407 10965 21419 10999
rect 21928 10996 21956 11036
rect 26786 11024 26792 11036
rect 26844 11024 26850 11076
rect 26896 11064 26924 11104
rect 27617 11101 27629 11135
rect 27663 11101 27675 11135
rect 27617 11095 27675 11101
rect 27632 11064 27660 11095
rect 28166 11092 28172 11144
rect 28224 11092 28230 11144
rect 26896 11036 27660 11064
rect 22186 10996 22192 11008
rect 21928 10968 22192 10996
rect 21361 10959 21419 10965
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 22922 10956 22928 11008
rect 22980 10996 22986 11008
rect 24670 10996 24676 11008
rect 22980 10968 24676 10996
rect 22980 10956 22986 10968
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 24946 10956 24952 11008
rect 25004 10996 25010 11008
rect 25145 10999 25203 11005
rect 25145 10996 25157 10999
rect 25004 10968 25157 10996
rect 25004 10956 25010 10968
rect 25145 10965 25157 10968
rect 25191 10965 25203 10999
rect 25145 10959 25203 10965
rect 29546 10956 29552 11008
rect 29604 10956 29610 11008
rect 30190 10956 30196 11008
rect 30248 10956 30254 11008
rect 552 10906 31648 10928
rect 552 10854 4285 10906
rect 4337 10854 4349 10906
rect 4401 10854 4413 10906
rect 4465 10854 4477 10906
rect 4529 10854 4541 10906
rect 4593 10854 12059 10906
rect 12111 10854 12123 10906
rect 12175 10854 12187 10906
rect 12239 10854 12251 10906
rect 12303 10854 12315 10906
rect 12367 10854 19833 10906
rect 19885 10854 19897 10906
rect 19949 10854 19961 10906
rect 20013 10854 20025 10906
rect 20077 10854 20089 10906
rect 20141 10854 27607 10906
rect 27659 10854 27671 10906
rect 27723 10854 27735 10906
rect 27787 10854 27799 10906
rect 27851 10854 27863 10906
rect 27915 10854 31648 10906
rect 552 10832 31648 10854
rect 2590 10752 2596 10804
rect 2648 10801 2654 10804
rect 2648 10795 2697 10801
rect 2648 10761 2651 10795
rect 2685 10792 2697 10795
rect 2685 10764 3924 10792
rect 2685 10761 2697 10764
rect 2648 10755 2697 10761
rect 2648 10752 2654 10755
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 3510 10724 3516 10736
rect 2188 10696 3516 10724
rect 2188 10684 2194 10696
rect 3510 10684 3516 10696
rect 3568 10684 3574 10736
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 2148 10656 2176 10684
rect 900 10628 2176 10656
rect 900 10616 906 10628
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 2372 10628 3801 10656
rect 2372 10616 2378 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3896 10656 3924 10764
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4890 10792 4896 10804
rect 4120 10764 4896 10792
rect 4120 10752 4126 10764
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5534 10752 5540 10804
rect 5592 10752 5598 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6917 10795 6975 10801
rect 6917 10792 6929 10795
rect 5960 10764 6929 10792
rect 5960 10752 5966 10764
rect 6917 10761 6929 10764
rect 6963 10792 6975 10795
rect 7466 10792 7472 10804
rect 6963 10764 7472 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 10042 10792 10048 10804
rect 7576 10764 10048 10792
rect 7576 10724 7604 10764
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10192 10764 12388 10792
rect 10192 10752 10198 10764
rect 6288 10696 7604 10724
rect 6288 10668 6316 10696
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 9401 10727 9459 10733
rect 9401 10724 9413 10727
rect 7800 10696 9413 10724
rect 7800 10684 7806 10696
rect 9401 10693 9413 10696
rect 9447 10693 9459 10727
rect 9401 10687 9459 10693
rect 9766 10684 9772 10736
rect 9824 10724 9830 10736
rect 9824 10696 10364 10724
rect 9824 10684 9830 10696
rect 6178 10656 6184 10668
rect 3896 10628 4569 10656
rect 3789 10619 3847 10625
rect 1213 10591 1271 10597
rect 1213 10588 1225 10591
rect 584 10560 1225 10588
rect 584 10520 612 10560
rect 1213 10557 1225 10560
rect 1259 10557 1271 10591
rect 1213 10551 1271 10557
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3804 10588 3832 10619
rect 4062 10588 4068 10600
rect 3007 10560 3280 10588
rect 3804 10560 4068 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 492 10492 612 10520
rect 492 10248 520 10492
rect 1762 10480 1768 10532
rect 1820 10480 1826 10532
rect 2774 10412 2780 10464
rect 2832 10412 2838 10464
rect 3252 10461 3280 10560
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4541 10597 4569 10628
rect 4632 10628 6184 10656
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4212 10560 4445 10588
rect 4212 10548 4218 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4526 10591 4584 10597
rect 4526 10557 4538 10591
rect 4572 10557 4584 10591
rect 4526 10551 4584 10557
rect 3326 10480 3332 10532
rect 3384 10520 3390 10532
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 3384 10492 3617 10520
rect 3384 10480 3390 10492
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 3605 10483 3663 10489
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10421 3295 10455
rect 3237 10415 3295 10421
rect 3694 10412 3700 10464
rect 3752 10412 3758 10464
rect 4632 10452 4660 10628
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 4913 10597 4941 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6270 10616 6276 10668
rect 6328 10616 6334 10668
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 10336 10665 10364 10696
rect 10321 10659 10379 10665
rect 9364 10628 10273 10656
rect 9364 10616 9370 10628
rect 4898 10591 4956 10597
rect 4898 10557 4910 10591
rect 4944 10557 4956 10591
rect 4898 10551 4956 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5997 10591 6055 10597
rect 5399 10560 5672 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 4709 10523 4767 10529
rect 4709 10489 4721 10523
rect 4755 10520 4767 10523
rect 4755 10492 5396 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 5368 10464 5396 10492
rect 4798 10452 4804 10464
rect 4632 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5074 10412 5080 10464
rect 5132 10412 5138 10464
rect 5350 10412 5356 10464
rect 5408 10412 5414 10464
rect 5644 10461 5672 10560
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6822 10588 6828 10600
rect 6043 10560 6828 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6089 10523 6147 10529
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 6932 10520 6960 10616
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 7708 10560 8401 10588
rect 7708 10548 7714 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8482 10591 8540 10597
rect 8482 10557 8494 10591
rect 8528 10557 8540 10591
rect 8482 10551 8540 10557
rect 6135 10492 6960 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 8076 10492 8217 10520
rect 8076 10480 8082 10492
rect 8205 10489 8217 10492
rect 8251 10489 8263 10523
rect 8205 10483 8263 10489
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8496 10452 8524 10551
rect 8754 10548 8760 10600
rect 8812 10548 8818 10600
rect 8938 10597 8944 10600
rect 8895 10591 8944 10597
rect 8895 10557 8907 10591
rect 8941 10557 8944 10591
rect 8895 10551 8944 10557
rect 8938 10548 8944 10551
rect 8996 10548 9002 10600
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 8665 10523 8723 10529
rect 8665 10489 8677 10523
rect 8711 10520 8723 10523
rect 8711 10492 8800 10520
rect 8711 10489 8723 10492
rect 8665 10483 8723 10489
rect 8772 10464 8800 10492
rect 9582 10480 9588 10532
rect 9640 10480 9646 10532
rect 10245 10520 10273 10628
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10560 10628 10609 10656
rect 10560 10616 10566 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 11606 10656 11612 10668
rect 10643 10628 11612 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12360 10665 12388 10764
rect 13170 10752 13176 10804
rect 13228 10752 13234 10804
rect 13538 10752 13544 10804
rect 13596 10792 13602 10804
rect 13722 10792 13728 10804
rect 13596 10764 13728 10792
rect 13596 10752 13602 10764
rect 13722 10752 13728 10764
rect 13780 10792 13786 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 13780 10764 15025 10792
rect 13780 10752 13786 10764
rect 15013 10761 15025 10764
rect 15059 10792 15071 10795
rect 15102 10792 15108 10804
rect 15059 10764 15108 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 16485 10795 16543 10801
rect 16485 10761 16497 10795
rect 16531 10792 16543 10795
rect 16942 10792 16948 10804
rect 16531 10764 16948 10792
rect 16531 10761 16543 10764
rect 16485 10755 16543 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17773 10795 17831 10801
rect 17773 10761 17785 10795
rect 17819 10792 17831 10795
rect 18230 10792 18236 10804
rect 17819 10764 18236 10792
rect 17819 10761 17831 10764
rect 17773 10755 17831 10761
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18690 10792 18696 10804
rect 18555 10764 18696 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19208 10764 19472 10792
rect 19208 10752 19214 10764
rect 14458 10724 14464 10736
rect 12544 10696 14464 10724
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12360 10588 12388 10619
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12544 10665 12572 10696
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 17221 10727 17279 10733
rect 17221 10724 17233 10727
rect 15856 10696 17233 10724
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 12492 10628 12541 10656
rect 12492 10616 12498 10628
rect 12529 10625 12541 10628
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 13262 10656 13268 10668
rect 12759 10628 13268 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15856 10665 15884 10696
rect 17221 10693 17233 10696
rect 17267 10693 17279 10727
rect 19334 10724 19340 10736
rect 17221 10687 17279 10693
rect 17788 10696 19340 10724
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 14792 10628 15853 10656
rect 14792 10616 14798 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 17788 10656 17816 10696
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 17954 10656 17960 10668
rect 15841 10619 15899 10625
rect 16132 10628 17816 10656
rect 17880 10628 17960 10656
rect 14826 10588 14832 10600
rect 12360 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 16132 10597 16160 10628
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 17402 10548 17408 10600
rect 17460 10548 17466 10600
rect 17880 10597 17908 10628
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 19444 10656 19472 10764
rect 20346 10752 20352 10804
rect 20404 10792 20410 10804
rect 21450 10792 21456 10804
rect 20404 10764 21456 10792
rect 20404 10752 20410 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 24213 10795 24271 10801
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24394 10792 24400 10804
rect 24259 10764 24400 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 24578 10752 24584 10804
rect 24636 10752 24642 10804
rect 26510 10684 26516 10736
rect 26568 10684 26574 10736
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 18187 10628 19196 10656
rect 19444 10628 20453 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10557 17923 10591
rect 17865 10551 17923 10557
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 18322 10548 18328 10600
rect 18380 10548 18386 10600
rect 18524 10597 18552 10628
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10588 18751 10591
rect 19058 10588 19064 10600
rect 18739 10560 19064 10588
rect 18739 10557 18751 10560
rect 18693 10551 18751 10557
rect 10873 10523 10931 10529
rect 10873 10520 10885 10523
rect 10245 10492 10885 10520
rect 10873 10489 10885 10492
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 11330 10480 11336 10532
rect 11388 10480 11394 10532
rect 12406 10492 12848 10520
rect 7616 10424 8524 10452
rect 7616 10412 7622 10424
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 9033 10455 9091 10461
rect 9033 10421 9045 10455
rect 9079 10452 9091 10455
rect 9122 10452 9128 10464
rect 9079 10424 9128 10452
rect 9079 10421 9091 10424
rect 9033 10415 9091 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9548 10424 9781 10452
rect 9548 10412 9554 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 9769 10415 9827 10421
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10962 10452 10968 10464
rect 10275 10424 10968 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12406 10452 12434 10492
rect 12820 10461 12848 10492
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 15654 10520 15660 10532
rect 13596 10492 15660 10520
rect 13596 10480 13602 10492
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 16669 10523 16727 10529
rect 16669 10520 16681 10523
rect 15804 10492 16681 10520
rect 15804 10480 15810 10492
rect 16669 10489 16681 10492
rect 16715 10489 16727 10523
rect 18064 10520 18092 10548
rect 18708 10520 18736 10551
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 18064 10492 18736 10520
rect 16669 10483 16727 10489
rect 11848 10424 12434 10452
rect 12805 10455 12863 10461
rect 11848 10412 11854 10424
rect 12805 10421 12817 10455
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 14976 10424 16037 10452
rect 14976 10412 14982 10424
rect 16025 10421 16037 10424
rect 16071 10452 16083 10455
rect 16390 10452 16396 10464
rect 16071 10424 16396 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16632 10424 16773 10452
rect 16632 10412 16638 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 18966 10452 18972 10464
rect 17368 10424 18972 10452
rect 17368 10412 17374 10424
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19168 10452 19196 10628
rect 20441 10625 20453 10628
rect 20487 10625 20499 10659
rect 20441 10619 20499 10625
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 23014 10656 23020 10668
rect 20763 10628 23020 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 23014 10616 23020 10628
rect 23072 10656 23078 10668
rect 23382 10656 23388 10668
rect 23072 10628 23388 10656
rect 23072 10616 23078 10628
rect 23382 10616 23388 10628
rect 23440 10656 23446 10668
rect 23661 10659 23719 10665
rect 23661 10656 23673 10659
rect 23440 10628 23673 10656
rect 23440 10616 23446 10628
rect 23661 10625 23673 10628
rect 23707 10656 23719 10659
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 23707 10628 26341 10656
rect 23707 10625 23719 10628
rect 23661 10619 23719 10625
rect 26329 10625 26341 10628
rect 26375 10656 26387 10659
rect 26786 10656 26792 10668
rect 26375 10628 26792 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 26786 10616 26792 10628
rect 26844 10656 26850 10668
rect 26844 10628 28304 10656
rect 26844 10616 26850 10628
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10557 21603 10591
rect 21545 10551 21603 10557
rect 20162 10520 20168 10532
rect 20010 10492 20168 10520
rect 20162 10480 20168 10492
rect 20220 10520 20226 10532
rect 20220 10492 20668 10520
rect 20220 10480 20226 10492
rect 20640 10464 20668 10492
rect 19518 10452 19524 10464
rect 19168 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 20898 10412 20904 10464
rect 20956 10412 20962 10464
rect 21560 10452 21588 10551
rect 21634 10548 21640 10600
rect 21692 10548 21698 10600
rect 28276 10597 28304 10628
rect 28261 10591 28319 10597
rect 28261 10557 28273 10591
rect 28307 10588 28319 10591
rect 28810 10588 28816 10600
rect 28307 10560 28816 10588
rect 28307 10557 28319 10560
rect 28261 10551 28319 10557
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 29365 10591 29423 10597
rect 29365 10588 29377 10591
rect 29144 10560 29377 10588
rect 29144 10548 29150 10560
rect 29365 10557 29377 10560
rect 29411 10557 29423 10591
rect 29365 10551 29423 10557
rect 29825 10591 29883 10597
rect 29825 10557 29837 10591
rect 29871 10588 29883 10591
rect 30190 10588 30196 10600
rect 29871 10560 30196 10588
rect 29871 10557 29883 10560
rect 29825 10551 29883 10557
rect 22922 10480 22928 10532
rect 22980 10480 22986 10532
rect 23385 10523 23443 10529
rect 23385 10489 23397 10523
rect 23431 10489 23443 10523
rect 23385 10483 23443 10489
rect 23106 10452 23112 10464
rect 21560 10424 23112 10452
rect 23106 10412 23112 10424
rect 23164 10412 23170 10464
rect 23400 10452 23428 10483
rect 23474 10480 23480 10532
rect 23532 10520 23538 10532
rect 23937 10523 23995 10529
rect 23937 10520 23949 10523
rect 23532 10492 23949 10520
rect 23532 10480 23538 10492
rect 23937 10489 23949 10492
rect 23983 10489 23995 10523
rect 25774 10520 25780 10532
rect 23937 10483 23995 10489
rect 24504 10492 24808 10520
rect 25622 10492 25780 10520
rect 24504 10452 24532 10492
rect 23400 10424 24532 10452
rect 24780 10452 24808 10492
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 26050 10480 26056 10532
rect 26108 10480 26114 10532
rect 27522 10480 27528 10532
rect 27580 10520 27586 10532
rect 27580 10492 27660 10520
rect 27580 10480 27586 10492
rect 25682 10452 25688 10464
rect 24780 10424 25688 10452
rect 25682 10412 25688 10424
rect 25740 10412 25746 10464
rect 27632 10452 27660 10492
rect 27706 10480 27712 10532
rect 27764 10520 27770 10532
rect 27985 10523 28043 10529
rect 27985 10520 27997 10523
rect 27764 10492 27997 10520
rect 27764 10480 27770 10492
rect 27985 10489 27997 10492
rect 28031 10489 28043 10523
rect 27985 10483 28043 10489
rect 28994 10480 29000 10532
rect 29052 10480 29058 10532
rect 29012 10452 29040 10480
rect 27632 10424 29040 10452
rect 29380 10452 29408 10551
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 29641 10455 29699 10461
rect 29641 10452 29653 10455
rect 29380 10424 29653 10452
rect 29641 10421 29653 10424
rect 29687 10421 29699 10455
rect 29641 10415 29699 10421
rect 552 10362 31808 10384
rect 552 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 15946 10362
rect 15998 10310 16010 10362
rect 16062 10310 16074 10362
rect 16126 10310 16138 10362
rect 16190 10310 16202 10362
rect 16254 10310 23720 10362
rect 23772 10310 23784 10362
rect 23836 10310 23848 10362
rect 23900 10310 23912 10362
rect 23964 10310 23976 10362
rect 24028 10310 31494 10362
rect 31546 10310 31558 10362
rect 31610 10310 31622 10362
rect 31674 10310 31686 10362
rect 31738 10310 31750 10362
rect 31802 10310 31808 10362
rect 552 10288 31808 10310
rect 1029 10251 1087 10257
rect 1029 10248 1041 10251
rect 492 10220 1041 10248
rect 1029 10217 1041 10220
rect 1075 10217 1087 10251
rect 1029 10211 1087 10217
rect 1305 10251 1363 10257
rect 1305 10217 1317 10251
rect 1351 10217 1363 10251
rect 1305 10211 1363 10217
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 2590 10248 2596 10260
rect 1811 10220 2596 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 1213 10115 1271 10121
rect 1213 10081 1225 10115
rect 1259 10112 1271 10115
rect 1320 10112 1348 10211
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 2774 10248 2780 10260
rect 2746 10208 2780 10248
rect 2832 10208 2838 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3973 10251 4031 10257
rect 3973 10248 3985 10251
rect 3752 10220 3985 10248
rect 3752 10208 3758 10220
rect 3973 10217 3985 10220
rect 4019 10217 4031 10251
rect 3973 10211 4031 10217
rect 4982 10208 4988 10260
rect 5040 10208 5046 10260
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7558 10248 7564 10260
rect 7064 10220 7564 10248
rect 7064 10208 7070 10220
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8294 10208 8300 10260
rect 8352 10208 8358 10260
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9088 10220 9812 10248
rect 9088 10208 9094 10220
rect 2314 10180 2320 10192
rect 1964 10152 2320 10180
rect 1259 10084 1348 10112
rect 1673 10115 1731 10121
rect 1259 10081 1271 10084
rect 1213 10075 1271 10081
rect 1673 10081 1685 10115
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 1688 9976 1716 10075
rect 1964 10053 1992 10152
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10180 2467 10183
rect 2746 10180 2774 10208
rect 5000 10180 5028 10208
rect 2455 10152 2774 10180
rect 4724 10152 5028 10180
rect 2455 10149 2467 10152
rect 2409 10143 2467 10149
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 4724 10121 4752 10152
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 9784 10189 9812 10220
rect 10226 10208 10232 10260
rect 10284 10208 10290 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10468 10220 10977 10248
rect 10468 10208 10474 10220
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 14553 10251 14611 10257
rect 11940 10220 13124 10248
rect 11940 10208 11946 10220
rect 9769 10183 9827 10189
rect 9769 10149 9781 10183
rect 9815 10149 9827 10183
rect 9769 10143 9827 10149
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 12161 10183 12219 10189
rect 10560 10152 11836 10180
rect 10560 10140 10566 10152
rect 4709 10115 4767 10121
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 2774 10044 2780 10056
rect 1949 10007 2007 10013
rect 2240 10016 2780 10044
rect 2240 9976 2268 10016
rect 2774 10004 2780 10016
rect 2832 10044 2838 10056
rect 3418 10044 3424 10056
rect 2832 10016 3424 10044
rect 2832 10004 2838 10016
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 1688 9948 2268 9976
rect 3528 9920 3556 10098
rect 4709 10081 4721 10115
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10081 5043 10115
rect 4985 10075 5043 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5350 10112 5356 10124
rect 5123 10084 5356 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 3927 10016 4537 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 4525 10013 4537 10016
rect 4571 10044 4583 10047
rect 5000 10044 5028 10075
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 7006 10112 7012 10124
rect 6227 10084 7012 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 7006 10072 7012 10084
rect 7064 10112 7070 10124
rect 7064 10084 7604 10112
rect 7064 10072 7070 10084
rect 4571 10016 5028 10044
rect 6365 10047 6423 10053
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7466 10044 7472 10056
rect 6411 10016 7472 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7576 10044 7604 10084
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10134 10112 10140 10124
rect 10091 10084 10140 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 10459 10084 11008 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 7926 10044 7932 10056
rect 7576 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10044 7990 10056
rect 8754 10044 8760 10056
rect 7984 10016 8760 10044
rect 7984 10004 7990 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 10870 10044 10876 10056
rect 10735 10016 10876 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 4890 9936 4896 9988
rect 4948 9976 4954 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 4948 9948 6009 9976
rect 4948 9936 4954 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 3510 9908 3516 9920
rect 1820 9880 3516 9908
rect 1820 9868 1826 9880
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 9950 9908 9956 9920
rect 7432 9880 9956 9908
rect 7432 9868 7438 9880
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10520 9908 10548 10007
rect 10612 9976 10640 10007
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 10980 10044 11008 10084
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11238 10112 11244 10124
rect 11112 10084 11244 10112
rect 11112 10072 11118 10084
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11422 10072 11428 10124
rect 11480 10072 11486 10124
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 11808 10121 11836 10152
rect 12161 10149 12173 10183
rect 12207 10180 12219 10183
rect 12618 10180 12624 10192
rect 12207 10152 12624 10180
rect 12207 10149 12219 10152
rect 12161 10143 12219 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13096 10189 13124 10220
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 14642 10248 14648 10260
rect 14599 10220 14648 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15194 10248 15200 10260
rect 15059 10220 15200 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15381 10251 15439 10257
rect 15381 10217 15393 10251
rect 15427 10248 15439 10251
rect 15427 10220 16804 10248
rect 15427 10217 15439 10220
rect 15381 10211 15439 10217
rect 13081 10183 13139 10189
rect 13081 10149 13093 10183
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 13814 10140 13820 10192
rect 13872 10140 13878 10192
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10180 15531 10183
rect 15746 10180 15752 10192
rect 15519 10152 15752 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12342 10112 12348 10124
rect 12115 10084 12348 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 15488 10112 15516 10143
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 15841 10183 15899 10189
rect 15841 10149 15853 10183
rect 15887 10180 15899 10183
rect 16298 10180 16304 10192
rect 15887 10152 16304 10180
rect 15887 10149 15899 10152
rect 15841 10143 15899 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 16390 10140 16396 10192
rect 16448 10180 16454 10192
rect 16776 10180 16804 10220
rect 16850 10208 16856 10260
rect 16908 10208 16914 10260
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 17862 10248 17868 10260
rect 17359 10220 17868 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18414 10208 18420 10260
rect 18472 10208 18478 10260
rect 18506 10208 18512 10260
rect 18564 10208 18570 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18656 10220 18889 10248
rect 18656 10208 18662 10220
rect 18877 10217 18889 10220
rect 18923 10248 18935 10251
rect 19150 10248 19156 10260
rect 18923 10220 19156 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 19702 10248 19708 10260
rect 19484 10220 19708 10248
rect 19484 10208 19490 10220
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 19904 10220 21312 10248
rect 18432 10180 18460 10208
rect 16448 10152 16528 10180
rect 16776 10152 18460 10180
rect 18524 10180 18552 10208
rect 19904 10189 19932 10220
rect 19061 10183 19119 10189
rect 19061 10180 19073 10183
rect 18524 10152 19073 10180
rect 16448 10140 16454 10152
rect 14148 10084 15516 10112
rect 14148 10072 14154 10084
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 16500 10121 16528 10152
rect 19061 10149 19073 10152
rect 19107 10149 19119 10183
rect 19061 10143 19119 10149
rect 19889 10183 19947 10189
rect 19889 10149 19901 10183
rect 19935 10149 19947 10183
rect 19889 10143 19947 10149
rect 16485 10115 16543 10121
rect 15620 10084 16344 10112
rect 15620 10072 15626 10084
rect 11146 10044 11152 10056
rect 10980 10016 11152 10044
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11348 9976 11376 10007
rect 11532 9976 11560 10072
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 11664 10016 12173 10044
rect 11664 10004 11670 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12584 10016 12817 10044
rect 12584 10004 12590 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 13722 10044 13728 10056
rect 12851 10016 13728 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 14734 10004 14740 10056
rect 14792 10004 14798 10056
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 10612 9948 11560 9976
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12342 9976 12348 9988
rect 11940 9948 12348 9976
rect 11940 9936 11946 9948
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 14476 9976 14504 10004
rect 16224 9976 16252 10007
rect 12544 9948 12941 9976
rect 14476 9948 16252 9976
rect 16316 9976 16344 10084
rect 16485 10081 16497 10115
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 17218 10072 17224 10124
rect 17276 10072 17282 10124
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17368 10084 17417 10112
rect 17368 10072 17374 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10112 17555 10115
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17543 10084 17969 10112
rect 17543 10081 17555 10084
rect 17497 10075 17555 10081
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 17236 10044 17264 10072
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17236 10016 17785 10044
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17972 10044 18000 10075
rect 18046 10072 18052 10124
rect 18104 10072 18110 10124
rect 18230 10072 18236 10124
rect 18288 10072 18294 10124
rect 18417 10115 18475 10121
rect 18417 10081 18429 10115
rect 18463 10112 18475 10115
rect 18693 10115 18751 10121
rect 18693 10112 18705 10115
rect 18463 10084 18705 10112
rect 18463 10081 18475 10084
rect 18417 10075 18475 10081
rect 18693 10081 18705 10084
rect 18739 10112 18751 10115
rect 18874 10112 18880 10124
rect 18739 10084 18880 10112
rect 18739 10081 18751 10084
rect 18693 10075 18751 10081
rect 18432 10044 18460 10075
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19904 10112 19932 10143
rect 20530 10140 20536 10192
rect 20588 10180 20594 10192
rect 20990 10180 20996 10192
rect 20588 10152 20996 10180
rect 20588 10140 20594 10152
rect 20990 10140 20996 10152
rect 21048 10140 21054 10192
rect 21284 10189 21312 10220
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 22646 10248 22652 10260
rect 21692 10220 22652 10248
rect 21692 10208 21698 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 24213 10251 24271 10257
rect 24213 10248 24225 10251
rect 23676 10220 24225 10248
rect 21269 10183 21327 10189
rect 21269 10149 21281 10183
rect 21315 10149 21327 10183
rect 22922 10180 22928 10192
rect 22586 10152 22928 10180
rect 21269 10143 21327 10149
rect 22922 10140 22928 10152
rect 22980 10140 22986 10192
rect 23017 10183 23075 10189
rect 23017 10149 23029 10183
rect 23063 10180 23075 10183
rect 23676 10180 23704 10220
rect 24213 10217 24225 10220
rect 24259 10217 24271 10251
rect 24213 10211 24271 10217
rect 24578 10208 24584 10260
rect 24636 10248 24642 10260
rect 25225 10251 25283 10257
rect 25225 10248 25237 10251
rect 24636 10220 25237 10248
rect 24636 10208 24642 10220
rect 25225 10217 25237 10220
rect 25271 10217 25283 10251
rect 25225 10211 25283 10217
rect 25593 10251 25651 10257
rect 25593 10217 25605 10251
rect 25639 10217 25651 10251
rect 25593 10211 25651 10217
rect 25608 10180 25636 10211
rect 25682 10208 25688 10260
rect 25740 10208 25746 10260
rect 26050 10208 26056 10260
rect 26108 10248 26114 10260
rect 26145 10251 26203 10257
rect 26145 10248 26157 10251
rect 26108 10220 26157 10248
rect 26108 10208 26114 10220
rect 26145 10217 26157 10220
rect 26191 10217 26203 10251
rect 26145 10211 26203 10217
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 26789 10251 26847 10257
rect 26789 10248 26801 10251
rect 26568 10220 26801 10248
rect 26568 10208 26574 10220
rect 26789 10217 26801 10220
rect 26835 10217 26847 10251
rect 26789 10211 26847 10217
rect 27157 10251 27215 10257
rect 27157 10217 27169 10251
rect 27203 10217 27215 10251
rect 27157 10211 27215 10217
rect 27433 10251 27491 10257
rect 27433 10217 27445 10251
rect 27479 10248 27491 10251
rect 27706 10248 27712 10260
rect 27479 10220 27712 10248
rect 27479 10217 27491 10220
rect 27433 10211 27491 10217
rect 23063 10152 23704 10180
rect 23860 10152 24992 10180
rect 25608 10152 26004 10180
rect 23063 10149 23075 10152
rect 23017 10143 23075 10149
rect 23860 10124 23888 10152
rect 19168 10084 19932 10112
rect 20257 10115 20315 10121
rect 17972 10016 18460 10044
rect 17773 10007 17831 10013
rect 17129 9979 17187 9985
rect 17129 9976 17141 9979
rect 16316 9948 17141 9976
rect 11054 9908 11060 9920
rect 10520 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 12544 9908 12572 9948
rect 11204 9880 12572 9908
rect 12621 9911 12679 9917
rect 11204 9868 11210 9880
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 12710 9908 12716 9920
rect 12667 9880 12716 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12913 9908 12941 9948
rect 15562 9908 15568 9920
rect 12913 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 16224 9908 16252 9948
rect 17129 9945 17141 9948
rect 17175 9945 17187 9979
rect 17129 9939 17187 9945
rect 17678 9936 17684 9988
rect 17736 9936 17742 9988
rect 19168 9976 19196 10084
rect 20257 10081 20269 10115
rect 20303 10112 20315 10115
rect 20717 10115 20775 10121
rect 20717 10112 20729 10115
rect 20303 10084 20729 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 20717 10081 20729 10084
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 23293 10115 23351 10121
rect 23293 10081 23305 10115
rect 23339 10112 23351 10115
rect 23382 10112 23388 10124
rect 23339 10084 23388 10112
rect 23339 10081 23351 10084
rect 23293 10075 23351 10081
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19392 10016 19625 10044
rect 19392 10004 19398 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 18064 9948 19196 9976
rect 18064 9908 18092 9948
rect 16224 9880 18092 9908
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 18196 9880 18337 9908
rect 18196 9868 18202 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 18966 9868 18972 9920
rect 19024 9908 19030 9920
rect 19242 9908 19248 9920
rect 19024 9880 19248 9908
rect 19024 9868 19030 9880
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 20272 9908 20300 10075
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 23753 10115 23811 10121
rect 23753 10112 23765 10115
rect 23492 10084 23765 10112
rect 20530 10004 20536 10056
rect 20588 10004 20594 10056
rect 20625 10047 20683 10053
rect 20625 10013 20637 10047
rect 20671 10044 20683 10047
rect 21634 10044 21640 10056
rect 20671 10016 21640 10044
rect 20671 10013 20683 10016
rect 20625 10007 20683 10013
rect 21634 10004 21640 10016
rect 21692 10044 21698 10056
rect 22462 10044 22468 10056
rect 21692 10016 22468 10044
rect 21692 10004 21698 10016
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 22646 10004 22652 10056
rect 22704 10044 22710 10056
rect 23492 10044 23520 10084
rect 23753 10081 23765 10084
rect 23799 10081 23811 10115
rect 23753 10075 23811 10081
rect 22704 10016 23520 10044
rect 23569 10047 23627 10053
rect 22704 10004 22710 10016
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23584 9976 23612 10007
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23768 10044 23796 10075
rect 23842 10072 23848 10124
rect 23900 10072 23906 10124
rect 23934 10072 23940 10124
rect 23992 10112 23998 10124
rect 24397 10115 24455 10121
rect 24397 10112 24409 10115
rect 23992 10084 24409 10112
rect 23992 10072 23998 10084
rect 24397 10081 24409 10084
rect 24443 10081 24455 10115
rect 24397 10075 24455 10081
rect 24489 10115 24547 10121
rect 24489 10081 24501 10115
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 24504 10044 24532 10075
rect 24578 10072 24584 10124
rect 24636 10072 24642 10124
rect 24673 10115 24731 10121
rect 24673 10081 24685 10115
rect 24719 10112 24731 10115
rect 24762 10112 24768 10124
rect 24719 10084 24768 10112
rect 24719 10081 24731 10084
rect 24673 10075 24731 10081
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 24964 10056 24992 10152
rect 25406 10072 25412 10124
rect 25464 10112 25470 10124
rect 25976 10121 26004 10152
rect 25869 10115 25927 10121
rect 25869 10112 25881 10115
rect 25464 10084 25881 10112
rect 25464 10072 25470 10084
rect 25869 10081 25881 10084
rect 25915 10081 25927 10115
rect 25869 10075 25927 10081
rect 25961 10115 26019 10121
rect 25961 10081 25973 10115
rect 26007 10081 26019 10115
rect 27172 10112 27200 10211
rect 27706 10208 27712 10220
rect 27764 10208 27770 10260
rect 28994 10248 29000 10260
rect 28736 10220 29000 10248
rect 28736 10180 28764 10220
rect 28994 10208 29000 10220
rect 29052 10208 29058 10260
rect 28658 10152 28764 10180
rect 28810 10140 28816 10192
rect 28868 10180 28874 10192
rect 28868 10152 29408 10180
rect 28868 10140 28874 10152
rect 29380 10121 29408 10152
rect 29546 10140 29552 10192
rect 29604 10140 29610 10192
rect 27249 10115 27307 10121
rect 27249 10112 27261 10115
rect 27172 10084 27261 10112
rect 25961 10075 26019 10081
rect 27249 10081 27261 10084
rect 27295 10081 27307 10115
rect 27249 10075 27307 10081
rect 29365 10115 29423 10121
rect 29365 10081 29377 10115
rect 29411 10081 29423 10115
rect 29365 10075 29423 10081
rect 23768 10016 24532 10044
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10044 25191 10047
rect 25222 10044 25228 10056
rect 25179 10016 25228 10044
rect 25179 10013 25191 10016
rect 25133 10007 25191 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 26050 10004 26056 10056
rect 26108 10044 26114 10056
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 26108 10016 26525 10044
rect 26108 10004 26114 10016
rect 26513 10013 26525 10016
rect 26559 10044 26571 10047
rect 26602 10044 26608 10056
rect 26559 10016 26608 10044
rect 26559 10013 26571 10016
rect 26513 10007 26571 10013
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 26694 10004 26700 10056
rect 26752 10004 26758 10056
rect 27614 10004 27620 10056
rect 27672 10004 27678 10056
rect 29089 10047 29147 10053
rect 29089 10013 29101 10047
rect 29135 10044 29147 10047
rect 29564 10044 29592 10140
rect 29135 10016 29592 10044
rect 29135 10013 29147 10016
rect 29089 10007 29147 10013
rect 23750 9976 23756 9988
rect 23348 9948 23756 9976
rect 23348 9936 23354 9948
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 24121 9979 24179 9985
rect 24121 9945 24133 9979
rect 24167 9976 24179 9979
rect 25406 9976 25412 9988
rect 24167 9948 25412 9976
rect 24167 9945 24179 9948
rect 24121 9939 24179 9945
rect 25406 9936 25412 9948
rect 25464 9936 25470 9988
rect 19300 9880 20300 9908
rect 21085 9911 21143 9917
rect 19300 9868 19306 9880
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 23934 9908 23940 9920
rect 21131 9880 23940 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 23934 9868 23940 9880
rect 23992 9868 23998 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25866 9908 25872 9920
rect 25004 9880 25872 9908
rect 25004 9868 25010 9880
rect 25866 9868 25872 9880
rect 25924 9868 25930 9920
rect 552 9818 31648 9840
rect 552 9766 4285 9818
rect 4337 9766 4349 9818
rect 4401 9766 4413 9818
rect 4465 9766 4477 9818
rect 4529 9766 4541 9818
rect 4593 9766 12059 9818
rect 12111 9766 12123 9818
rect 12175 9766 12187 9818
rect 12239 9766 12251 9818
rect 12303 9766 12315 9818
rect 12367 9766 19833 9818
rect 19885 9766 19897 9818
rect 19949 9766 19961 9818
rect 20013 9766 20025 9818
rect 20077 9766 20089 9818
rect 20141 9766 27607 9818
rect 27659 9766 27671 9818
rect 27723 9766 27735 9818
rect 27787 9766 27799 9818
rect 27851 9766 27863 9818
rect 27915 9766 31648 9818
rect 552 9744 31648 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 6270 9704 6276 9716
rect 3936 9676 6276 9704
rect 3936 9664 3942 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7006 9664 7012 9716
rect 7064 9664 7070 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8938 9704 8944 9716
rect 8076 9676 8944 9704
rect 8076 9664 8082 9676
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 11514 9704 11520 9716
rect 10980 9676 11520 9704
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 2556 9608 3740 9636
rect 2556 9596 2562 9608
rect 3712 9577 3740 9608
rect 3896 9577 3924 9664
rect 4982 9636 4988 9648
rect 4448 9608 4988 9636
rect 845 9571 903 9577
rect 845 9537 857 9571
rect 891 9568 903 9571
rect 2593 9571 2651 9577
rect 891 9540 2176 9568
rect 891 9537 903 9540
rect 845 9531 903 9537
rect 2148 9512 2176 9540
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3697 9571 3755 9577
rect 2639 9540 3648 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2130 9460 2136 9512
rect 2188 9460 2194 9512
rect 3620 9509 3648 9540
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9500 2927 9503
rect 3605 9503 3663 9509
rect 2915 9472 3280 9500
rect 2915 9469 2927 9472
rect 2869 9463 2927 9469
rect 1121 9435 1179 9441
rect 1121 9401 1133 9435
rect 1167 9401 1179 9435
rect 1121 9395 1179 9401
rect 1136 9364 1164 9395
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 3252 9373 3280 9472
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4448 9500 4476 9608
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 6454 9636 6460 9648
rect 6012 9608 6460 9636
rect 5000 9568 5028 9596
rect 6012 9577 6040 9608
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 6546 9596 6552 9648
rect 6604 9596 6610 9648
rect 5997 9571 6055 9577
rect 5000 9540 5304 9568
rect 3651 9472 4476 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4522 9460 4528 9512
rect 4580 9460 4586 9512
rect 4706 9509 4712 9512
rect 4673 9503 4712 9509
rect 4673 9469 4685 9503
rect 4673 9463 4712 9469
rect 4706 9460 4712 9463
rect 4764 9460 4770 9512
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5031 9503 5089 9509
rect 5031 9469 5043 9503
rect 5077 9500 5089 9503
rect 5166 9500 5172 9512
rect 5077 9472 5172 9500
rect 5077 9469 5089 9472
rect 5031 9463 5089 9469
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 4801 9435 4859 9441
rect 4801 9432 4813 9435
rect 4212 9404 4813 9432
rect 4212 9392 4218 9404
rect 4724 9376 4752 9404
rect 4801 9401 4813 9404
rect 4847 9401 4859 9435
rect 4908 9432 4936 9463
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5276 9500 5304 9540
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 7024 9568 7052 9664
rect 7558 9596 7564 9648
rect 7616 9596 7622 9648
rect 8389 9639 8447 9645
rect 8389 9605 8401 9639
rect 8435 9636 8447 9639
rect 8846 9636 8852 9648
rect 8435 9608 8852 9636
rect 8435 9605 8447 9608
rect 8389 9599 8447 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 10505 9639 10563 9645
rect 10505 9605 10517 9639
rect 10551 9636 10563 9639
rect 10980 9636 11008 9676
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11790 9704 11796 9716
rect 11664 9676 11796 9704
rect 11664 9664 11670 9676
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12032 9676 12664 9704
rect 12032 9664 12038 9676
rect 12526 9636 12532 9648
rect 10551 9608 11008 9636
rect 12268 9608 12532 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 7576 9568 7604 9596
rect 7024 9540 7144 9568
rect 7576 9540 7697 9568
rect 5997 9531 6055 9537
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5276 9472 6101 9500
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 6089 9463 6147 9469
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 7006 9509 7012 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6512 9472 6837 9500
rect 6512 9460 6518 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 6973 9503 7012 9509
rect 6973 9469 6985 9503
rect 6973 9463 7012 9469
rect 7006 9460 7012 9463
rect 7064 9460 7070 9512
rect 7116 9509 7144 9540
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7190 9460 7196 9512
rect 7248 9460 7254 9512
rect 7374 9509 7380 9512
rect 7331 9503 7380 9509
rect 7331 9469 7343 9503
rect 7377 9469 7380 9503
rect 7331 9463 7380 9469
rect 7374 9460 7380 9463
rect 7432 9460 7438 9512
rect 7669 9509 7697 9540
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 7984 9540 8156 9568
rect 7984 9528 7990 9540
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7654 9503 7712 9509
rect 7654 9469 7666 9503
rect 7700 9469 7712 9503
rect 8026 9503 8084 9509
rect 7654 9463 7712 9469
rect 7760 9472 7972 9500
rect 5442 9432 5448 9444
rect 4908 9404 5448 9432
rect 4801 9395 4859 9401
rect 5442 9392 5448 9404
rect 5500 9432 5506 9444
rect 6181 9435 6239 9441
rect 6181 9432 6193 9435
rect 5500 9404 6193 9432
rect 5500 9392 5506 9404
rect 6181 9401 6193 9404
rect 6227 9401 6239 9435
rect 7576 9432 7604 9463
rect 6181 9395 6239 9401
rect 7484 9404 7604 9432
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 1136 9336 2697 9364
rect 2685 9333 2697 9336
rect 2731 9333 2743 9367
rect 2685 9327 2743 9333
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9333 3295 9367
rect 3237 9327 3295 9333
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 7484 9373 7512 9404
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9333 7527 9367
rect 7469 9327 7527 9333
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 7760 9364 7788 9472
rect 7944 9441 7972 9472
rect 8026 9469 8038 9503
rect 8072 9469 8084 9503
rect 8128 9500 8156 9540
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9766 9568 9772 9580
rect 9088 9540 9772 9568
rect 9088 9528 9094 9540
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 8294 9500 8300 9512
rect 8128 9472 8300 9500
rect 8026 9463 8084 9469
rect 7837 9435 7895 9441
rect 7837 9401 7849 9435
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9401 7987 9435
rect 8041 9432 8069 9463
rect 8294 9460 8300 9472
rect 8352 9500 8358 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 8352 9472 8769 9500
rect 8352 9460 8358 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9263 9472 9996 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 8041 9404 8800 9432
rect 7929 9395 7987 9401
rect 7616 9336 7788 9364
rect 7852 9364 7880 9395
rect 8018 9364 8024 9376
rect 7852 9336 8024 9364
rect 7616 9324 7622 9336
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9364 8263 9367
rect 8662 9364 8668 9376
rect 8251 9336 8668 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8772 9364 8800 9404
rect 8846 9392 8852 9444
rect 8904 9392 8910 9444
rect 9398 9392 9404 9444
rect 9456 9392 9462 9444
rect 9585 9435 9643 9441
rect 9585 9401 9597 9435
rect 9631 9432 9643 9435
rect 9858 9432 9864 9444
rect 9631 9404 9864 9432
rect 9631 9401 9643 9404
rect 9585 9395 9643 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 9968 9432 9996 9472
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10520 9500 10548 9599
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 12268 9577 12296 9608
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11664 9540 11989 9568
rect 11664 9528 11670 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12636 9568 12664 9676
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13630 9704 13636 9716
rect 12768 9676 13636 9704
rect 12768 9664 12774 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13722 9664 13728 9716
rect 13780 9664 13786 9716
rect 17313 9707 17371 9713
rect 17313 9673 17325 9707
rect 17359 9704 17371 9707
rect 17402 9704 17408 9716
rect 17359 9676 17408 9704
rect 17359 9673 17371 9676
rect 17313 9667 17371 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 17678 9664 17684 9716
rect 17736 9704 17742 9716
rect 18230 9704 18236 9716
rect 17736 9676 18236 9704
rect 17736 9664 17742 9676
rect 18230 9664 18236 9676
rect 18288 9704 18294 9716
rect 18288 9676 19104 9704
rect 18288 9664 18294 9676
rect 13078 9596 13084 9648
rect 13136 9636 13142 9648
rect 13740 9636 13768 9664
rect 13136 9608 13768 9636
rect 13136 9596 13142 9608
rect 12894 9568 12900 9580
rect 12636 9540 12900 9568
rect 12253 9531 12311 9537
rect 12894 9528 12900 9540
rect 12952 9568 12958 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12952 9540 13185 9568
rect 12952 9528 12958 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9568 13691 9571
rect 13740 9568 13768 9608
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 16390 9636 16396 9648
rect 15764 9608 16396 9636
rect 13679 9540 13768 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 10100 9472 10548 9500
rect 10100 9460 10106 9472
rect 12342 9460 12348 9512
rect 12400 9460 12406 9512
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12584 9472 13308 9500
rect 12584 9460 12590 9472
rect 9968 9404 10732 9432
rect 8938 9364 8944 9376
rect 8772 9336 8944 9364
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10502 9364 10508 9376
rect 10459 9336 10508 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10704 9364 10732 9404
rect 11514 9392 11520 9444
rect 11572 9392 11578 9444
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 13170 9432 13176 9444
rect 11756 9404 12664 9432
rect 11756 9392 11762 9404
rect 11974 9364 11980 9376
rect 10704 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12526 9324 12532 9376
rect 12584 9324 12590 9376
rect 12636 9373 12664 9404
rect 12820 9404 13176 9432
rect 12820 9376 12848 9404
rect 12621 9367 12679 9373
rect 12621 9333 12633 9367
rect 12667 9333 12679 9367
rect 12621 9327 12679 9333
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 12986 9324 12992 9376
rect 13044 9324 13050 9376
rect 13096 9373 13124 9404
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 13081 9367 13139 9373
rect 13081 9333 13093 9367
rect 13127 9333 13139 9367
rect 13280 9364 13308 9472
rect 13648 9432 13676 9531
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14056 9540 15056 9568
rect 14056 9528 14062 9540
rect 15028 9500 15056 9540
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15764 9568 15792 9608
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 16669 9639 16727 9645
rect 16669 9605 16681 9639
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 15436 9540 15792 9568
rect 15436 9528 15442 9540
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 15896 9540 15945 9568
rect 15896 9528 15902 9540
rect 15933 9537 15945 9540
rect 15979 9537 15991 9571
rect 16684 9568 16712 9599
rect 16758 9596 16764 9648
rect 16816 9596 16822 9648
rect 17221 9639 17279 9645
rect 17221 9605 17233 9639
rect 17267 9636 17279 9639
rect 17267 9608 18092 9636
rect 17267 9605 17279 9608
rect 17221 9599 17279 9605
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16684 9540 16865 9568
rect 15933 9531 15991 9537
rect 16853 9537 16865 9540
rect 16899 9568 16911 9571
rect 17586 9568 17592 9580
rect 16899 9540 17592 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 15470 9500 15476 9512
rect 15028 9486 15476 9500
rect 15042 9472 15476 9486
rect 15470 9460 15476 9472
rect 15528 9500 15534 9512
rect 16574 9500 16580 9512
rect 15528 9472 16580 9500
rect 15528 9460 15534 9472
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 17402 9460 17408 9512
rect 17460 9460 17466 9512
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 18064 9509 18092 9608
rect 19076 9568 19104 9676
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 21361 9707 21419 9713
rect 21361 9704 21373 9707
rect 21232 9676 21373 9704
rect 21232 9664 21238 9676
rect 21361 9673 21373 9676
rect 21407 9673 21419 9707
rect 21361 9667 21419 9673
rect 21726 9664 21732 9716
rect 21784 9664 21790 9716
rect 23382 9664 23388 9716
rect 23440 9704 23446 9716
rect 30190 9704 30196 9716
rect 23440 9676 30196 9704
rect 23440 9664 23446 9676
rect 30190 9664 30196 9676
rect 30248 9664 30254 9716
rect 20990 9596 20996 9648
rect 21048 9636 21054 9648
rect 21818 9636 21824 9648
rect 21048 9608 21824 9636
rect 21048 9596 21054 9608
rect 21818 9596 21824 9608
rect 21876 9636 21882 9648
rect 23474 9636 23480 9648
rect 21876 9608 23480 9636
rect 21876 9596 21882 9608
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 23566 9596 23572 9648
rect 23624 9636 23630 9648
rect 23624 9608 24532 9636
rect 23624 9596 23630 9608
rect 19076 9540 24256 9568
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18598 9500 18604 9512
rect 18095 9472 18604 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19076 9509 19104 9540
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 13814 9432 13820 9444
rect 13648 9404 13820 9432
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9432 16175 9435
rect 16298 9432 16304 9444
rect 16163 9404 16304 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 13924 9364 13952 9395
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 18892 9432 18920 9463
rect 19150 9460 19156 9512
rect 19208 9460 19214 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 21284 9509 21312 9540
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19300 9472 19441 9500
rect 19300 9460 19306 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9469 21327 9503
rect 21269 9463 21327 9469
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 23382 9500 23388 9512
rect 22020 9472 23388 9500
rect 22020 9444 22048 9472
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24118 9460 24124 9512
rect 24176 9500 24182 9512
rect 24228 9509 24256 9540
rect 24394 9528 24400 9580
rect 24452 9528 24458 9580
rect 24504 9568 24532 9608
rect 24946 9596 24952 9648
rect 25004 9636 25010 9648
rect 25961 9639 26019 9645
rect 25961 9636 25973 9639
rect 25004 9608 25973 9636
rect 25004 9596 25010 9608
rect 25961 9605 25973 9608
rect 26007 9605 26019 9639
rect 25961 9599 26019 9605
rect 27065 9571 27123 9577
rect 27065 9568 27077 9571
rect 24504 9540 26188 9568
rect 24213 9503 24271 9509
rect 24213 9500 24225 9503
rect 24176 9472 24225 9500
rect 24176 9460 24182 9472
rect 24213 9469 24225 9472
rect 24259 9469 24271 9503
rect 24213 9463 24271 9469
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 24673 9503 24731 9509
rect 24673 9500 24685 9503
rect 24360 9472 24685 9500
rect 24360 9460 24366 9472
rect 24673 9469 24685 9472
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 25682 9460 25688 9512
rect 25740 9460 25746 9512
rect 26160 9509 26188 9540
rect 26252 9540 27077 9568
rect 26145 9503 26203 9509
rect 26145 9469 26157 9503
rect 26191 9469 26203 9503
rect 26145 9463 26203 9469
rect 19610 9432 19616 9444
rect 16448 9404 18828 9432
rect 18892 9404 19616 9432
rect 16448 9392 16454 9404
rect 13280 9336 13952 9364
rect 13081 9327 13139 9333
rect 15378 9324 15384 9376
rect 15436 9324 15442 9376
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16574 9364 16580 9376
rect 16071 9336 16580 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16574 9324 16580 9336
rect 16632 9364 16638 9376
rect 17310 9364 17316 9376
rect 16632 9336 17316 9364
rect 16632 9324 16638 9336
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9364 17647 9367
rect 17770 9364 17776 9376
rect 17635 9336 17776 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 17862 9324 17868 9376
rect 17920 9324 17926 9376
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 18564 9336 18705 9364
rect 18564 9324 18570 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 18800 9364 18828 9404
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 19705 9435 19763 9441
rect 19705 9401 19717 9435
rect 19751 9432 19763 9435
rect 19978 9432 19984 9444
rect 19751 9404 19984 9432
rect 19751 9401 19763 9404
rect 19705 9395 19763 9401
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 20990 9432 20996 9444
rect 20930 9404 20996 9432
rect 20990 9392 20996 9404
rect 21048 9432 21054 9444
rect 22002 9432 22008 9444
rect 21048 9404 22008 9432
rect 21048 9392 21054 9404
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 24949 9435 25007 9441
rect 22480 9404 24348 9432
rect 19334 9364 19340 9376
rect 18800 9336 19340 9364
rect 18693 9327 18751 9333
rect 19334 9324 19340 9336
rect 19392 9364 19398 9376
rect 20530 9364 20536 9376
rect 19392 9336 20536 9364
rect 19392 9324 19398 9336
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 21726 9364 21732 9376
rect 20680 9336 21732 9364
rect 20680 9324 20686 9336
rect 21726 9324 21732 9336
rect 21784 9364 21790 9376
rect 22480 9364 22508 9404
rect 21784 9336 22508 9364
rect 21784 9324 21790 9336
rect 22554 9324 22560 9376
rect 22612 9364 22618 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 22612 9336 23213 9364
rect 22612 9324 22618 9336
rect 23201 9333 23213 9336
rect 23247 9333 23259 9367
rect 23201 9327 23259 9333
rect 23290 9324 23296 9376
rect 23348 9364 23354 9376
rect 24320 9373 24348 9404
rect 24949 9401 24961 9435
rect 24995 9432 25007 9435
rect 25130 9432 25136 9444
rect 24995 9404 25136 9432
rect 24995 9401 25007 9404
rect 24949 9395 25007 9401
rect 25130 9392 25136 9404
rect 25188 9392 25194 9444
rect 25225 9435 25283 9441
rect 25225 9401 25237 9435
rect 25271 9432 25283 9435
rect 25314 9432 25320 9444
rect 25271 9404 25320 9432
rect 25271 9401 25283 9404
rect 25225 9395 25283 9401
rect 25314 9392 25320 9404
rect 25372 9392 25378 9444
rect 25406 9392 25412 9444
rect 25464 9392 25470 9444
rect 25777 9435 25835 9441
rect 25777 9432 25789 9435
rect 25516 9404 25789 9432
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23348 9336 23857 9364
rect 23348 9324 23354 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 24305 9367 24363 9373
rect 24305 9333 24317 9367
rect 24351 9333 24363 9367
rect 24305 9327 24363 9333
rect 24394 9324 24400 9376
rect 24452 9364 24458 9376
rect 25516 9364 25544 9404
rect 25777 9401 25789 9404
rect 25823 9401 25835 9435
rect 25777 9395 25835 9401
rect 25866 9392 25872 9444
rect 25924 9432 25930 9444
rect 26252 9432 26280 9540
rect 27065 9537 27077 9540
rect 27111 9568 27123 9571
rect 28077 9571 28135 9577
rect 28077 9568 28089 9571
rect 27111 9540 28089 9568
rect 27111 9537 27123 9540
rect 27065 9531 27123 9537
rect 28077 9537 28089 9540
rect 28123 9568 28135 9571
rect 28166 9568 28172 9580
rect 28123 9540 28172 9568
rect 28123 9537 28135 9540
rect 28077 9531 28135 9537
rect 28166 9528 28172 9540
rect 28224 9528 28230 9580
rect 28902 9528 28908 9580
rect 28960 9528 28966 9580
rect 26694 9460 26700 9512
rect 26752 9500 26758 9512
rect 27893 9503 27951 9509
rect 27893 9500 27905 9503
rect 26752 9472 27905 9500
rect 26752 9460 26758 9472
rect 27893 9469 27905 9472
rect 27939 9500 27951 9503
rect 28920 9500 28948 9528
rect 27939 9472 28948 9500
rect 27939 9469 27951 9472
rect 27893 9463 27951 9469
rect 27154 9432 27160 9444
rect 25924 9404 26280 9432
rect 26344 9404 27160 9432
rect 25924 9392 25930 9404
rect 26344 9376 26372 9404
rect 24452 9336 25544 9364
rect 25593 9367 25651 9373
rect 24452 9324 24458 9336
rect 25593 9333 25605 9367
rect 25639 9364 25651 9367
rect 26050 9364 26056 9376
rect 25639 9336 26056 9364
rect 25639 9333 25651 9336
rect 25593 9327 25651 9333
rect 26050 9324 26056 9336
rect 26108 9324 26114 9376
rect 26326 9324 26332 9376
rect 26384 9324 26390 9376
rect 26418 9324 26424 9376
rect 26476 9324 26482 9376
rect 26786 9324 26792 9376
rect 26844 9324 26850 9376
rect 26896 9373 26924 9404
rect 27154 9392 27160 9404
rect 27212 9392 27218 9444
rect 26881 9367 26939 9373
rect 26881 9333 26893 9367
rect 26927 9333 26939 9367
rect 26881 9327 26939 9333
rect 27433 9367 27491 9373
rect 27433 9333 27445 9367
rect 27479 9364 27491 9367
rect 27522 9364 27528 9376
rect 27479 9336 27528 9364
rect 27479 9333 27491 9336
rect 27433 9327 27491 9333
rect 27522 9324 27528 9336
rect 27580 9324 27586 9376
rect 27798 9324 27804 9376
rect 27856 9364 27862 9376
rect 28350 9364 28356 9376
rect 27856 9336 28356 9364
rect 27856 9324 27862 9336
rect 28350 9324 28356 9336
rect 28408 9324 28414 9376
rect 552 9274 31808 9296
rect 552 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 15946 9274
rect 15998 9222 16010 9274
rect 16062 9222 16074 9274
rect 16126 9222 16138 9274
rect 16190 9222 16202 9274
rect 16254 9222 23720 9274
rect 23772 9222 23784 9274
rect 23836 9222 23848 9274
rect 23900 9222 23912 9274
rect 23964 9222 23976 9274
rect 24028 9222 31494 9274
rect 31546 9222 31558 9274
rect 31610 9222 31622 9274
rect 31674 9222 31686 9274
rect 31738 9222 31750 9274
rect 31802 9222 31808 9274
rect 552 9200 31808 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 2038 9160 2044 9172
rect 1627 9132 2044 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 2038 9120 2044 9132
rect 2096 9160 2102 9172
rect 2590 9160 2596 9172
rect 2096 9132 2596 9160
rect 2096 9120 2102 9132
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2746 9132 3924 9160
rect 2746 9092 2774 9132
rect 3896 9104 3924 9132
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4580 9132 4721 9160
rect 4580 9120 4586 9132
rect 4709 9129 4721 9132
rect 4755 9129 4767 9163
rect 5534 9160 5540 9172
rect 4709 9123 4767 9129
rect 4816 9132 5540 9160
rect 1504 9064 2774 9092
rect 1504 8965 1532 9064
rect 3878 9052 3884 9104
rect 3936 9052 3942 9104
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8925 1547 8959
rect 1688 8956 1716 8987
rect 2130 8984 2136 9036
rect 2188 8984 2194 9036
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4816 9024 4844 9132
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 4908 9064 5396 9092
rect 4908 9033 4936 9064
rect 3568 8996 4844 9024
rect 4893 9027 4951 9033
rect 3568 8984 3574 8996
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 1688 8928 2176 8956
rect 1489 8919 1547 8925
rect 2038 8780 2044 8832
rect 2096 8780 2102 8832
rect 2148 8820 2176 8928
rect 2406 8916 2412 8968
rect 2464 8916 2470 8968
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8956 3939 8959
rect 4154 8956 4160 8968
rect 3927 8928 4160 8956
rect 3927 8925 3939 8928
rect 3881 8919 3939 8925
rect 4154 8916 4160 8928
rect 4212 8956 4218 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4212 8928 4537 8956
rect 4212 8916 4218 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 4908 8956 4936 8987
rect 4982 8984 4988 9036
rect 5040 8984 5046 9036
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5092 8956 5120 8987
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 5224 8996 5273 9024
rect 5224 8984 5230 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 4856 8928 4936 8956
rect 5000 8928 5120 8956
rect 5368 8956 5396 9064
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5828 9024 5856 9123
rect 7650 9120 7656 9172
rect 7708 9120 7714 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 9226 9163 9284 9169
rect 9226 9160 9238 9163
rect 8536 9132 9238 9160
rect 8536 9120 8542 9132
rect 9226 9129 9238 9132
rect 9272 9129 9284 9163
rect 9226 9123 9284 9129
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6362 9092 6368 9104
rect 6227 9064 6368 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 5583 8996 5856 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 5626 8956 5632 8968
rect 5368 8928 5632 8956
rect 4856 8916 4862 8928
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 4816 8888 4844 8916
rect 3660 8860 4844 8888
rect 5000 8888 5028 8928
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 6196 8888 6224 9055
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 7668 9092 7696 9120
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 6840 9064 7757 9092
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6840 9033 6868 9064
rect 7745 9061 7757 9064
rect 7791 9061 7803 9095
rect 7745 9055 7803 9061
rect 8389 9095 8447 9101
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 8570 9092 8576 9104
rect 8435 9064 8576 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 8757 9095 8815 9101
rect 8757 9061 8769 9095
rect 8803 9092 8815 9095
rect 9030 9092 9036 9104
rect 8803 9064 9036 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9241 9092 9269 9123
rect 9582 9120 9588 9172
rect 9640 9120 9646 9172
rect 10502 9160 10508 9172
rect 9692 9132 10508 9160
rect 9692 9092 9720 9132
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10836 9132 11069 9160
rect 10836 9120 10842 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11057 9123 11115 9129
rect 11238 9120 11244 9172
rect 11296 9120 11302 9172
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 12710 9120 12716 9172
rect 12768 9120 12774 9172
rect 16390 9160 16396 9172
rect 12820 9132 15608 9160
rect 10226 9092 10232 9104
rect 9241 9064 9720 9092
rect 9877 9064 10232 9092
rect 7006 9033 7012 9036
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6512 8996 6837 9024
rect 6512 8984 6518 8996
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 6973 9027 7012 9033
rect 6973 8993 6985 9027
rect 6973 8987 7012 8993
rect 7006 8984 7012 8987
rect 7064 8984 7070 9036
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 7116 8900 7144 8987
rect 7208 8956 7236 8987
rect 7282 8984 7288 9036
rect 7340 9033 7346 9036
rect 7340 9024 7348 9033
rect 7340 8996 7385 9024
rect 7340 8987 7348 8996
rect 7340 8984 7346 8987
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 7650 9024 7656 9036
rect 7524 8996 7656 9024
rect 7524 8984 7530 8996
rect 7650 8984 7656 8996
rect 7708 9024 7714 9036
rect 8849 9027 8907 9033
rect 8849 9024 8861 9027
rect 7708 8996 8861 9024
rect 7708 8984 7714 8996
rect 8849 8993 8861 8996
rect 8895 9024 8907 9027
rect 9877 9024 9905 9064
rect 10226 9052 10232 9064
rect 10284 9092 10290 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 10284 9064 10701 9092
rect 10284 9052 10290 9064
rect 10689 9061 10701 9064
rect 10735 9092 10747 9095
rect 11425 9095 11483 9101
rect 11425 9092 11437 9095
rect 10735 9064 11437 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 11425 9061 11437 9064
rect 11471 9092 11483 9095
rect 12820 9092 12848 9132
rect 15580 9104 15608 9132
rect 15672 9132 16396 9160
rect 11471 9064 12848 9092
rect 11471 9061 11483 9064
rect 11425 9055 11483 9061
rect 14090 9052 14096 9104
rect 14148 9052 14154 9104
rect 15562 9052 15568 9104
rect 15620 9052 15626 9104
rect 8895 9022 9444 9024
rect 9508 9022 9905 9024
rect 8895 8996 9905 9022
rect 10137 9027 10195 9033
rect 8895 8993 8907 8996
rect 9416 8994 9536 8996
rect 8849 8987 8907 8993
rect 10137 8993 10149 9027
rect 10183 9024 10195 9027
rect 10318 9024 10324 9036
rect 10183 8996 10324 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 10318 8984 10324 8996
rect 10376 9024 10382 9036
rect 11146 9024 11152 9036
rect 10376 8996 11152 9024
rect 10376 8984 10382 8996
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 11974 9024 11980 9036
rect 11747 8996 11980 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12308 8996 12817 9024
rect 12308 8984 12314 8996
rect 12805 8993 12817 8996
rect 12851 9024 12863 9027
rect 12986 9024 12992 9036
rect 12851 8996 12992 9024
rect 12851 8993 12863 8996
rect 12805 8987 12863 8993
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 13136 8996 13185 9024
rect 13136 8984 13142 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 7208 8928 9826 8956
rect 6822 8888 6828 8900
rect 5000 8860 6132 8888
rect 6196 8860 6828 8888
rect 3660 8848 3666 8860
rect 5000 8832 5028 8860
rect 3142 8820 3148 8832
rect 2148 8792 3148 8820
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4798 8820 4804 8832
rect 4672 8792 4804 8820
rect 4672 8780 4678 8792
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4982 8780 4988 8832
rect 5040 8780 5046 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5353 8823 5411 8829
rect 5353 8820 5365 8823
rect 5224 8792 5365 8820
rect 5224 8780 5230 8792
rect 5353 8789 5365 8792
rect 5399 8789 5411 8823
rect 6104 8820 6132 8860
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 7098 8848 7104 8900
rect 7156 8848 7162 8900
rect 8018 8888 8024 8900
rect 7392 8860 8024 8888
rect 7392 8820 7420 8860
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8570 8888 8576 8900
rect 8168 8860 8576 8888
rect 8168 8848 8174 8860
rect 8570 8848 8576 8860
rect 8628 8888 8634 8900
rect 8754 8888 8760 8900
rect 8628 8860 8760 8888
rect 8628 8848 8634 8860
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8996 8860 9413 8888
rect 8996 8848 9002 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9798 8888 9826 8928
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 11054 8956 11060 8968
rect 9916 8928 11060 8956
rect 9916 8916 9922 8928
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13906 8956 13912 8968
rect 13596 8928 13912 8956
rect 13596 8916 13602 8928
rect 13906 8916 13912 8928
rect 13964 8956 13970 8968
rect 14921 8959 14979 8965
rect 14921 8956 14933 8959
rect 13964 8928 14933 8956
rect 13964 8916 13970 8928
rect 14921 8925 14933 8928
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15672 8965 15700 9132
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 19889 9163 19947 9169
rect 17828 9132 18092 9160
rect 17828 9120 17834 9132
rect 15749 9095 15807 9101
rect 15749 9061 15761 9095
rect 15795 9092 15807 9095
rect 15795 9064 16252 9092
rect 15795 9061 15807 9064
rect 15749 9055 15807 9061
rect 16224 9033 16252 9064
rect 17034 9052 17040 9104
rect 17092 9052 17098 9104
rect 18064 9101 18092 9132
rect 18524 9132 19334 9160
rect 18049 9095 18107 9101
rect 18049 9061 18061 9095
rect 18095 9061 18107 9095
rect 18049 9055 18107 9061
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15436 8928 15669 8956
rect 15436 8916 15442 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 16224 8956 16252 8987
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 18325 9027 18383 9033
rect 16356 8996 16712 9024
rect 16356 8984 16362 8996
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16224 8928 16589 8956
rect 15841 8919 15899 8925
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 16684 8956 16712 8996
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18414 9024 18420 9036
rect 18371 8996 18420 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18524 9033 18552 9132
rect 19306 9092 19334 9132
rect 19889 9129 19901 9163
rect 19935 9129 19947 9163
rect 19889 9123 19947 9129
rect 19306 9064 19840 9092
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 8993 18567 9027
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 18509 8987 18567 8993
rect 18800 8996 19533 9024
rect 18524 8956 18552 8987
rect 16684 8928 18552 8956
rect 12710 8888 12716 8900
rect 9798 8860 12716 8888
rect 9401 8851 9459 8857
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 12912 8888 12940 8916
rect 13078 8888 13084 8900
rect 12912 8860 13084 8888
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 15856 8888 15884 8919
rect 16684 8888 16712 8928
rect 18598 8916 18604 8968
rect 18656 8956 18662 8968
rect 18800 8965 18828 8996
rect 19521 8993 19533 8996
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 18656 8928 18797 8956
rect 18656 8916 18662 8928
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 19242 8916 19248 8968
rect 19300 8916 19306 8968
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 19702 8956 19708 8968
rect 19475 8928 19708 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 15856 8860 16712 8888
rect 18414 8848 18420 8900
rect 18472 8888 18478 8900
rect 18690 8888 18696 8900
rect 18472 8860 18696 8888
rect 18472 8848 18478 8860
rect 18690 8848 18696 8860
rect 18748 8888 18754 8900
rect 19260 8888 19288 8916
rect 18748 8860 19288 8888
rect 19352 8888 19380 8919
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19812 8956 19840 9064
rect 19904 9024 19932 9123
rect 19978 9120 19984 9172
rect 20036 9120 20042 9172
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 20533 9163 20591 9169
rect 20533 9160 20545 9163
rect 20312 9132 20545 9160
rect 20312 9120 20318 9132
rect 20533 9129 20545 9132
rect 20579 9129 20591 9163
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20533 9123 20591 9129
rect 20732 9132 21281 9160
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 19904 8996 20177 9024
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20732 9024 20760 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 21637 9163 21695 9169
rect 21637 9160 21649 9163
rect 21416 9132 21649 9160
rect 21416 9120 21422 9132
rect 21637 9129 21649 9132
rect 21683 9129 21695 9163
rect 21637 9123 21695 9129
rect 21726 9120 21732 9172
rect 21784 9120 21790 9172
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 24176 9132 24593 9160
rect 24176 9120 24182 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 25593 9163 25651 9169
rect 25593 9129 25605 9163
rect 25639 9160 25651 9163
rect 25958 9160 25964 9172
rect 25639 9132 25964 9160
rect 25639 9129 25651 9132
rect 25593 9123 25651 9129
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26418 9120 26424 9172
rect 26476 9120 26482 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 30101 9163 30159 9169
rect 30101 9160 30113 9163
rect 28408 9132 30113 9160
rect 28408 9120 28414 9132
rect 30101 9129 30113 9132
rect 30147 9129 30159 9163
rect 30101 9123 30159 9129
rect 20993 9095 21051 9101
rect 20993 9061 21005 9095
rect 21039 9092 21051 9095
rect 21174 9092 21180 9104
rect 21039 9064 21180 9092
rect 21039 9061 21051 9064
rect 20993 9055 21051 9061
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 22554 9052 22560 9104
rect 22612 9092 22618 9104
rect 22612 9064 22876 9092
rect 22612 9052 22618 9064
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 20395 8996 20760 9024
rect 20824 8996 22293 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 20717 8959 20775 8965
rect 20717 8956 20729 8959
rect 19812 8928 20729 8956
rect 20717 8925 20729 8928
rect 20763 8956 20775 8959
rect 20824 8956 20852 8996
rect 22281 8993 22293 8996
rect 22327 9024 22339 9027
rect 22370 9024 22376 9036
rect 22327 8996 22376 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 22370 8984 22376 8996
rect 22428 8984 22434 9036
rect 22465 9027 22523 9033
rect 22465 8993 22477 9027
rect 22511 9024 22523 9027
rect 22738 9024 22744 9036
rect 22511 8996 22744 9024
rect 22511 8993 22523 8996
rect 22465 8987 22523 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 22848 9033 22876 9064
rect 23106 9052 23112 9104
rect 23164 9052 23170 9104
rect 24486 9092 24492 9104
rect 24334 9064 24492 9092
rect 24486 9052 24492 9064
rect 24544 9052 24550 9104
rect 24854 9052 24860 9104
rect 24912 9092 24918 9104
rect 25501 9095 25559 9101
rect 25501 9092 25513 9095
rect 24912 9064 25513 9092
rect 24912 9052 24918 9064
rect 25501 9061 25513 9064
rect 25547 9092 25559 9095
rect 25547 9064 26004 9092
rect 25547 9061 25559 9064
rect 25501 9055 25559 9061
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 8993 22891 9027
rect 22833 8987 22891 8993
rect 25041 9027 25099 9033
rect 25041 8993 25053 9027
rect 25087 9024 25099 9027
rect 25087 8996 25176 9024
rect 25087 8993 25099 8996
rect 25041 8987 25099 8993
rect 20763 8928 20852 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 21818 8916 21824 8968
rect 21876 8916 21882 8968
rect 22186 8916 22192 8968
rect 22244 8956 22250 8968
rect 23750 8956 23756 8968
rect 22244 8928 23756 8956
rect 22244 8916 22250 8928
rect 22756 8897 22784 8928
rect 23750 8916 23756 8928
rect 23808 8916 23814 8968
rect 25148 8897 25176 8996
rect 25866 8984 25872 9036
rect 25924 8984 25930 9036
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8956 25835 8959
rect 25884 8956 25912 8984
rect 25823 8928 25912 8956
rect 25976 8956 26004 9064
rect 26053 9027 26111 9033
rect 26053 8993 26065 9027
rect 26099 9024 26111 9027
rect 26436 9024 26464 9120
rect 27430 9052 27436 9104
rect 27488 9052 27494 9104
rect 29086 9052 29092 9104
rect 29144 9052 29150 9104
rect 26099 8996 26464 9024
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 26142 8956 26148 8968
rect 25976 8928 26148 8956
rect 25823 8925 25835 8928
rect 25777 8919 25835 8925
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 27985 8959 28043 8965
rect 27985 8956 27997 8959
rect 26252 8928 27997 8956
rect 26252 8897 26280 8928
rect 27985 8925 27997 8928
rect 28031 8925 28043 8959
rect 28261 8959 28319 8965
rect 28261 8956 28273 8959
rect 27985 8919 28043 8925
rect 28184 8928 28273 8956
rect 22741 8891 22799 8897
rect 19352 8860 19472 8888
rect 18748 8848 18754 8860
rect 6104 8792 7420 8820
rect 5353 8783 5411 8789
rect 7466 8780 7472 8832
rect 7524 8780 7530 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 8444 8792 9229 8820
rect 8444 8780 8450 8792
rect 9217 8789 9229 8792
rect 9263 8820 9275 8823
rect 9490 8820 9496 8832
rect 9263 8792 9496 8820
rect 9263 8789 9275 8792
rect 9217 8783 9275 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9732 8792 9781 8820
rect 9732 8780 9738 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10321 8823 10379 8829
rect 10321 8820 10333 8823
rect 10008 8792 10333 8820
rect 10008 8780 10014 8792
rect 10321 8789 10333 8792
rect 10367 8789 10379 8823
rect 10321 8783 10379 8789
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 10686 8820 10692 8832
rect 10551 8792 10692 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 10686 8780 10692 8792
rect 10744 8820 10750 8832
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 10744 8792 11253 8820
rect 10744 8780 10750 8792
rect 11241 8789 11253 8792
rect 11287 8820 11299 8823
rect 11330 8820 11336 8832
rect 11287 8792 11336 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 11330 8780 11336 8792
rect 11388 8820 11394 8832
rect 15289 8823 15347 8829
rect 15289 8820 15301 8823
rect 11388 8792 15301 8820
rect 11388 8780 11394 8792
rect 15289 8789 15301 8792
rect 15335 8789 15347 8823
rect 15289 8783 15347 8789
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 16758 8820 16764 8832
rect 16448 8792 16764 8820
rect 16448 8780 16454 8792
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 19444 8820 19472 8860
rect 22741 8857 22753 8891
rect 22787 8857 22799 8891
rect 25133 8891 25191 8897
rect 22741 8851 22799 8857
rect 24780 8860 24992 8888
rect 24780 8832 24808 8860
rect 20714 8820 20720 8832
rect 16908 8792 20720 8820
rect 16908 8780 16914 8792
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 24854 8780 24860 8832
rect 24912 8780 24918 8832
rect 24964 8820 24992 8860
rect 25133 8857 25145 8891
rect 25179 8857 25191 8891
rect 25133 8851 25191 8857
rect 26237 8891 26295 8897
rect 26237 8857 26249 8891
rect 26283 8857 26295 8891
rect 26237 8851 26295 8857
rect 26602 8848 26608 8900
rect 26660 8888 26666 8900
rect 26660 8860 27016 8888
rect 26660 8848 26666 8860
rect 26513 8823 26571 8829
rect 26513 8820 26525 8823
rect 24964 8792 26525 8820
rect 26513 8789 26525 8792
rect 26559 8820 26571 8823
rect 26786 8820 26792 8832
rect 26559 8792 26792 8820
rect 26559 8789 26571 8792
rect 26513 8783 26571 8789
rect 26786 8780 26792 8792
rect 26844 8780 26850 8832
rect 26988 8820 27016 8860
rect 28184 8820 28212 8928
rect 28261 8925 28273 8928
rect 28307 8956 28319 8959
rect 28353 8959 28411 8965
rect 28353 8956 28365 8959
rect 28307 8928 28365 8956
rect 28307 8925 28319 8928
rect 28261 8919 28319 8925
rect 28353 8925 28365 8928
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 28626 8916 28632 8968
rect 28684 8916 28690 8968
rect 26988 8792 28212 8820
rect 552 8730 31648 8752
rect 552 8678 4285 8730
rect 4337 8678 4349 8730
rect 4401 8678 4413 8730
rect 4465 8678 4477 8730
rect 4529 8678 4541 8730
rect 4593 8678 12059 8730
rect 12111 8678 12123 8730
rect 12175 8678 12187 8730
rect 12239 8678 12251 8730
rect 12303 8678 12315 8730
rect 12367 8678 19833 8730
rect 19885 8678 19897 8730
rect 19949 8678 19961 8730
rect 20013 8678 20025 8730
rect 20077 8678 20089 8730
rect 20141 8678 27607 8730
rect 27659 8678 27671 8730
rect 27723 8678 27735 8730
rect 27787 8678 27799 8730
rect 27851 8678 27863 8730
rect 27915 8678 31648 8730
rect 552 8656 31648 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2464 8588 2697 8616
rect 2464 8576 2470 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 3160 8588 3648 8616
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 3160 8548 3188 8588
rect 2556 8520 3188 8548
rect 3237 8551 3295 8557
rect 2556 8508 2562 8520
rect 3237 8517 3249 8551
rect 3283 8517 3295 8551
rect 3237 8511 3295 8517
rect 842 8372 848 8424
rect 900 8372 906 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3252 8412 3280 8511
rect 3620 8421 3648 8588
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4890 8616 4896 8628
rect 4304 8588 4896 8616
rect 4304 8576 4310 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5064 8619 5122 8625
rect 5064 8585 5076 8619
rect 5110 8616 5122 8619
rect 5166 8616 5172 8628
rect 5110 8588 5172 8616
rect 5110 8585 5122 8588
rect 5064 8579 5122 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 6328 8588 6653 8616
rect 6328 8576 6334 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7098 8616 7104 8628
rect 6880 8588 7104 8616
rect 6880 8576 6886 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7558 8576 7564 8628
rect 7616 8576 7622 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8018 8616 8024 8628
rect 7975 8588 8024 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 3988 8548 4016 8576
rect 3712 8520 4016 8548
rect 3712 8489 3740 8520
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 2915 8384 3280 8412
rect 3605 8415 3663 8421
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 4172 8412 4200 8576
rect 6549 8551 6607 8557
rect 6549 8517 6561 8551
rect 6595 8548 6607 8551
rect 6595 8520 7328 8548
rect 6595 8517 6607 8520
rect 6549 8511 6607 8517
rect 7300 8489 7328 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 7285 8483 7343 8489
rect 4847 8452 6960 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 6932 8424 6960 8452
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7576 8480 7604 8576
rect 7760 8548 7788 8579
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8386 8576 8392 8628
rect 8444 8576 8450 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 9030 8616 9036 8628
rect 8711 8588 9036 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9306 8576 9312 8628
rect 9364 8576 9370 8628
rect 9858 8576 9864 8628
rect 9916 8576 9922 8628
rect 10226 8616 10232 8628
rect 9968 8588 10232 8616
rect 8404 8548 8432 8576
rect 7760 8520 8432 8548
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8517 8539 8551
rect 9968 8548 9996 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10318 8576 10324 8628
rect 10376 8576 10382 8628
rect 11330 8616 11336 8628
rect 11164 8588 11336 8616
rect 10336 8548 10364 8576
rect 10686 8548 10692 8560
rect 8481 8511 8539 8517
rect 9048 8520 9996 8548
rect 10060 8520 10364 8548
rect 10428 8520 10692 8548
rect 7331 8452 7604 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8496 8480 8524 8511
rect 8444 8452 8524 8480
rect 8444 8440 8450 8452
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8720 8452 8800 8480
rect 8720 8440 8726 8452
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4172 8384 4353 8412
rect 4065 8375 4123 8381
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 1121 8347 1179 8353
rect 1121 8313 1133 8347
rect 1167 8344 1179 8347
rect 1210 8344 1216 8356
rect 1167 8316 1216 8344
rect 1167 8313 1179 8316
rect 1121 8307 1179 8313
rect 1210 8304 1216 8316
rect 1268 8304 1274 8356
rect 2958 8344 2964 8356
rect 2346 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3050 8304 3056 8356
rect 3108 8344 3114 8356
rect 4080 8344 4108 8375
rect 3108 8316 4108 8344
rect 3108 8304 3114 8316
rect 4246 8304 4252 8356
rect 4304 8304 4310 8356
rect 4448 8344 4476 8375
rect 6914 8372 6920 8424
rect 6972 8372 6978 8424
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8412 7435 8415
rect 7650 8412 7656 8424
rect 7423 8384 7656 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 4706 8344 4712 8356
rect 4448 8316 4712 8344
rect 2593 8279 2651 8285
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 3142 8276 3148 8288
rect 2639 8248 3148 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 4448 8276 4476 8316
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5534 8304 5540 8356
rect 5592 8304 5598 8356
rect 7006 8304 7012 8356
rect 7064 8344 7070 8356
rect 7791 8347 7849 8353
rect 7791 8344 7803 8347
rect 7064 8316 7803 8344
rect 7064 8304 7070 8316
rect 7791 8313 7803 8316
rect 7837 8344 7849 8347
rect 8386 8344 8392 8356
rect 7837 8316 8392 8344
rect 7837 8313 7849 8316
rect 7791 8307 7849 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 3476 8248 4476 8276
rect 3476 8236 3482 8248
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5350 8276 5356 8288
rect 5224 8248 5356 8276
rect 5224 8236 5230 8248
rect 5350 8236 5356 8248
rect 5408 8276 5414 8288
rect 6730 8276 6736 8288
rect 5408 8248 6736 8276
rect 5408 8236 5414 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8478 8276 8484 8288
rect 7708 8248 8484 8276
rect 7708 8236 7714 8248
rect 8478 8236 8484 8248
rect 8536 8276 8542 8288
rect 8656 8279 8714 8285
rect 8656 8276 8668 8279
rect 8536 8248 8668 8276
rect 8536 8236 8542 8248
rect 8656 8245 8668 8248
rect 8702 8245 8714 8279
rect 8772 8276 8800 8452
rect 9048 8421 9076 8520
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 10060 8480 10088 8520
rect 10428 8480 10456 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 10873 8551 10931 8557
rect 10873 8517 10885 8551
rect 10919 8548 10931 8551
rect 11164 8548 11192 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12342 8616 12348 8628
rect 11572 8588 12348 8616
rect 11572 8576 11578 8588
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13262 8616 13268 8628
rect 13219 8588 13268 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13403 8588 15056 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13446 8548 13452 8560
rect 10919 8520 11192 8548
rect 12360 8520 13452 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 9723 8452 10088 8480
rect 10152 8452 10456 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9582 8412 9588 8424
rect 9171 8384 9588 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 9950 8412 9956 8424
rect 9824 8384 9956 8412
rect 9824 8372 9830 8384
rect 9950 8372 9956 8384
rect 10008 8412 10014 8424
rect 10152 8412 10180 8452
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 11057 8483 11115 8489
rect 10560 8452 11008 8480
rect 10560 8440 10566 8452
rect 10980 8421 11008 8452
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 11974 8480 11980 8492
rect 11103 8452 11980 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12360 8480 12388 8520
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 12124 8452 12388 8480
rect 12124 8440 12130 8452
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13078 8440 13084 8492
rect 13136 8480 13142 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13136 8452 14105 8480
rect 13136 8440 13142 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10008 8384 10180 8412
rect 10336 8384 10701 8412
rect 10008 8372 10014 8384
rect 10336 8356 10364 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8381 11023 8415
rect 10965 8375 11023 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 13354 8412 13360 8424
rect 13219 8384 13360 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14366 8372 14372 8424
rect 14424 8372 14430 8424
rect 14826 8372 14832 8424
rect 14884 8372 14890 8424
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 15028 8412 15056 8588
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15160 8588 15669 8616
rect 15160 8576 15166 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15804 8588 16037 8616
rect 15804 8576 15810 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16482 8576 16488 8628
rect 16540 8576 16546 8628
rect 16574 8576 16580 8628
rect 16632 8576 16638 8628
rect 17402 8576 17408 8628
rect 17460 8576 17466 8628
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17736 8588 17785 8616
rect 17736 8576 17742 8588
rect 17773 8585 17785 8588
rect 17819 8585 17831 8619
rect 17773 8579 17831 8585
rect 19150 8576 19156 8628
rect 19208 8576 19214 8628
rect 20257 8619 20315 8625
rect 20257 8585 20269 8619
rect 20303 8616 20315 8619
rect 20346 8616 20352 8628
rect 20303 8588 20352 8616
rect 20303 8585 20315 8588
rect 20257 8579 20315 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 21416 8588 22477 8616
rect 21416 8576 21422 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 22833 8619 22891 8625
rect 22833 8585 22845 8619
rect 22879 8616 22891 8619
rect 23106 8616 23112 8628
rect 22879 8588 23112 8616
rect 22879 8585 22891 8588
rect 22833 8579 22891 8585
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23661 8619 23719 8625
rect 23661 8616 23673 8619
rect 23624 8588 23673 8616
rect 23624 8576 23630 8588
rect 23661 8585 23673 8588
rect 23707 8585 23719 8619
rect 23661 8579 23719 8585
rect 23934 8576 23940 8628
rect 23992 8576 23998 8628
rect 24302 8576 24308 8628
rect 24360 8576 24366 8628
rect 24660 8619 24718 8625
rect 24660 8585 24672 8619
rect 24706 8616 24718 8619
rect 24854 8616 24860 8628
rect 24706 8588 24860 8616
rect 24706 8585 24718 8588
rect 24660 8579 24718 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 26142 8576 26148 8628
rect 26200 8576 26206 8628
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26421 8619 26479 8625
rect 26421 8616 26433 8619
rect 26292 8588 26433 8616
rect 26292 8576 26298 8588
rect 26421 8585 26433 8588
rect 26467 8585 26479 8619
rect 26421 8579 26479 8585
rect 15194 8508 15200 8560
rect 15252 8548 15258 8560
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 15252 8520 16129 8548
rect 15252 8508 15258 8520
rect 16117 8517 16129 8520
rect 16163 8517 16175 8551
rect 16592 8548 16620 8576
rect 16117 8511 16175 8517
rect 16408 8520 16620 8548
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 16408 8489 16436 8520
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 16724 8520 18705 8548
rect 16724 8508 16730 8520
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 18693 8511 18751 8517
rect 16393 8483 16451 8489
rect 15344 8452 15884 8480
rect 15344 8440 15350 8452
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15028 8384 15669 8412
rect 14921 8375 14979 8381
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 15856 8412 15884 8452
rect 16393 8449 16405 8483
rect 16439 8449 16451 8483
rect 16393 8443 16451 8449
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 17144 8452 18337 8480
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 15856 8384 16497 8412
rect 15749 8375 15807 8381
rect 16485 8381 16497 8384
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 10229 8347 10287 8353
rect 10229 8313 10241 8347
rect 10275 8313 10287 8347
rect 10229 8307 10287 8313
rect 9306 8276 9312 8288
rect 8772 8248 9312 8276
rect 8656 8239 8714 8245
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10244 8276 10272 8307
rect 10318 8304 10324 8356
rect 10376 8344 10382 8356
rect 10502 8344 10508 8356
rect 10376 8316 10508 8344
rect 10376 8304 10382 8316
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 11330 8304 11336 8356
rect 11388 8304 11394 8356
rect 12710 8344 12716 8356
rect 12558 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 12894 8304 12900 8356
rect 12952 8304 12958 8356
rect 14182 8344 14188 8356
rect 13556 8316 14188 8344
rect 10192 8248 10272 8276
rect 10192 8236 10198 8248
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 12802 8276 12808 8288
rect 10836 8248 12808 8276
rect 10836 8236 10842 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13556 8285 13584 8316
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 14844 8344 14872 8372
rect 14476 8316 14872 8344
rect 14936 8344 14964 8375
rect 14936 8316 15332 8344
rect 13541 8279 13599 8285
rect 13541 8245 13553 8279
rect 13587 8245 13599 8279
rect 13541 8239 13599 8245
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 13906 8276 13912 8288
rect 13688 8248 13912 8276
rect 13688 8236 13694 8248
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 13998 8236 14004 8288
rect 14056 8276 14062 8288
rect 14476 8276 14504 8316
rect 14056 8248 14504 8276
rect 14056 8236 14062 8248
rect 15194 8236 15200 8288
rect 15252 8236 15258 8288
rect 15304 8276 15332 8316
rect 15470 8304 15476 8356
rect 15528 8304 15534 8356
rect 15764 8344 15792 8375
rect 15764 8316 16436 8344
rect 16408 8288 16436 8316
rect 15562 8276 15568 8288
rect 15304 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16390 8236 16396 8288
rect 16448 8236 16454 8288
rect 16500 8276 16528 8375
rect 16758 8372 16764 8424
rect 16816 8412 16822 8424
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16816 8384 17049 8412
rect 16816 8372 16822 8384
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17144 8344 17172 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 17954 8372 17960 8424
rect 18012 8372 18018 8424
rect 18046 8372 18052 8424
rect 18104 8412 18110 8424
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 18104 8384 18889 8412
rect 18104 8372 18110 8384
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 17972 8344 18000 8372
rect 18141 8347 18199 8353
rect 18141 8344 18153 8347
rect 16632 8316 17172 8344
rect 17236 8316 18000 8344
rect 18064 8316 18153 8344
rect 16632 8304 16638 8316
rect 17236 8276 17264 8316
rect 16500 8248 17264 8276
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18064 8276 18092 8316
rect 18141 8313 18153 8316
rect 18187 8313 18199 8347
rect 18141 8307 18199 8313
rect 18233 8347 18291 8353
rect 18233 8313 18245 8347
rect 18279 8344 18291 8347
rect 18414 8344 18420 8356
rect 18279 8316 18420 8344
rect 18279 8313 18291 8316
rect 18233 8307 18291 8313
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 19168 8344 19196 8576
rect 19242 8508 19248 8560
rect 19300 8548 19306 8560
rect 19300 8520 20760 8548
rect 19300 8508 19306 8520
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 19720 8412 19748 8443
rect 19794 8440 19800 8492
rect 19852 8440 19858 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 20732 8489 20760 8520
rect 22572 8520 24440 8548
rect 22572 8492 22600 8520
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8480 20775 8483
rect 22554 8480 22560 8492
rect 20763 8452 22560 8480
rect 20763 8449 20775 8452
rect 20717 8443 20775 8449
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23198 8440 23204 8492
rect 23256 8440 23262 8492
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 24412 8489 24440 8520
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24670 8480 24676 8492
rect 24443 8452 24676 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 26436 8480 26464 8579
rect 27522 8576 27528 8628
rect 27580 8576 27586 8628
rect 27801 8619 27859 8625
rect 27801 8585 27813 8619
rect 27847 8616 27859 8619
rect 28626 8616 28632 8628
rect 27847 8588 28632 8616
rect 27847 8585 27859 8588
rect 27801 8579 27859 8585
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 27430 8508 27436 8560
rect 27488 8508 27494 8560
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26436 8452 26985 8480
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 20456 8412 20484 8440
rect 19720 8384 20484 8412
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22060 8384 22126 8412
rect 22060 8372 22066 8384
rect 22462 8372 22468 8424
rect 22520 8372 22526 8424
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8412 22707 8415
rect 23308 8412 23336 8440
rect 22695 8384 23336 8412
rect 23768 8412 23796 8440
rect 23850 8415 23908 8421
rect 23850 8412 23862 8415
rect 23768 8384 23862 8412
rect 22695 8381 22707 8384
rect 22649 8375 22707 8381
rect 23850 8381 23862 8384
rect 23896 8412 23908 8415
rect 23896 8384 24440 8412
rect 23896 8381 23908 8384
rect 23850 8375 23908 8381
rect 19889 8347 19947 8353
rect 19889 8344 19901 8347
rect 19168 8316 19901 8344
rect 19889 8313 19901 8316
rect 19935 8313 19947 8347
rect 19889 8307 19947 8313
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 20993 8347 21051 8353
rect 20993 8344 21005 8347
rect 20312 8316 21005 8344
rect 20312 8304 20318 8316
rect 20993 8313 21005 8316
rect 21039 8313 21051 8347
rect 22480 8344 22508 8372
rect 23934 8344 23940 8356
rect 22480 8316 23940 8344
rect 20993 8307 21051 8313
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 24412 8344 24440 8384
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 27540 8412 27568 8576
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 26712 8384 27016 8412
rect 27540 8384 27629 8412
rect 26712 8356 26740 8384
rect 24762 8344 24768 8356
rect 24412 8316 24768 8344
rect 24762 8304 24768 8316
rect 24820 8304 24826 8356
rect 26694 8304 26700 8356
rect 26752 8304 26758 8356
rect 26988 8353 27016 8384
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 28077 8415 28135 8421
rect 28077 8381 28089 8415
rect 28123 8412 28135 8415
rect 28166 8412 28172 8424
rect 28123 8384 28172 8412
rect 28123 8381 28135 8384
rect 28077 8375 28135 8381
rect 28166 8372 28172 8384
rect 28224 8372 28230 8424
rect 26881 8347 26939 8353
rect 26881 8313 26893 8347
rect 26927 8313 26939 8347
rect 26881 8307 26939 8313
rect 26973 8347 27031 8353
rect 26973 8313 26985 8347
rect 27019 8313 27031 8347
rect 26973 8307 27031 8313
rect 18012 8248 18092 8276
rect 18012 8236 18018 8248
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 21726 8276 21732 8288
rect 19576 8248 21732 8276
rect 19576 8236 19582 8248
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 23293 8279 23351 8285
rect 23293 8245 23305 8279
rect 23339 8276 23351 8279
rect 23382 8276 23388 8288
rect 23339 8248 23388 8276
rect 23339 8245 23351 8248
rect 23293 8239 23351 8245
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 25314 8276 25320 8288
rect 23624 8248 25320 8276
rect 23624 8236 23630 8248
rect 25314 8236 25320 8248
rect 25372 8276 25378 8288
rect 26896 8276 26924 8307
rect 25372 8248 26924 8276
rect 27893 8279 27951 8285
rect 25372 8236 25378 8248
rect 27893 8245 27905 8279
rect 27939 8276 27951 8279
rect 27982 8276 27988 8288
rect 27939 8248 27988 8276
rect 27939 8245 27951 8248
rect 27893 8239 27951 8245
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 552 8186 31808 8208
rect 552 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 15946 8186
rect 15998 8134 16010 8186
rect 16062 8134 16074 8186
rect 16126 8134 16138 8186
rect 16190 8134 16202 8186
rect 16254 8134 23720 8186
rect 23772 8134 23784 8186
rect 23836 8134 23848 8186
rect 23900 8134 23912 8186
rect 23964 8134 23976 8186
rect 24028 8134 31494 8186
rect 31546 8134 31558 8186
rect 31610 8134 31622 8186
rect 31674 8134 31686 8186
rect 31738 8134 31750 8186
rect 31802 8134 31808 8186
rect 552 8112 31808 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 3694 8072 3700 8084
rect 1636 8044 3700 8072
rect 1636 8032 1642 8044
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 7006 8072 7012 8084
rect 4847 8044 7012 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8846 8072 8852 8084
rect 7616 8044 8852 8072
rect 7616 8032 7622 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 10042 8072 10048 8084
rect 9048 8044 9904 8072
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 2225 8007 2283 8013
rect 2225 8004 2237 8007
rect 1820 7976 2237 8004
rect 1820 7964 1826 7976
rect 2225 7973 2237 7976
rect 2271 7973 2283 8007
rect 7650 8004 7656 8016
rect 2225 7967 2283 7973
rect 4908 7976 7656 8004
rect 1029 7939 1087 7945
rect 1029 7936 1041 7939
rect 768 7908 1041 7936
rect 768 7732 796 7908
rect 1029 7905 1041 7908
rect 1075 7905 1087 7939
rect 1029 7899 1087 7905
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 1305 7939 1363 7945
rect 1305 7936 1317 7939
rect 1176 7908 1317 7936
rect 1176 7896 1182 7908
rect 1305 7905 1317 7908
rect 1351 7905 1363 7939
rect 1305 7899 1363 7905
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1578 7896 1584 7948
rect 1636 7896 1642 7948
rect 4908 7945 4936 7976
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 8352 7976 8585 8004
rect 8352 7964 8358 7976
rect 8573 7973 8585 7976
rect 8619 8004 8631 8007
rect 8619 7976 8708 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 8680 7948 8708 7976
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7905 1731 7939
rect 4893 7939 4951 7945
rect 1673 7899 1731 7905
rect 1688 7812 1716 7899
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 3344 7868 3372 7922
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 4893 7899 4951 7905
rect 5258 7896 5264 7948
rect 5316 7896 5322 7948
rect 5350 7896 5356 7948
rect 5408 7896 5414 7948
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5500 7908 5580 7936
rect 5500 7896 5506 7908
rect 2280 7840 3372 7868
rect 2280 7828 2286 7840
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3697 7871 3755 7877
rect 3697 7868 3709 7871
rect 3568 7840 3709 7868
rect 3568 7828 3574 7840
rect 3697 7837 3709 7840
rect 3743 7868 3755 7871
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 3743 7840 4353 7868
rect 3743 7837 3755 7840
rect 3697 7831 3755 7837
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 5552 7868 5580 7908
rect 5718 7896 5724 7948
rect 5776 7896 5782 7948
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5868 7908 6101 7936
rect 5868 7896 5874 7908
rect 6089 7905 6101 7908
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 6227 7908 6316 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 5552 7840 5641 7868
rect 4341 7831 4399 7837
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5736 7868 5764 7896
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 5736 7840 5917 7868
rect 5629 7831 5687 7837
rect 5905 7837 5917 7840
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 1213 7803 1271 7809
rect 1213 7769 1225 7803
rect 1259 7769 1271 7803
rect 1213 7763 1271 7769
rect 492 7704 796 7732
rect 1228 7732 1256 7763
rect 1670 7760 1676 7812
rect 1728 7760 1734 7812
rect 3970 7800 3976 7812
rect 3712 7772 3976 7800
rect 1762 7732 1768 7744
rect 1228 7704 1768 7732
rect 492 7528 520 7704
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7732 1915 7735
rect 3712 7732 3740 7772
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 5258 7760 5264 7812
rect 5316 7800 5322 7812
rect 6288 7800 6316 7908
rect 6454 7896 6460 7948
rect 6512 7896 6518 7948
rect 6730 7896 6736 7948
rect 6788 7896 6794 7948
rect 6822 7896 6828 7948
rect 6880 7896 6886 7948
rect 7006 7896 7012 7948
rect 7064 7896 7070 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 7116 7868 7144 7899
rect 7374 7868 7380 7880
rect 6411 7840 6914 7868
rect 7116 7840 7380 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 5316 7772 6316 7800
rect 5316 7760 5322 7772
rect 1903 7704 3740 7732
rect 1903 7701 1915 7704
rect 1857 7695 1915 7701
rect 3786 7692 3792 7744
rect 3844 7692 3850 7744
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 4890 7732 4896 7744
rect 4764 7704 4896 7732
rect 4764 7692 4770 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5442 7732 5448 7744
rect 5123 7704 5448 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5718 7732 5724 7744
rect 5583 7704 5724 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5718 7692 5724 7704
rect 5776 7732 5782 7744
rect 6380 7732 6408 7831
rect 6886 7800 6914 7840
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7944 7868 7972 7899
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8076 7908 8401 7936
rect 8076 7896 8082 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 7524 7840 7972 7868
rect 8404 7868 8432 7899
rect 8478 7896 8484 7948
rect 8536 7896 8542 7948
rect 8662 7896 8668 7948
rect 8720 7896 8726 7948
rect 8754 7896 8760 7948
rect 8812 7896 8818 7948
rect 8864 7936 8892 8032
rect 8864 7908 8948 7936
rect 8570 7868 8576 7880
rect 8404 7840 8576 7868
rect 7524 7828 7530 7840
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8920 7868 8948 7908
rect 9048 7868 9076 8044
rect 9876 8013 9904 8044
rect 9968 8044 10048 8072
rect 9968 8013 9996 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 11054 8032 11060 8084
rect 11112 8032 11118 8084
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 12066 8072 12072 8084
rect 11195 8044 12072 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12986 8072 12992 8084
rect 12483 8044 12992 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12986 8032 12992 8044
rect 13044 8072 13050 8084
rect 13170 8072 13176 8084
rect 13044 8044 13176 8072
rect 13044 8032 13050 8044
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 16574 8072 16580 8084
rect 15620 8044 16580 8072
rect 15620 8032 15626 8044
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 24118 8072 24124 8084
rect 16816 8044 24124 8072
rect 16816 8032 16822 8044
rect 24118 8032 24124 8044
rect 24176 8032 24182 8084
rect 24486 8032 24492 8084
rect 24544 8032 24550 8084
rect 24670 8032 24676 8084
rect 24728 8072 24734 8084
rect 25409 8075 25467 8081
rect 24728 8044 25176 8072
rect 24728 8032 24734 8044
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 7973 9919 8007
rect 9861 7967 9919 7973
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 7973 10011 8007
rect 11072 8004 11100 8032
rect 12529 8007 12587 8013
rect 12529 8004 12541 8007
rect 11072 7976 12541 8004
rect 9953 7967 10011 7973
rect 12529 7973 12541 7976
rect 12575 7973 12587 8007
rect 12529 7967 12587 7973
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9306 7936 9312 7948
rect 9263 7908 9312 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 8920 7840 9076 7868
rect 7006 7800 7012 7812
rect 6886 7772 7012 7800
rect 7006 7760 7012 7772
rect 7064 7760 7070 7812
rect 7926 7800 7932 7812
rect 7116 7772 7932 7800
rect 7116 7744 7144 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 9140 7800 9168 7899
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9876 7908 10057 7936
rect 9876 7880 9904 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10045 7899 10103 7905
rect 10244 7908 10517 7936
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 8720 7772 9168 7800
rect 9508 7800 9536 7831
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 9968 7800 9996 7828
rect 10244 7809 10272 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10778 7896 10784 7948
rect 10836 7896 10842 7948
rect 10962 7896 10968 7948
rect 11020 7896 11026 7948
rect 11609 7939 11667 7945
rect 11072 7908 11560 7936
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10686 7868 10692 7880
rect 10376 7840 10692 7868
rect 10376 7828 10382 7840
rect 10686 7828 10692 7840
rect 10744 7868 10750 7880
rect 11072 7868 11100 7908
rect 10744 7840 11100 7868
rect 11532 7868 11560 7908
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 12544 7936 12572 7967
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 12860 7976 13124 8004
rect 12860 7964 12866 7976
rect 12986 7936 12992 7948
rect 11655 7908 12434 7936
rect 12544 7908 12992 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11532 7840 11713 7868
rect 10744 7828 10750 7840
rect 11701 7837 11713 7840
rect 11747 7868 11759 7871
rect 11790 7868 11796 7880
rect 11747 7840 11796 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 9508 7772 9996 7800
rect 10229 7803 10287 7809
rect 8720 7760 8726 7772
rect 10229 7769 10241 7803
rect 10275 7769 10287 7803
rect 10229 7763 10287 7769
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 12069 7803 12127 7809
rect 12069 7800 12081 7803
rect 11112 7772 12081 7800
rect 11112 7760 11118 7772
rect 12069 7769 12081 7772
rect 12115 7769 12127 7803
rect 12406 7800 12434 7908
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 12618 7828 12624 7880
rect 12676 7828 12682 7880
rect 13096 7868 13124 7976
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13412 7908 13645 7936
rect 13412 7896 13418 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 14384 7936 14412 8032
rect 15654 7964 15660 8016
rect 15712 7964 15718 8016
rect 16393 8007 16451 8013
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 16666 8004 16672 8016
rect 16439 7976 16672 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 17034 7964 17040 8016
rect 17092 7964 17098 8016
rect 18966 8004 18972 8016
rect 18340 7976 18972 8004
rect 13863 7908 14412 7936
rect 17604 7908 18184 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 13096 7840 13461 7868
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13648 7868 13676 7899
rect 17604 7880 17632 7908
rect 15286 7868 15292 7880
rect 13648 7840 15292 7868
rect 13449 7831 13507 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 12897 7803 12955 7809
rect 12897 7800 12909 7803
rect 12406 7772 12909 7800
rect 12069 7763 12127 7769
rect 12897 7769 12909 7772
rect 12943 7769 12955 7803
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 12897 7763 12955 7769
rect 13464 7772 14381 7800
rect 13464 7744 13492 7772
rect 14369 7769 14381 7772
rect 14415 7800 14427 7803
rect 16132 7800 16160 7831
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17092 7840 17540 7868
rect 17092 7828 17098 7840
rect 14415 7772 16160 7800
rect 17512 7800 17540 7840
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17736 7840 17877 7868
rect 17736 7828 17742 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 18156 7868 18184 7908
rect 18230 7896 18236 7948
rect 18288 7896 18294 7948
rect 18340 7945 18368 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 19702 8013 19708 8016
rect 19687 8007 19708 8013
rect 19687 7973 19699 8007
rect 19687 7967 19708 7973
rect 19702 7964 19708 7967
rect 19760 7964 19766 8016
rect 20165 8007 20223 8013
rect 20165 7973 20177 8007
rect 20211 7973 20223 8007
rect 20165 7967 20223 7973
rect 20257 8007 20315 8013
rect 20257 7973 20269 8007
rect 20303 8004 20315 8007
rect 20438 8004 20444 8016
rect 20303 7976 20444 8004
rect 20303 7973 20315 7976
rect 20257 7967 20315 7973
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 18509 7939 18567 7945
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18598 7936 18604 7948
rect 18555 7908 18604 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18524 7868 18552 7899
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 19392 7908 19993 7936
rect 19392 7896 19398 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 20180 7936 20208 7967
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 20530 7964 20536 8016
rect 20588 8004 20594 8016
rect 20625 8007 20683 8013
rect 20625 8004 20637 8007
rect 20588 7976 20637 8004
rect 20588 7964 20594 7976
rect 20625 7973 20637 7976
rect 20671 8004 20683 8007
rect 21453 8007 21511 8013
rect 21453 8004 21465 8007
rect 20671 7976 21465 8004
rect 20671 7973 20683 7976
rect 20625 7967 20683 7973
rect 21453 7973 21465 7976
rect 21499 7973 21511 8007
rect 21453 7967 21511 7973
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 22833 8007 22891 8013
rect 22833 8004 22845 8007
rect 22796 7976 22845 8004
rect 22796 7964 22802 7976
rect 22833 7973 22845 7976
rect 22879 8004 22891 8007
rect 23566 8004 23572 8016
rect 22879 7976 23572 8004
rect 22879 7973 22891 7976
rect 22833 7967 22891 7973
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 24504 8004 24532 8032
rect 24426 7976 24532 8004
rect 24857 8007 24915 8013
rect 24857 7973 24869 8007
rect 24903 8004 24915 8007
rect 24946 8004 24952 8016
rect 24903 7976 24952 8004
rect 24903 7973 24915 7976
rect 24857 7967 24915 7973
rect 24946 7964 24952 7976
rect 25004 7964 25010 8016
rect 25148 8004 25176 8044
rect 25409 8041 25421 8075
rect 25455 8072 25467 8075
rect 25682 8072 25688 8084
rect 25455 8044 25688 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 25682 8032 25688 8044
rect 25740 8032 25746 8084
rect 25774 8032 25780 8084
rect 25832 8072 25838 8084
rect 28258 8072 28264 8084
rect 25832 8044 26648 8072
rect 25832 8032 25838 8044
rect 26620 8004 26648 8044
rect 27172 8044 28264 8072
rect 27172 8004 27200 8044
rect 28258 8032 28264 8044
rect 28316 8072 28322 8084
rect 29086 8072 29092 8084
rect 28316 8044 29092 8072
rect 28316 8032 28322 8044
rect 29086 8032 29092 8044
rect 29144 8032 29150 8084
rect 25148 7976 26556 8004
rect 26620 7976 27278 8004
rect 20180 7908 20668 7936
rect 19981 7899 20039 7905
rect 20640 7880 20668 7908
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 21821 7939 21879 7945
rect 21821 7936 21833 7939
rect 21232 7908 21833 7936
rect 21232 7896 21238 7908
rect 21821 7905 21833 7908
rect 21867 7905 21879 7939
rect 21821 7899 21879 7905
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 25148 7945 25176 7976
rect 26528 7948 26556 7976
rect 23017 7939 23075 7945
rect 23017 7905 23029 7939
rect 23063 7905 23075 7939
rect 23017 7899 23075 7905
rect 25133 7939 25191 7945
rect 25133 7905 25145 7939
rect 25179 7905 25191 7939
rect 25133 7899 25191 7905
rect 25225 7939 25283 7945
rect 25225 7905 25237 7939
rect 25271 7905 25283 7939
rect 25225 7899 25283 7905
rect 18156 7840 18552 7868
rect 18969 7871 19027 7877
rect 17865 7831 17923 7837
rect 18969 7837 18981 7871
rect 19015 7868 19027 7871
rect 19058 7868 19064 7880
rect 19015 7840 19064 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19208 7840 20300 7868
rect 19208 7828 19214 7840
rect 20162 7800 20168 7812
rect 17512 7772 20168 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 20272 7800 20300 7840
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21637 7871 21695 7877
rect 21637 7868 21649 7871
rect 21048 7840 21649 7868
rect 21048 7828 21054 7840
rect 21637 7837 21649 7840
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 21968 7840 22569 7868
rect 21968 7828 21974 7840
rect 22557 7837 22569 7840
rect 22603 7868 22615 7871
rect 22922 7868 22928 7880
rect 22603 7840 22928 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 20272 7772 20944 7800
rect 5776 7704 6408 7732
rect 6549 7735 6607 7741
rect 5776 7692 5782 7704
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 6638 7732 6644 7744
rect 6595 7704 6644 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7098 7692 7104 7744
rect 7156 7692 7162 7744
rect 7374 7692 7380 7744
rect 7432 7692 7438 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 8168 7704 8217 7732
rect 8168 7692 8174 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9364 7704 9413 7732
rect 9364 7692 9370 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 9916 7704 10333 7732
rect 9916 7692 9922 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 11238 7692 11244 7744
rect 11296 7692 11302 7744
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 13446 7732 13452 7744
rect 12032 7704 13452 7732
rect 12032 7692 12038 7704
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 13998 7732 14004 7744
rect 13771 7704 14004 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 16482 7692 16488 7744
rect 16540 7732 16546 7744
rect 20714 7732 20720 7744
rect 16540 7704 20720 7732
rect 16540 7692 16546 7704
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 20806 7692 20812 7744
rect 20864 7692 20870 7744
rect 20916 7732 20944 7772
rect 23032 7732 23060 7899
rect 23382 7828 23388 7880
rect 23440 7828 23446 7880
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24394 7868 24400 7880
rect 23900 7840 24400 7868
rect 23900 7828 23906 7840
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 25240 7868 25268 7899
rect 25406 7896 25412 7948
rect 25464 7896 25470 7948
rect 25866 7896 25872 7948
rect 25924 7896 25930 7948
rect 26510 7896 26516 7948
rect 26568 7896 26574 7948
rect 28718 7896 28724 7948
rect 28776 7896 28782 7948
rect 25148 7840 25268 7868
rect 25148 7812 25176 7840
rect 25498 7828 25504 7880
rect 25556 7868 25562 7880
rect 25593 7871 25651 7877
rect 25593 7868 25605 7871
rect 25556 7840 25605 7868
rect 25556 7828 25562 7840
rect 25593 7837 25605 7840
rect 25639 7837 25651 7871
rect 25777 7871 25835 7877
rect 25777 7868 25789 7871
rect 25593 7831 25651 7837
rect 25700 7840 25789 7868
rect 23124 7772 23888 7800
rect 23124 7744 23152 7772
rect 20916 7704 23060 7732
rect 23106 7692 23112 7744
rect 23164 7692 23170 7744
rect 23201 7735 23259 7741
rect 23201 7701 23213 7735
rect 23247 7732 23259 7735
rect 23566 7732 23572 7744
rect 23247 7704 23572 7732
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 23860 7732 23888 7772
rect 25130 7760 25136 7812
rect 25188 7760 25194 7812
rect 25222 7732 25228 7744
rect 23860 7704 25228 7732
rect 25222 7692 25228 7704
rect 25280 7732 25286 7744
rect 25700 7732 25728 7840
rect 25777 7837 25789 7840
rect 25823 7837 25835 7871
rect 25777 7831 25835 7837
rect 26789 7871 26847 7877
rect 26789 7837 26801 7871
rect 26835 7868 26847 7871
rect 28074 7868 28080 7880
rect 26835 7840 28080 7868
rect 26835 7837 26847 7840
rect 26789 7831 26847 7837
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7868 28319 7871
rect 28736 7868 28764 7896
rect 28307 7840 28764 7868
rect 28307 7837 28319 7840
rect 28261 7831 28319 7837
rect 28350 7760 28356 7812
rect 28408 7800 28414 7812
rect 28445 7803 28503 7809
rect 28445 7800 28457 7803
rect 28408 7772 28457 7800
rect 28408 7760 28414 7772
rect 28445 7769 28457 7772
rect 28491 7769 28503 7803
rect 28445 7763 28503 7769
rect 25280 7704 25728 7732
rect 26237 7735 26295 7741
rect 25280 7692 25286 7704
rect 26237 7701 26249 7735
rect 26283 7732 26295 7735
rect 28534 7732 28540 7744
rect 26283 7704 28540 7732
rect 26283 7701 26295 7704
rect 26237 7695 26295 7701
rect 28534 7692 28540 7704
rect 28592 7692 28598 7744
rect 552 7642 31648 7664
rect 552 7590 4285 7642
rect 4337 7590 4349 7642
rect 4401 7590 4413 7642
rect 4465 7590 4477 7642
rect 4529 7590 4541 7642
rect 4593 7590 12059 7642
rect 12111 7590 12123 7642
rect 12175 7590 12187 7642
rect 12239 7590 12251 7642
rect 12303 7590 12315 7642
rect 12367 7590 19833 7642
rect 19885 7590 19897 7642
rect 19949 7590 19961 7642
rect 20013 7590 20025 7642
rect 20077 7590 20089 7642
rect 20141 7590 27607 7642
rect 27659 7590 27671 7642
rect 27723 7590 27735 7642
rect 27787 7590 27799 7642
rect 27851 7590 27863 7642
rect 27915 7590 31648 7642
rect 552 7568 31648 7590
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 492 7500 3249 7528
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 3786 7488 3792 7540
rect 3844 7488 3850 7540
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5721 7531 5779 7537
rect 4948 7500 5488 7528
rect 4948 7488 4954 7500
rect 2685 7463 2743 7469
rect 2685 7460 2697 7463
rect 2148 7432 2697 7460
rect 1210 7352 1216 7404
rect 1268 7392 1274 7404
rect 2148 7392 2176 7432
rect 2685 7429 2697 7432
rect 2731 7429 2743 7463
rect 2685 7423 2743 7429
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 2958 7460 2964 7472
rect 2832 7432 2964 7460
rect 2832 7420 2838 7432
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3804 7460 3832 7488
rect 3712 7432 3832 7460
rect 3712 7401 3740 7432
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 5460 7460 5488 7500
rect 5721 7497 5733 7531
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 5736 7460 5764 7491
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5960 7500 6377 7528
rect 5960 7488 5966 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6549 7531 6607 7537
rect 6549 7497 6561 7531
rect 6595 7528 6607 7531
rect 6730 7528 6736 7540
rect 6595 7500 6736 7528
rect 6595 7497 6607 7500
rect 6549 7491 6607 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 9306 7528 9312 7540
rect 7064 7500 9312 7528
rect 7064 7488 7070 7500
rect 9306 7488 9312 7500
rect 9364 7528 9370 7540
rect 9677 7531 9735 7537
rect 9364 7500 9444 7528
rect 9364 7488 9370 7500
rect 4856 7432 5212 7460
rect 5460 7432 5580 7460
rect 5736 7432 6592 7460
rect 4856 7420 4862 7432
rect 1268 7364 2176 7392
rect 2593 7395 2651 7401
rect 1268 7352 1274 7364
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3697 7395 3755 7401
rect 2639 7364 3648 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 842 7284 848 7336
rect 900 7284 906 7336
rect 2222 7284 2228 7336
rect 2280 7284 2286 7336
rect 2866 7284 2872 7336
rect 2924 7284 2930 7336
rect 3620 7324 3648 7364
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3786 7352 3792 7404
rect 3844 7352 3850 7404
rect 4816 7364 5107 7392
rect 4816 7336 4844 7364
rect 4154 7324 4160 7336
rect 3620 7296 4160 7324
rect 4154 7284 4160 7296
rect 4212 7324 4218 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4212 7296 4629 7324
rect 4212 7284 4218 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7320 5043 7327
rect 5079 7320 5107 7364
rect 5184 7333 5212 7432
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 5552 7392 5580 7432
rect 5552 7364 6500 7392
rect 5031 7293 5107 7320
rect 4985 7292 5107 7293
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7293 5227 7327
rect 5460 7324 5488 7352
rect 5552 7333 5580 7364
rect 4985 7287 5043 7292
rect 5169 7287 5227 7293
rect 5368 7296 5488 7324
rect 5537 7327 5595 7333
rect 1121 7259 1179 7265
rect 1121 7225 1133 7259
rect 1167 7225 1179 7259
rect 1121 7219 1179 7225
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 1136 7188 1164 7219
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 2832 7228 4108 7256
rect 2832 7216 2838 7228
rect 992 7160 1164 7188
rect 992 7148 998 7160
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 2648 7160 3617 7188
rect 2648 7148 2654 7160
rect 3605 7157 3617 7160
rect 3651 7188 3663 7191
rect 3878 7188 3884 7200
rect 3651 7160 3884 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4080 7197 4108 7228
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4890 7256 4896 7268
rect 4580 7228 4896 7256
rect 4580 7216 4586 7228
rect 4890 7216 4896 7228
rect 4948 7256 4954 7268
rect 5368 7265 5396 7296
rect 5537 7293 5549 7327
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 5353 7259 5411 7265
rect 4948 7228 5304 7256
rect 4948 7216 4954 7228
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4764 7160 4813 7188
rect 4764 7148 4770 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 5276 7188 5304 7228
rect 5353 7225 5365 7259
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 5441 7259 5499 7265
rect 5441 7225 5453 7259
rect 5487 7256 5499 7259
rect 5626 7256 5632 7268
rect 5487 7228 5632 7256
rect 5487 7225 5499 7228
rect 5441 7219 5499 7225
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7225 6055 7259
rect 6472 7256 6500 7364
rect 6564 7320 6592 7432
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 6696 7432 6868 7460
rect 6696 7420 6702 7432
rect 6840 7333 6868 7432
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 7892 7432 8161 7460
rect 7892 7420 7898 7432
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7282 7352 7288 7404
rect 7340 7392 7346 7404
rect 8133 7392 8161 7432
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8260 7432 8493 7460
rect 8260 7420 8266 7432
rect 8481 7429 8493 7432
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 8904 7432 9357 7460
rect 8904 7420 8910 7432
rect 9214 7392 9220 7404
rect 7340 7364 7972 7392
rect 8133 7364 8248 7392
rect 7340 7352 7346 7364
rect 7944 7336 7972 7364
rect 6733 7327 6791 7333
rect 6733 7324 6745 7327
rect 6656 7320 6745 7324
rect 6564 7296 6745 7320
rect 6564 7292 6684 7296
rect 6733 7293 6745 7296
rect 6779 7293 6791 7327
rect 6733 7287 6791 7293
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 7558 7324 7564 7336
rect 6825 7287 6883 7293
rect 7024 7296 7564 7324
rect 7024 7256 7052 7296
rect 7558 7284 7564 7296
rect 7616 7324 7622 7336
rect 7699 7327 7757 7333
rect 7699 7324 7711 7327
rect 7616 7296 7711 7324
rect 7616 7284 7622 7296
rect 7699 7293 7711 7296
rect 7745 7293 7757 7327
rect 7699 7287 7757 7293
rect 7926 7284 7932 7336
rect 7984 7284 7990 7336
rect 8018 7284 8024 7336
rect 8076 7333 8082 7336
rect 8220 7333 8248 7364
rect 8312 7364 8616 7392
rect 8312 7336 8340 7364
rect 8076 7327 8115 7333
rect 8103 7293 8115 7327
rect 8076 7287 8115 7293
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8076 7284 8082 7287
rect 8294 7284 8300 7336
rect 8352 7284 8358 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8404 7296 8493 7324
rect 7285 7259 7343 7265
rect 7285 7256 7297 7259
rect 6472 7228 7052 7256
rect 7116 7228 7297 7256
rect 5997 7219 6055 7225
rect 6012 7188 6040 7219
rect 5276 7160 6040 7188
rect 4801 7151 4859 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 7116 7188 7144 7228
rect 7285 7225 7297 7228
rect 7331 7225 7343 7259
rect 7285 7219 7343 7225
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7524 7228 7849 7256
rect 7524 7216 7530 7228
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 6604 7160 7144 7188
rect 6604 7148 6610 7160
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 7248 7160 7389 7188
rect 7248 7148 7254 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8404 7188 8432 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8588 7256 8616 7364
rect 8864 7364 9220 7392
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 8864 7333 8892 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9030 7333 9036 7336
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 8997 7327 9036 7333
rect 8997 7293 9009 7327
rect 8997 7287 9036 7293
rect 9030 7284 9036 7287
rect 9088 7284 9094 7336
rect 9329 7333 9357 7432
rect 9416 7392 9444 7500
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10226 7528 10232 7540
rect 9723 7500 10232 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10413 7531 10471 7537
rect 10413 7497 10425 7531
rect 10459 7528 10471 7531
rect 10962 7528 10968 7540
rect 10459 7500 10968 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11146 7488 11152 7540
rect 11204 7488 11210 7540
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 11606 7528 11612 7540
rect 11563 7500 11612 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11606 7488 11612 7500
rect 11664 7528 11670 7540
rect 11664 7500 15884 7528
rect 11664 7488 11670 7500
rect 9493 7463 9551 7469
rect 9493 7429 9505 7463
rect 9539 7460 9551 7463
rect 9766 7460 9772 7472
rect 9539 7432 9772 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 11164 7460 11192 7488
rect 11698 7460 11704 7472
rect 11164 7432 11704 7460
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 13354 7460 13360 7472
rect 13188 7432 13360 7460
rect 10134 7392 10140 7404
rect 9416 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10192 7364 10885 7392
rect 10192 7352 10198 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 11422 7392 11428 7404
rect 10873 7355 10931 7361
rect 11072 7364 11428 7392
rect 9314 7327 9372 7333
rect 9314 7293 9326 7327
rect 9360 7293 9372 7327
rect 9314 7287 9372 7293
rect 9858 7284 9864 7336
rect 9916 7284 9922 7336
rect 9950 7284 9956 7336
rect 10008 7284 10014 7336
rect 10042 7284 10048 7336
rect 10100 7284 10106 7336
rect 10226 7284 10232 7336
rect 10284 7284 10290 7336
rect 10594 7284 10600 7336
rect 10652 7284 10658 7336
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 10962 7284 10968 7336
rect 11020 7284 11026 7336
rect 11072 7333 11100 7364
rect 11422 7352 11428 7364
rect 11480 7392 11486 7404
rect 11480 7364 11547 7392
rect 11480 7352 11486 7364
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8588 7228 9137 7256
rect 8588 7200 8616 7228
rect 9125 7225 9137 7228
rect 9171 7225 9183 7259
rect 9125 7219 9183 7225
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 10060 7256 10088 7284
rect 10870 7256 10876 7268
rect 9263 7228 9996 7256
rect 10060 7228 10876 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9968 7200 9996 7228
rect 10870 7216 10876 7228
rect 10928 7256 10934 7268
rect 11164 7256 11192 7287
rect 10928 7228 11192 7256
rect 10928 7216 10934 7228
rect 7708 7160 8432 7188
rect 7708 7148 7714 7160
rect 8570 7148 8576 7200
rect 8628 7148 8634 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9306 7188 9312 7200
rect 9088 7160 9312 7188
rect 9088 7148 9094 7160
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11146 7188 11152 7200
rect 11020 7160 11152 7188
rect 11020 7148 11026 7160
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 11422 7148 11428 7200
rect 11480 7148 11486 7200
rect 11519 7188 11547 7364
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 13188 7392 13216 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13541 7463 13599 7469
rect 13541 7429 13553 7463
rect 13587 7460 13599 7463
rect 13587 7432 13676 7460
rect 13587 7429 13599 7432
rect 13541 7423 13599 7429
rect 12492 7364 13216 7392
rect 13265 7395 13323 7401
rect 12492 7352 12498 7364
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13446 7392 13452 7404
rect 13311 7364 13452 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13648 7324 13676 7432
rect 15562 7420 15568 7472
rect 15620 7420 15626 7472
rect 15749 7463 15807 7469
rect 15749 7429 15761 7463
rect 15795 7429 15807 7463
rect 15749 7423 15807 7429
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 15764 7392 15792 7423
rect 14516 7364 15792 7392
rect 14516 7352 14522 7364
rect 13280 7296 13676 7324
rect 13725 7327 13783 7333
rect 12894 7256 12900 7268
rect 12558 7228 12900 7256
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7256 13047 7259
rect 13280 7256 13308 7296
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13035 7228 13308 7256
rect 13035 7225 13047 7228
rect 12989 7219 13047 7225
rect 13354 7216 13360 7268
rect 13412 7256 13418 7268
rect 13740 7256 13768 7287
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 13412 7228 13768 7256
rect 13412 7216 13418 7228
rect 14090 7216 14096 7268
rect 14148 7216 14154 7268
rect 15102 7188 15108 7200
rect 11519 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15856 7188 15884 7500
rect 18046 7488 18052 7540
rect 18104 7488 18110 7540
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 20441 7531 20499 7537
rect 20441 7528 20453 7531
rect 19668 7500 20453 7528
rect 19668 7488 19674 7500
rect 20441 7497 20453 7500
rect 20487 7528 20499 7531
rect 23198 7528 23204 7540
rect 20487 7500 23204 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 23658 7488 23664 7540
rect 23716 7488 23722 7540
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 24394 7528 24400 7540
rect 23808 7500 24400 7528
rect 23808 7488 23814 7500
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 26053 7531 26111 7537
rect 25149 7500 26004 7528
rect 16482 7460 16488 7472
rect 16132 7432 16488 7460
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 16132 7401 16160 7432
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7460 17279 7463
rect 18064 7460 18092 7488
rect 17267 7432 18092 7460
rect 17267 7429 17279 7432
rect 17221 7423 17279 7429
rect 20806 7420 20812 7472
rect 20864 7420 20870 7472
rect 23014 7460 23020 7472
rect 21652 7432 23020 7460
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 15988 7364 16129 7392
rect 15988 7352 15994 7364
rect 16117 7361 16129 7364
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16298 7352 16304 7404
rect 16356 7352 16362 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 16850 7392 16856 7404
rect 16715 7364 16856 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 17920 7364 18245 7392
rect 17920 7352 17926 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 18690 7352 18696 7404
rect 18748 7352 18754 7404
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 19024 7364 20760 7392
rect 19024 7352 19030 7364
rect 17678 7324 17684 7336
rect 16224 7296 17684 7324
rect 16224 7265 16252 7296
rect 17678 7284 17684 7296
rect 17736 7324 17742 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 17736 7296 17785 7324
rect 17736 7284 17742 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 18138 7284 18144 7336
rect 18196 7284 18202 7336
rect 18322 7284 18328 7336
rect 18380 7284 18386 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 20070 7284 20076 7336
rect 20128 7284 20134 7336
rect 16209 7259 16267 7265
rect 16209 7225 16221 7259
rect 16255 7225 16267 7259
rect 17957 7259 18015 7265
rect 16209 7219 16267 7225
rect 16316 7228 17724 7256
rect 16316 7188 16344 7228
rect 15856 7160 16344 7188
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 16942 7188 16948 7200
rect 16899 7160 16948 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 16942 7148 16948 7160
rect 17000 7188 17006 7200
rect 17589 7191 17647 7197
rect 17589 7188 17601 7191
rect 17000 7160 17601 7188
rect 17000 7148 17006 7160
rect 17589 7157 17601 7160
rect 17635 7157 17647 7191
rect 17696 7188 17724 7228
rect 17957 7225 17969 7259
rect 18003 7256 18015 7259
rect 18969 7259 19027 7265
rect 18969 7256 18981 7259
rect 18003 7228 18981 7256
rect 18003 7225 18015 7228
rect 17957 7219 18015 7225
rect 18969 7225 18981 7228
rect 19015 7225 19027 7259
rect 20732 7256 20760 7364
rect 20824 7324 20852 7420
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7392 21235 7395
rect 21542 7392 21548 7404
rect 21223 7364 21548 7392
rect 21223 7361 21235 7364
rect 21177 7355 21235 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20824 7296 21097 7324
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 21453 7327 21511 7333
rect 21453 7324 21465 7327
rect 21324 7296 21465 7324
rect 21324 7284 21330 7296
rect 21453 7293 21465 7296
rect 21499 7324 21511 7327
rect 21652 7324 21680 7432
rect 23014 7420 23020 7432
rect 23072 7420 23078 7472
rect 23109 7463 23167 7469
rect 23109 7429 23121 7463
rect 23155 7429 23167 7463
rect 23676 7460 23704 7488
rect 23676 7432 24164 7460
rect 23109 7423 23167 7429
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22066 7364 22661 7392
rect 21499 7296 21680 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 21910 7284 21916 7336
rect 21968 7284 21974 7336
rect 21634 7256 21640 7268
rect 20732 7228 21640 7256
rect 18969 7219 19027 7225
rect 21634 7216 21640 7228
rect 21692 7216 21698 7268
rect 22066 7188 22094 7364
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 23124 7392 23152 7423
rect 23124 7364 23704 7392
rect 22189 7327 22247 7333
rect 22189 7293 22201 7327
rect 22235 7324 22247 7327
rect 22278 7324 22284 7336
rect 22235 7296 22284 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 17696 7160 22094 7188
rect 17589 7151 17647 7157
rect 22278 7148 22284 7200
rect 22336 7148 22342 7200
rect 22388 7188 22416 7287
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22520 7296 22569 7324
rect 22520 7284 22526 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 22646 7216 22652 7268
rect 22704 7216 22710 7268
rect 22554 7188 22560 7200
rect 22388 7160 22560 7188
rect 22554 7148 22560 7160
rect 22612 7188 22618 7200
rect 23124 7188 23152 7364
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 23676 7333 23704 7364
rect 23860 7364 24072 7392
rect 23860 7336 23888 7364
rect 23477 7327 23535 7333
rect 23477 7324 23489 7327
rect 23256 7296 23489 7324
rect 23256 7284 23262 7296
rect 23477 7293 23489 7296
rect 23523 7293 23535 7327
rect 23477 7287 23535 7293
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 23750 7324 23756 7336
rect 23707 7296 23756 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 23842 7284 23848 7336
rect 23900 7284 23906 7336
rect 24044 7333 24072 7364
rect 24136 7333 24164 7432
rect 24210 7420 24216 7472
rect 24268 7420 24274 7472
rect 24228 7392 24256 7420
rect 25149 7392 25177 7500
rect 25225 7463 25283 7469
rect 25225 7429 25237 7463
rect 25271 7460 25283 7463
rect 25774 7460 25780 7472
rect 25271 7432 25780 7460
rect 25271 7429 25283 7432
rect 25225 7423 25283 7429
rect 25774 7420 25780 7432
rect 25832 7420 25838 7472
rect 25976 7460 26004 7500
rect 26053 7497 26065 7531
rect 26099 7528 26111 7531
rect 28994 7528 29000 7540
rect 26099 7500 29000 7528
rect 26099 7497 26111 7500
rect 26053 7491 26111 7497
rect 28994 7488 29000 7500
rect 29052 7488 29058 7540
rect 26326 7460 26332 7472
rect 25976 7432 26332 7460
rect 26326 7420 26332 7432
rect 26384 7420 26390 7472
rect 28258 7420 28264 7472
rect 28316 7420 28322 7472
rect 24228 7364 25177 7392
rect 23937 7327 23995 7333
rect 23937 7293 23949 7327
rect 23983 7293 23995 7327
rect 23937 7287 23995 7293
rect 24029 7327 24087 7333
rect 24029 7293 24041 7327
rect 24075 7293 24087 7327
rect 24136 7327 24198 7333
rect 24136 7296 24152 7327
rect 24029 7287 24087 7293
rect 24140 7293 24152 7296
rect 24186 7293 24198 7327
rect 24228 7324 24256 7364
rect 24305 7327 24363 7333
rect 24305 7324 24317 7327
rect 24228 7296 24317 7324
rect 24140 7287 24198 7293
rect 24305 7293 24317 7296
rect 24351 7293 24363 7327
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24305 7287 24363 7293
rect 24412 7296 24593 7324
rect 23952 7256 23980 7287
rect 24412 7256 24440 7296
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 24581 7287 24639 7293
rect 24670 7284 24676 7336
rect 24728 7324 24734 7336
rect 24872 7333 24900 7364
rect 25498 7352 25504 7404
rect 25556 7352 25562 7404
rect 26510 7352 26516 7404
rect 26568 7392 26574 7404
rect 26786 7392 26792 7404
rect 26568 7364 26792 7392
rect 26568 7352 26574 7364
rect 26786 7352 26792 7364
rect 26844 7352 26850 7404
rect 24765 7327 24823 7333
rect 24765 7324 24777 7327
rect 24728 7296 24777 7324
rect 24728 7284 24734 7296
rect 24765 7293 24777 7296
rect 24811 7293 24823 7327
rect 24765 7287 24823 7293
rect 24857 7327 24915 7333
rect 24857 7293 24869 7327
rect 24903 7293 24915 7327
rect 24857 7287 24915 7293
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 26234 7324 26240 7336
rect 25521 7296 26240 7324
rect 23492 7228 24440 7256
rect 23492 7200 23520 7228
rect 22612 7160 23152 7188
rect 22612 7148 22618 7160
rect 23474 7148 23480 7200
rect 23532 7148 23538 7200
rect 23569 7191 23627 7197
rect 23569 7157 23581 7191
rect 23615 7188 23627 7191
rect 24118 7188 24124 7200
rect 23615 7160 24124 7188
rect 23615 7157 23627 7160
rect 23569 7151 23627 7157
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24412 7188 24440 7228
rect 24489 7259 24547 7265
rect 24489 7225 24501 7259
rect 24535 7256 24547 7259
rect 25314 7256 25320 7268
rect 24535 7228 25320 7256
rect 24535 7225 24547 7228
rect 24489 7219 24547 7225
rect 25314 7216 25320 7228
rect 25372 7216 25378 7268
rect 25222 7188 25228 7200
rect 24412 7160 25228 7188
rect 25222 7148 25228 7160
rect 25280 7188 25286 7200
rect 25521 7188 25549 7296
rect 26234 7284 26240 7296
rect 26292 7324 26298 7336
rect 26329 7327 26387 7333
rect 26329 7324 26341 7327
rect 26292 7296 26341 7324
rect 26292 7284 26298 7296
rect 26329 7293 26341 7296
rect 26375 7293 26387 7327
rect 26329 7287 26387 7293
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 28276 7324 28304 7420
rect 26467 7296 26740 7324
rect 28198 7296 28304 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 26712 7268 26740 7296
rect 26605 7259 26663 7265
rect 26605 7256 26617 7259
rect 26160 7228 26617 7256
rect 26160 7200 26188 7228
rect 26605 7225 26617 7228
rect 26651 7225 26663 7259
rect 26605 7219 26663 7225
rect 26694 7216 26700 7268
rect 26752 7216 26758 7268
rect 27065 7259 27123 7265
rect 27065 7225 27077 7259
rect 27111 7225 27123 7259
rect 27065 7219 27123 7225
rect 25280 7160 25549 7188
rect 25280 7148 25286 7160
rect 25590 7148 25596 7200
rect 25648 7148 25654 7200
rect 25682 7148 25688 7200
rect 25740 7148 25746 7200
rect 26142 7148 26148 7200
rect 26200 7148 26206 7200
rect 26513 7191 26571 7197
rect 26513 7157 26525 7191
rect 26559 7188 26571 7191
rect 26878 7188 26884 7200
rect 26559 7160 26884 7188
rect 26559 7157 26571 7160
rect 26513 7151 26571 7157
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 27080 7188 27108 7219
rect 28810 7216 28816 7268
rect 28868 7216 28874 7268
rect 27982 7188 27988 7200
rect 27080 7160 27988 7188
rect 27982 7148 27988 7160
rect 28040 7148 28046 7200
rect 552 7098 31808 7120
rect 552 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 15946 7098
rect 15998 7046 16010 7098
rect 16062 7046 16074 7098
rect 16126 7046 16138 7098
rect 16190 7046 16202 7098
rect 16254 7046 23720 7098
rect 23772 7046 23784 7098
rect 23836 7046 23848 7098
rect 23900 7046 23912 7098
rect 23964 7046 23976 7098
rect 24028 7046 31494 7098
rect 31546 7046 31558 7098
rect 31610 7046 31622 7098
rect 31674 7046 31686 7098
rect 31738 7046 31750 7098
rect 31802 7046 31808 7098
rect 552 7024 31808 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 3418 6984 3424 6996
rect 1728 6956 3424 6984
rect 1728 6944 1734 6956
rect 3418 6944 3424 6956
rect 3476 6984 3482 6996
rect 3476 6956 3556 6984
rect 3476 6944 3482 6956
rect 1688 6916 1716 6944
rect 1228 6888 1716 6916
rect 2041 6919 2099 6925
rect 1026 6808 1032 6860
rect 1084 6808 1090 6860
rect 1228 6857 1256 6888
rect 2041 6885 2053 6919
rect 2087 6916 2099 6919
rect 2498 6916 2504 6928
rect 2087 6888 2504 6916
rect 2087 6885 2099 6888
rect 2041 6879 2099 6885
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 3528 6872 3556 6956
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4617 6987 4675 6993
rect 4028 6956 4568 6984
rect 4028 6944 4034 6956
rect 4540 6916 4568 6956
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 5258 6984 5264 6996
rect 4663 6956 5264 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6546 6984 6552 6996
rect 5592 6956 6552 6984
rect 5592 6944 5598 6956
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7466 6984 7472 6996
rect 7340 6956 7472 6984
rect 7340 6944 7346 6956
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 10042 6984 10048 6996
rect 7616 6956 10048 6984
rect 7616 6944 7622 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10410 6944 10416 6996
rect 10468 6944 10474 6996
rect 11238 6944 11244 6996
rect 11296 6944 11302 6996
rect 11422 6944 11428 6996
rect 11480 6944 11486 6996
rect 11606 6944 11612 6996
rect 11664 6944 11670 6996
rect 11701 6987 11759 6993
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 11790 6984 11796 6996
rect 11747 6956 11796 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 11790 6944 11796 6956
rect 11848 6984 11854 6996
rect 11974 6984 11980 6996
rect 11848 6956 11980 6984
rect 11848 6944 11854 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12434 6984 12440 6996
rect 12115 6956 12440 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 13446 6984 13452 6996
rect 12544 6956 13452 6984
rect 4540 6888 5396 6916
rect 1213 6851 1271 6857
rect 1213 6817 1225 6851
rect 1259 6817 1271 6851
rect 1213 6811 1271 6817
rect 1305 6851 1363 6857
rect 1305 6817 1317 6851
rect 1351 6848 1363 6851
rect 1394 6848 1400 6860
rect 1351 6820 1400 6848
rect 1351 6817 1363 6820
rect 1305 6811 1363 6817
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1486 6808 1492 6860
rect 1544 6808 1550 6860
rect 1578 6808 1584 6860
rect 1636 6808 1642 6860
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 2774 6848 2780 6860
rect 2179 6820 2780 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 2866 6808 2872 6860
rect 2924 6808 2930 6860
rect 3418 6808 3424 6860
rect 3476 6808 3482 6860
rect 3528 6857 3648 6872
rect 3528 6851 3663 6857
rect 3528 6844 3617 6851
rect 3605 6817 3617 6844
rect 3651 6817 3663 6851
rect 3605 6811 3663 6817
rect 3697 6851 3755 6857
rect 3697 6817 3709 6851
rect 3743 6817 3755 6851
rect 3697 6811 3755 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6817 3847 6851
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3789 6811 3847 6817
rect 3896 6820 4077 6848
rect 1504 6780 1532 6808
rect 1504 6752 2268 6780
rect 1670 6672 1676 6724
rect 1728 6672 1734 6724
rect 2240 6712 2268 6752
rect 2314 6740 2320 6792
rect 2372 6740 2378 6792
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3712 6780 3740 6811
rect 3200 6752 3740 6780
rect 3200 6740 3206 6752
rect 2240 6684 3556 6712
rect 1026 6604 1032 6656
rect 1084 6644 1090 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 1084 6616 2513 6644
rect 1084 6604 1090 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 3528 6644 3556 6684
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 3804 6712 3832 6811
rect 3660 6684 3832 6712
rect 3660 6672 3666 6684
rect 3896 6644 3924 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4709 6851 4767 6857
rect 4479 6820 4568 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4172 6780 4200 6811
rect 3988 6752 4200 6780
rect 3988 6721 4016 6752
rect 3973 6715 4031 6721
rect 3973 6681 3985 6715
rect 4019 6681 4031 6715
rect 4356 6712 4384 6811
rect 4540 6792 4568 6820
rect 4709 6817 4721 6851
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4724 6780 4752 6811
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 5040 6820 5089 6848
rect 5040 6808 5046 6820
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 5368 6857 5396 6888
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 8021 6919 8079 6925
rect 5868 6888 6316 6916
rect 5868 6876 5874 6888
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6817 6239 6851
rect 6288 6848 6316 6888
rect 8021 6885 8033 6919
rect 8067 6916 8079 6919
rect 8110 6916 8116 6928
rect 8067 6888 8116 6916
rect 8067 6885 8079 6888
rect 8021 6879 8079 6885
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 10428 6916 10456 6944
rect 11256 6916 11284 6944
rect 9646 6888 10456 6916
rect 10888 6888 11284 6916
rect 11440 6916 11468 6944
rect 11440 6888 12204 6916
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 6288 6820 6868 6848
rect 6181 6811 6239 6817
rect 5534 6780 5540 6792
rect 4724 6752 5540 6780
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5810 6780 5816 6792
rect 5675 6752 5816 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 4798 6712 4804 6724
rect 4356 6684 4804 6712
rect 3973 6675 4031 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 4893 6715 4951 6721
rect 4893 6681 4905 6715
rect 4939 6712 4951 6715
rect 5442 6712 5448 6724
rect 4939 6684 5448 6712
rect 4939 6681 4951 6684
rect 4893 6675 4951 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5718 6672 5724 6724
rect 5776 6672 5782 6724
rect 6196 6712 6224 6811
rect 6840 6792 6868 6820
rect 7024 6820 7757 6848
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7024 6780 7052 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 9646 6848 9674 6888
rect 9232 6820 9674 6848
rect 6972 6752 7052 6780
rect 7101 6783 7159 6789
rect 6972 6740 6978 6752
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7558 6780 7564 6792
rect 7147 6752 7564 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 8754 6780 8760 6792
rect 7852 6752 8760 6780
rect 7852 6712 7880 6752
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9232 6780 9260 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9824 6820 9965 6848
rect 9824 6808 9830 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 10597 6851 10655 6857
rect 10244 6820 10456 6848
rect 9088 6752 9260 6780
rect 9493 6783 9551 6789
rect 9088 6740 9094 6752
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 9674 6780 9680 6792
rect 9539 6752 9680 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10244 6712 10272 6820
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10428 6780 10456 6820
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10888 6848 10916 6888
rect 10643 6820 10916 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 12176 6857 12204 6888
rect 12544 6860 12572 6956
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 13688 6956 14749 6984
rect 13688 6944 13694 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 14737 6947 14795 6953
rect 14844 6956 16497 6984
rect 14182 6876 14188 6928
rect 14240 6916 14246 6928
rect 14844 6916 14872 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 19426 6984 19432 6996
rect 16485 6947 16543 6953
rect 16592 6956 19432 6984
rect 14240 6888 14872 6916
rect 14240 6876 14246 6888
rect 15102 6876 15108 6928
rect 15160 6916 15166 6928
rect 15381 6919 15439 6925
rect 15381 6916 15393 6919
rect 15160 6888 15393 6916
rect 15160 6876 15166 6888
rect 15381 6885 15393 6888
rect 15427 6916 15439 6919
rect 16592 6916 16620 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 20809 6987 20867 6993
rect 20809 6984 20821 6987
rect 20312 6956 20821 6984
rect 20312 6944 20318 6956
rect 20809 6953 20821 6956
rect 20855 6953 20867 6987
rect 25590 6984 25596 6996
rect 20809 6947 20867 6953
rect 22296 6956 25596 6984
rect 17494 6916 17500 6928
rect 15427 6888 16620 6916
rect 17236 6888 17500 6916
rect 15427 6885 15439 6888
rect 15381 6879 15439 6885
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6848 11207 6851
rect 12161 6851 12219 6857
rect 11195 6820 11652 6848
rect 11195 6817 11207 6820
rect 11149 6811 11207 6817
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10428 6752 11069 6780
rect 10321 6743 10379 6749
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 6196 6684 7880 6712
rect 9508 6684 10272 6712
rect 4062 6644 4068 6656
rect 3528 6616 4068 6644
rect 2501 6607 2559 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5258 6644 5264 6656
rect 5132 6616 5264 6644
rect 5132 6604 5138 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 5736 6644 5764 6672
rect 9508 6656 9536 6684
rect 5583 6616 5764 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6086 6604 6092 6656
rect 6144 6604 6150 6656
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 7742 6644 7748 6656
rect 7699 6616 7748 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 10192 6616 10241 6644
rect 10192 6604 10198 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10336 6644 10364 6743
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11624 6780 11652 6820
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 11698 6780 11704 6792
rect 11624 6752 11704 6780
rect 11517 6743 11575 6749
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 11348 6712 11376 6740
rect 10827 6684 11376 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 11532 6656 11560 6743
rect 11698 6740 11704 6752
rect 11756 6780 11762 6792
rect 12434 6780 12440 6792
rect 11756 6752 12440 6780
rect 11756 6740 11762 6752
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13924 6780 13952 6834
rect 14844 6820 15301 6848
rect 14461 6783 14519 6789
rect 12952 6752 14412 6780
rect 12952 6740 12958 6752
rect 11422 6644 11428 6656
rect 10336 6616 11428 6644
rect 10229 6607 10287 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 11572 6616 12357 6644
rect 11572 6604 11578 6616
rect 12345 6613 12357 6616
rect 12391 6644 12403 6647
rect 12618 6644 12624 6656
rect 12391 6616 12624 6644
rect 12391 6613 12403 6616
rect 12345 6607 12403 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 13446 6604 13452 6656
rect 13504 6644 13510 6656
rect 14182 6644 14188 6656
rect 13504 6616 14188 6644
rect 13504 6604 13510 6616
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 14274 6604 14280 6656
rect 14332 6604 14338 6656
rect 14384 6644 14412 6752
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14476 6712 14504 6743
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14608 6752 14657 6780
rect 14608 6740 14614 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14844 6712 14872 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 17236 6848 17264 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 18322 6876 18328 6928
rect 18380 6916 18386 6928
rect 18417 6919 18475 6925
rect 18417 6916 18429 6919
rect 18380 6888 18429 6916
rect 18380 6876 18386 6888
rect 18417 6885 18429 6888
rect 18463 6885 18475 6919
rect 21910 6916 21916 6928
rect 18417 6879 18475 6885
rect 20548 6888 21916 6916
rect 20548 6860 20576 6888
rect 21910 6876 21916 6888
rect 21968 6916 21974 6928
rect 21968 6888 22232 6916
rect 21968 6876 21974 6888
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 15335 6820 17264 6848
rect 17328 6820 17417 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 16224 6789 16252 6820
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 14976 6752 15393 6780
rect 14976 6740 14982 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6780 16451 6783
rect 16482 6780 16488 6792
rect 16439 6752 16488 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 15010 6712 15016 6724
rect 14476 6684 15016 6712
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15105 6715 15163 6721
rect 15105 6681 15117 6715
rect 15151 6712 15163 6715
rect 17328 6712 17356 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 17604 6780 17632 6811
rect 17678 6808 17684 6860
rect 17736 6848 17742 6860
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17736 6820 17969 6848
rect 17736 6808 17742 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 18785 6851 18843 6857
rect 18785 6817 18797 6851
rect 18831 6848 18843 6851
rect 18831 6820 19334 6848
rect 18831 6817 18843 6820
rect 18785 6811 18843 6817
rect 18138 6780 18144 6792
rect 17604 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6780 18383 6783
rect 18414 6780 18420 6792
rect 18371 6752 18420 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6749 19119 6783
rect 19306 6780 19334 6820
rect 19794 6808 19800 6860
rect 19852 6848 19858 6860
rect 19889 6851 19947 6857
rect 19889 6848 19901 6851
rect 19852 6820 19901 6848
rect 19852 6808 19858 6820
rect 19889 6817 19901 6820
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 20162 6848 20168 6860
rect 20119 6820 20168 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 20254 6808 20260 6860
rect 20312 6848 20318 6860
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 20312 6820 20361 6848
rect 20312 6808 20318 6820
rect 20349 6817 20361 6820
rect 20395 6817 20407 6851
rect 20349 6811 20407 6817
rect 20530 6808 20536 6860
rect 20588 6808 20594 6860
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19306 6752 19717 6780
rect 19061 6743 19119 6749
rect 19705 6749 19717 6752
rect 19751 6780 19763 6783
rect 21468 6780 21496 6811
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 22204 6857 22232 6888
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 21692 6820 21833 6848
rect 21692 6808 21698 6820
rect 21821 6817 21833 6820
rect 21867 6817 21879 6851
rect 21821 6811 21879 6817
rect 22189 6851 22247 6857
rect 22189 6817 22201 6851
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 19751 6752 21496 6780
rect 21836 6780 21864 6811
rect 22296 6780 22324 6956
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 25869 6987 25927 6993
rect 25869 6953 25881 6987
rect 25915 6984 25927 6987
rect 26326 6984 26332 6996
rect 25915 6956 26332 6984
rect 25915 6953 25927 6956
rect 25869 6947 25927 6953
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 22557 6919 22615 6925
rect 22557 6916 22569 6919
rect 22520 6888 22569 6916
rect 22520 6876 22526 6888
rect 22557 6885 22569 6888
rect 22603 6885 22615 6919
rect 22557 6879 22615 6885
rect 22649 6919 22707 6925
rect 22649 6885 22661 6919
rect 22695 6885 22707 6919
rect 22649 6879 22707 6885
rect 22664 6848 22692 6879
rect 22922 6876 22928 6928
rect 22980 6916 22986 6928
rect 23290 6916 23296 6928
rect 22980 6888 23296 6916
rect 22980 6876 22986 6888
rect 23290 6876 23296 6888
rect 23348 6916 23354 6928
rect 24946 6916 24952 6928
rect 23348 6888 24952 6916
rect 23348 6876 23354 6888
rect 24946 6876 24952 6888
rect 25004 6916 25010 6928
rect 25004 6888 25084 6916
rect 25004 6876 25010 6888
rect 21836 6752 22324 6780
rect 22388 6820 22692 6848
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 17954 6712 17960 6724
rect 15151 6684 17960 6712
rect 15151 6681 15163 6684
rect 15105 6675 15163 6681
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 18248 6712 18276 6740
rect 18874 6712 18880 6724
rect 18248 6684 18880 6712
rect 18874 6672 18880 6684
rect 18932 6672 18938 6724
rect 18966 6672 18972 6724
rect 19024 6672 19030 6724
rect 19076 6712 19104 6743
rect 20438 6712 20444 6724
rect 19076 6684 20444 6712
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 20533 6715 20591 6721
rect 20533 6681 20545 6715
rect 20579 6712 20591 6715
rect 21174 6712 21180 6724
rect 20579 6684 21180 6712
rect 20579 6681 20591 6684
rect 20533 6675 20591 6681
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 21453 6715 21511 6721
rect 21453 6681 21465 6715
rect 21499 6681 21511 6715
rect 21453 6675 21511 6681
rect 15194 6644 15200 6656
rect 14384 6616 15200 6644
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15838 6604 15844 6656
rect 15896 6604 15902 6656
rect 16850 6604 16856 6656
rect 16908 6604 16914 6656
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 18598 6604 18604 6656
rect 18656 6604 18662 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19794 6644 19800 6656
rect 19392 6616 19800 6644
rect 19392 6604 19398 6616
rect 19794 6604 19800 6616
rect 19852 6604 19858 6656
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 21468 6644 21496 6675
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 22388 6712 22416 6820
rect 23566 6808 23572 6860
rect 23624 6808 23630 6860
rect 24118 6808 24124 6860
rect 24176 6808 24182 6860
rect 24210 6808 24216 6860
rect 24268 6808 24274 6860
rect 24302 6808 24308 6860
rect 24360 6848 24366 6860
rect 24486 6848 24492 6860
rect 24360 6820 24492 6848
rect 24360 6808 24366 6820
rect 24486 6808 24492 6820
rect 24544 6848 24550 6860
rect 25056 6857 25084 6888
rect 25406 6876 25412 6928
rect 25464 6916 25470 6928
rect 25884 6916 25912 6947
rect 26326 6944 26332 6956
rect 26384 6944 26390 6996
rect 26634 6993 26640 6996
rect 26605 6987 26640 6993
rect 26605 6953 26617 6987
rect 26605 6947 26640 6953
rect 26634 6944 26640 6947
rect 26692 6944 26698 6996
rect 28074 6944 28080 6996
rect 28132 6984 28138 6996
rect 28721 6987 28779 6993
rect 28721 6984 28733 6987
rect 28132 6956 28733 6984
rect 28132 6944 28138 6956
rect 28721 6953 28733 6956
rect 28767 6953 28779 6987
rect 28721 6947 28779 6953
rect 28994 6944 29000 6996
rect 29052 6944 29058 6996
rect 25464 6888 25912 6916
rect 26160 6888 26740 6916
rect 25464 6876 25470 6888
rect 26160 6860 26188 6888
rect 24673 6851 24731 6857
rect 24673 6848 24685 6851
rect 24544 6820 24685 6848
rect 24544 6808 24550 6820
rect 24673 6817 24685 6820
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 25041 6851 25099 6857
rect 25041 6817 25053 6851
rect 25087 6817 25099 6851
rect 26142 6848 26148 6860
rect 25041 6811 25099 6817
rect 25148 6820 26148 6848
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 22244 6684 22416 6712
rect 23109 6715 23167 6721
rect 22244 6672 22250 6684
rect 23109 6681 23121 6715
rect 23155 6712 23167 6715
rect 23474 6712 23480 6724
rect 23155 6684 23480 6712
rect 23155 6681 23167 6684
rect 23109 6675 23167 6681
rect 23474 6672 23480 6684
rect 23532 6672 23538 6724
rect 24136 6712 24164 6808
rect 25148 6792 25176 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26234 6808 26240 6860
rect 26292 6848 26298 6860
rect 26712 6857 26740 6888
rect 28534 6876 28540 6928
rect 28592 6876 28598 6928
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 26292 6820 26433 6848
rect 26292 6808 26298 6820
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 26697 6851 26755 6857
rect 26697 6817 26709 6851
rect 26743 6817 26755 6851
rect 26697 6811 26755 6817
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 26881 6851 26939 6857
rect 26881 6848 26893 6851
rect 26844 6820 26893 6848
rect 26844 6808 26850 6820
rect 26881 6817 26893 6820
rect 26927 6817 26939 6851
rect 26881 6811 26939 6817
rect 28258 6808 28264 6860
rect 28316 6808 28322 6860
rect 28552 6848 28580 6876
rect 28905 6851 28963 6857
rect 28905 6848 28917 6851
rect 28552 6820 28917 6848
rect 28905 6817 28917 6820
rect 28951 6817 28963 6851
rect 29012 6848 29040 6944
rect 29181 6851 29239 6857
rect 29181 6848 29193 6851
rect 29012 6820 29193 6848
rect 28905 6811 28963 6817
rect 29181 6817 29193 6820
rect 29227 6817 29239 6851
rect 29181 6811 29239 6817
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 25130 6780 25136 6792
rect 24627 6752 25136 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25556 6752 25605 6780
rect 25556 6740 25562 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 25593 6743 25651 6749
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 25866 6780 25872 6792
rect 25823 6752 25872 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 25866 6740 25872 6752
rect 25924 6740 25930 6792
rect 26326 6740 26332 6792
rect 26384 6740 26390 6792
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6780 27215 6783
rect 27203 6752 28212 6780
rect 27203 6749 27215 6752
rect 27157 6743 27215 6749
rect 24762 6712 24768 6724
rect 24136 6684 24768 6712
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 26344 6712 26372 6740
rect 28184 6712 28212 6752
rect 28997 6715 29055 6721
rect 28997 6712 29009 6715
rect 26344 6684 26551 6712
rect 28184 6684 29009 6712
rect 20220 6616 21496 6644
rect 20220 6604 20226 6616
rect 24670 6604 24676 6656
rect 24728 6644 24734 6656
rect 26142 6644 26148 6656
rect 24728 6616 26148 6644
rect 24728 6604 24734 6616
rect 26142 6604 26148 6616
rect 26200 6604 26206 6656
rect 26234 6604 26240 6656
rect 26292 6604 26298 6656
rect 26326 6604 26332 6656
rect 26384 6644 26390 6656
rect 26421 6647 26479 6653
rect 26421 6644 26433 6647
rect 26384 6616 26433 6644
rect 26384 6604 26390 6616
rect 26421 6613 26433 6616
rect 26467 6613 26479 6647
rect 26523 6644 26551 6684
rect 28997 6681 29009 6684
rect 29043 6681 29055 6715
rect 28997 6675 29055 6681
rect 27154 6644 27160 6656
rect 26523 6616 27160 6644
rect 26421 6607 26479 6613
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 28626 6604 28632 6656
rect 28684 6604 28690 6656
rect 552 6554 31648 6576
rect 552 6502 4285 6554
rect 4337 6502 4349 6554
rect 4401 6502 4413 6554
rect 4465 6502 4477 6554
rect 4529 6502 4541 6554
rect 4593 6502 12059 6554
rect 12111 6502 12123 6554
rect 12175 6502 12187 6554
rect 12239 6502 12251 6554
rect 12303 6502 12315 6554
rect 12367 6502 19833 6554
rect 19885 6502 19897 6554
rect 19949 6502 19961 6554
rect 20013 6502 20025 6554
rect 20077 6502 20089 6554
rect 20141 6502 27607 6554
rect 27659 6502 27671 6554
rect 27723 6502 27735 6554
rect 27787 6502 27799 6554
rect 27851 6502 27863 6554
rect 27915 6502 31648 6554
rect 552 6480 31648 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 2639 6443 2697 6449
rect 1452 6412 2084 6440
rect 1452 6400 1458 6412
rect 2056 6372 2084 6412
rect 2639 6409 2651 6443
rect 2685 6440 2697 6443
rect 2958 6440 2964 6452
rect 2685 6412 2964 6440
rect 2685 6409 2697 6412
rect 2639 6403 2697 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4246 6440 4252 6452
rect 3160 6412 4252 6440
rect 3160 6372 3188 6412
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 5350 6440 5356 6452
rect 4755 6412 5356 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5592 6412 7236 6440
rect 5592 6400 5598 6412
rect 2056 6344 3188 6372
rect 3237 6375 3295 6381
rect 3237 6341 3249 6375
rect 3283 6341 3295 6375
rect 3237 6335 3295 6341
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 3252 6304 3280 6335
rect 4062 6332 4068 6384
rect 4120 6332 4126 6384
rect 7208 6372 7236 6412
rect 7282 6400 7288 6452
rect 7340 6440 7346 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7340 6412 7665 6440
rect 7340 6400 7346 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8478 6440 8484 6452
rect 8251 6412 8484 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 9490 6440 9496 6452
rect 8628 6412 9496 6440
rect 8628 6400 8634 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 9916 6412 10609 6440
rect 9916 6400 9922 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 11514 6440 11520 6452
rect 10597 6403 10655 6409
rect 10888 6412 11520 6440
rect 8389 6375 8447 6381
rect 8389 6372 8401 6375
rect 7208 6344 8401 6372
rect 8389 6341 8401 6344
rect 8435 6341 8447 6375
rect 8389 6335 8447 6341
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 8904 6344 10180 6372
rect 8904 6332 8910 6344
rect 900 6276 2084 6304
rect 900 6264 906 6276
rect 2056 6248 2084 6276
rect 3160 6276 3280 6304
rect 1210 6196 1216 6248
rect 1268 6196 1274 6248
rect 2038 6196 2044 6248
rect 2096 6196 2102 6248
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3160 6236 3188 6276
rect 3694 6264 3700 6316
rect 3752 6264 3758 6316
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 3007 6208 3188 6236
rect 4080 6236 4108 6332
rect 5905 6307 5963 6313
rect 4264 6276 4660 6304
rect 4264 6245 4292 6276
rect 4632 6248 4660 6276
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6914 6304 6920 6316
rect 5951 6276 6920 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6914 6264 6920 6276
rect 6972 6304 6978 6316
rect 6972 6276 7512 6304
rect 6972 6264 6978 6276
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 4080 6208 4169 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 2222 6128 2228 6180
rect 2280 6128 2286 6180
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 3970 6168 3976 6180
rect 3651 6140 3976 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3620 6100 3648 6131
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4448 6168 4476 6199
rect 4172 6140 4476 6168
rect 4540 6168 4568 6199
rect 4614 6196 4620 6248
rect 4672 6196 4678 6248
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 5166 6236 5172 6248
rect 4908 6208 5172 6236
rect 4908 6168 4936 6208
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5684 6208 5733 6236
rect 5684 6196 5690 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7248 6208 7314 6236
rect 7248 6196 7254 6208
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 4540 6140 4936 6168
rect 5000 6140 6193 6168
rect 4172 6112 4200 6140
rect 2924 6072 3648 6100
rect 2924 6060 2930 6072
rect 4154 6060 4160 6112
rect 4212 6060 4218 6112
rect 5000 6109 5028 6140
rect 6181 6137 6193 6140
rect 6227 6137 6239 6171
rect 6181 6131 6239 6137
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6069 5043 6103
rect 4985 6063 5043 6069
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 7484 6100 7512 6276
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7616 6276 8156 6304
rect 7616 6264 7622 6276
rect 7742 6196 7748 6248
rect 7800 6196 7806 6248
rect 7834 6196 7840 6248
rect 7892 6196 7898 6248
rect 8018 6196 8024 6248
rect 8076 6196 8082 6248
rect 8128 6168 8156 6276
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9030 6304 9036 6316
rect 8628 6276 9036 6304
rect 8628 6264 8634 6276
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9732 6276 9781 6304
rect 9732 6264 9738 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9272 6208 9965 6236
rect 9272 6196 9278 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10046 6239 10104 6245
rect 10046 6205 10058 6239
rect 10092 6205 10104 6239
rect 10152 6236 10180 6344
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10888 6313 10916 6412
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12986 6440 12992 6452
rect 12032 6412 12992 6440
rect 12032 6400 12038 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 14001 6443 14059 6449
rect 14001 6409 14013 6443
rect 14047 6440 14059 6443
rect 14090 6440 14096 6452
rect 14047 6412 14096 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 14734 6440 14740 6452
rect 14424 6412 14740 6440
rect 14424 6400 14430 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 15746 6400 15752 6452
rect 15804 6400 15810 6452
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6409 16635 6443
rect 16577 6403 16635 6409
rect 16761 6443 16819 6449
rect 16761 6409 16773 6443
rect 16807 6440 16819 6443
rect 17678 6440 17684 6452
rect 16807 6412 17684 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 11425 6375 11483 6381
rect 11425 6341 11437 6375
rect 11471 6372 11483 6375
rect 11882 6372 11888 6384
rect 11471 6344 11888 6372
rect 11471 6341 11483 6344
rect 11425 6335 11483 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 15764 6372 15792 6400
rect 13955 6344 15792 6372
rect 15841 6375 15899 6381
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 15841 6341 15853 6375
rect 15887 6341 15899 6375
rect 16592 6372 16620 6403
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 17770 6400 17776 6452
rect 17828 6400 17834 6452
rect 17862 6400 17868 6452
rect 17920 6400 17926 6452
rect 18046 6400 18052 6452
rect 18104 6400 18110 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18656 6412 21128 6440
rect 18656 6400 18662 6412
rect 16592 6344 17080 6372
rect 15841 6335 15899 6341
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10284 6276 10885 6304
rect 10284 6264 10290 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11238 6304 11244 6316
rect 11011 6276 11244 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11238 6264 11244 6276
rect 11296 6304 11302 6316
rect 11563 6307 11621 6313
rect 11563 6304 11575 6307
rect 11296 6276 11575 6304
rect 11296 6264 11302 6276
rect 11563 6273 11575 6276
rect 11609 6273 11621 6307
rect 11563 6267 11621 6273
rect 13354 6264 13360 6316
rect 13412 6264 13418 6316
rect 13707 6307 13765 6313
rect 13707 6273 13719 6307
rect 13753 6304 13765 6307
rect 14182 6304 14188 6316
rect 13753 6276 14188 6304
rect 13753 6273 13765 6276
rect 13707 6267 13765 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14608 6276 14657 6304
rect 14608 6264 14614 6276
rect 14645 6273 14657 6276
rect 14691 6304 14703 6307
rect 15010 6304 15016 6316
rect 14691 6276 15016 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 15010 6264 15016 6276
rect 15068 6304 15074 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15068 6276 15301 6304
rect 15068 6264 15074 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15856 6304 15884 6335
rect 16666 6304 16672 6316
rect 15856 6276 16672 6304
rect 15289 6267 15347 6273
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 10418 6239 10476 6245
rect 10418 6236 10430 6239
rect 10152 6208 10430 6236
rect 10046 6199 10104 6205
rect 10418 6205 10430 6208
rect 10464 6205 10476 6239
rect 12989 6239 13047 6245
rect 10418 6199 10476 6205
rect 10612 6208 11376 6236
rect 10060 6168 10088 6199
rect 8128 6140 10088 6168
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 10321 6171 10379 6177
rect 10321 6137 10333 6171
rect 10367 6168 10379 6171
rect 10612 6168 10640 6208
rect 11348 6180 11376 6208
rect 12989 6205 13001 6239
rect 13035 6236 13047 6239
rect 13078 6236 13084 6248
rect 13035 6208 13084 6236
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13648 6208 13829 6236
rect 10367 6140 10640 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 8018 6100 8024 6112
rect 7484 6072 8024 6100
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8754 6060 8760 6112
rect 8812 6060 8818 6112
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 8895 6072 9229 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10244 6100 10272 6131
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10744 6140 11069 6168
rect 10744 6128 10750 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 9548 6072 10272 6100
rect 11072 6100 11100 6131
rect 11330 6128 11336 6180
rect 11388 6128 11394 6180
rect 12618 6128 12624 6180
rect 12676 6128 12682 6180
rect 13648 6112 13676 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 14056 6208 14105 6236
rect 14056 6196 14062 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14332 6208 14381 6236
rect 14332 6196 14338 6208
rect 14369 6205 14381 6208
rect 14415 6233 14427 6239
rect 15102 6236 15108 6248
rect 14567 6233 15108 6236
rect 14415 6208 15108 6233
rect 14415 6205 14595 6208
rect 14369 6199 14427 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 15378 6128 15384 6180
rect 15436 6128 15442 6180
rect 15562 6128 15568 6180
rect 15620 6128 15626 6180
rect 16316 6112 16344 6199
rect 17052 6180 17080 6344
rect 17788 6304 17816 6400
rect 18064 6304 18092 6400
rect 18138 6332 18144 6384
rect 18196 6372 18202 6384
rect 19702 6372 19708 6384
rect 18196 6344 19708 6372
rect 18196 6332 18202 6344
rect 19702 6332 19708 6344
rect 19760 6372 19766 6384
rect 21100 6372 21128 6412
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 23385 6443 23443 6449
rect 21232 6412 23060 6440
rect 21232 6400 21238 6412
rect 21266 6372 21272 6384
rect 19760 6344 20024 6372
rect 21100 6344 21272 6372
rect 19760 6332 19766 6344
rect 19996 6304 20024 6344
rect 21266 6332 21272 6344
rect 21324 6332 21330 6384
rect 21358 6332 21364 6384
rect 21416 6372 21422 6384
rect 23032 6372 23060 6412
rect 23385 6409 23397 6443
rect 23431 6440 23443 6443
rect 25866 6440 25872 6452
rect 23431 6412 25872 6440
rect 23431 6409 23443 6412
rect 23385 6403 23443 6409
rect 25866 6400 25872 6412
rect 25924 6400 25930 6452
rect 26234 6400 26240 6452
rect 26292 6440 26298 6452
rect 28166 6440 28172 6452
rect 26292 6412 28172 6440
rect 26292 6400 26298 6412
rect 28166 6400 28172 6412
rect 28224 6400 28230 6452
rect 28350 6400 28356 6452
rect 28408 6400 28414 6452
rect 28626 6400 28632 6452
rect 28684 6400 28690 6452
rect 21416 6344 22968 6372
rect 23032 6344 24067 6372
rect 21416 6332 21422 6344
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 17604 6276 17816 6304
rect 17972 6276 19932 6304
rect 19996 6276 20085 6304
rect 17604 6245 17632 6276
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17773 6239 17831 6245
rect 17773 6205 17785 6239
rect 17819 6236 17831 6239
rect 17972 6236 18000 6276
rect 17819 6208 18000 6236
rect 18049 6239 18107 6245
rect 17819 6205 17831 6208
rect 17773 6199 17831 6205
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 18187 6208 18368 6236
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 17034 6128 17040 6180
rect 17092 6168 17098 6180
rect 17405 6171 17463 6177
rect 17405 6168 17417 6171
rect 17092 6140 17417 6168
rect 17092 6128 17098 6140
rect 17405 6137 17417 6140
rect 17451 6137 17463 6171
rect 17405 6131 17463 6137
rect 13630 6100 13636 6112
rect 11072 6072 13636 6100
rect 9548 6060 9554 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 14918 6060 14924 6112
rect 14976 6060 14982 6112
rect 16298 6060 16304 6112
rect 16356 6060 16362 6112
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 18064 6100 18092 6199
rect 18340 6180 18368 6208
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18564 6208 19748 6236
rect 18564 6196 18570 6208
rect 18230 6128 18236 6180
rect 18288 6128 18294 6180
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 19242 6168 19248 6180
rect 18380 6140 19248 6168
rect 18380 6128 18386 6140
rect 19242 6128 19248 6140
rect 19300 6128 19306 6180
rect 16540 6072 18092 6100
rect 16540 6060 16546 6072
rect 19610 6060 19616 6112
rect 19668 6060 19674 6112
rect 19720 6100 19748 6208
rect 19794 6196 19800 6248
rect 19852 6196 19858 6248
rect 19904 6168 19932 6276
rect 20073 6273 20085 6276
rect 20119 6304 20131 6307
rect 20254 6304 20260 6316
rect 20119 6276 20260 6304
rect 20119 6273 20131 6276
rect 20073 6267 20131 6273
rect 20254 6264 20260 6276
rect 20312 6304 20318 6316
rect 20312 6276 20392 6304
rect 20312 6264 20318 6276
rect 19978 6196 19984 6248
rect 20036 6236 20042 6248
rect 20364 6245 20392 6276
rect 21726 6264 21732 6316
rect 21784 6264 21790 6316
rect 22462 6264 22468 6316
rect 22520 6304 22526 6316
rect 22940 6313 22968 6344
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 22520 6276 22845 6304
rect 22520 6264 22526 6276
rect 22833 6273 22845 6276
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6273 22983 6307
rect 22925 6267 22983 6273
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 20036 6208 20177 6236
rect 20036 6196 20042 6208
rect 20165 6205 20177 6208
rect 20211 6205 20223 6239
rect 20165 6199 20223 6205
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20349 6199 20407 6205
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6236 21051 6239
rect 21082 6236 21088 6248
rect 21039 6208 21088 6236
rect 21039 6205 21051 6208
rect 20993 6199 21051 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 21315 6208 21373 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21361 6205 21373 6208
rect 21407 6236 21419 6239
rect 21744 6236 21772 6264
rect 24039 6248 24067 6344
rect 25130 6332 25136 6384
rect 25188 6372 25194 6384
rect 25958 6372 25964 6384
rect 25188 6344 25964 6372
rect 25188 6332 25194 6344
rect 25958 6332 25964 6344
rect 26016 6332 26022 6384
rect 28368 6372 28396 6400
rect 27448 6344 28396 6372
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 24504 6276 24593 6304
rect 21407 6208 21772 6236
rect 21407 6205 21419 6208
rect 21361 6199 21419 6205
rect 20070 6168 20076 6180
rect 19904 6140 20076 6168
rect 20070 6128 20076 6140
rect 20128 6168 20134 6180
rect 20257 6171 20315 6177
rect 20257 6168 20269 6171
rect 20128 6140 20269 6168
rect 20128 6128 20134 6140
rect 20257 6137 20269 6140
rect 20303 6168 20315 6171
rect 20530 6168 20536 6180
rect 20303 6140 20536 6168
rect 20303 6137 20315 6140
rect 20257 6131 20315 6137
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 21192 6168 21220 6199
rect 21818 6196 21824 6248
rect 21876 6196 21882 6248
rect 22002 6196 22008 6248
rect 22060 6196 22066 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 24026 6245 24032 6248
rect 24024 6236 24032 6245
rect 22152 6208 23888 6236
rect 23987 6208 24032 6236
rect 22152 6196 22158 6208
rect 21634 6168 21640 6180
rect 20732 6140 21640 6168
rect 20732 6100 20760 6140
rect 21634 6128 21640 6140
rect 21692 6168 21698 6180
rect 22020 6168 22048 6196
rect 21692 6140 22048 6168
rect 21692 6128 21698 6140
rect 22830 6128 22836 6180
rect 22888 6168 22894 6180
rect 22925 6171 22983 6177
rect 22925 6168 22937 6171
rect 22888 6140 22937 6168
rect 22888 6128 22894 6140
rect 22925 6137 22937 6140
rect 22971 6137 22983 6171
rect 22925 6131 22983 6137
rect 19720 6072 20760 6100
rect 20809 6103 20867 6109
rect 20809 6069 20821 6103
rect 20855 6100 20867 6103
rect 22186 6100 22192 6112
rect 20855 6072 22192 6100
rect 20855 6069 20867 6072
rect 20809 6063 20867 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22462 6060 22468 6112
rect 22520 6100 22526 6112
rect 23860 6109 23888 6208
rect 24024 6199 24032 6208
rect 24026 6196 24032 6199
rect 24084 6196 24090 6248
rect 24394 6236 24400 6248
rect 24355 6208 24400 6236
rect 24394 6196 24400 6208
rect 24452 6196 24458 6248
rect 24504 6245 24532 6276
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 24581 6267 24639 6273
rect 24762 6264 24768 6316
rect 24820 6304 24826 6316
rect 24820 6276 26464 6304
rect 24820 6264 24826 6276
rect 24489 6239 24547 6245
rect 24489 6205 24501 6239
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24728 6208 24869 6236
rect 24728 6196 24734 6208
rect 24857 6205 24869 6208
rect 24903 6205 24915 6239
rect 24857 6199 24915 6205
rect 24946 6196 24952 6248
rect 25004 6196 25010 6248
rect 25041 6239 25099 6245
rect 25041 6205 25053 6239
rect 25087 6205 25099 6239
rect 25041 6199 25099 6205
rect 24118 6128 24124 6180
rect 24176 6128 24182 6180
rect 24213 6171 24271 6177
rect 24213 6137 24225 6171
rect 24259 6137 24271 6171
rect 25056 6168 25084 6199
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25188 6208 25237 6236
rect 25188 6196 25194 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 25314 6196 25320 6248
rect 25372 6236 25378 6248
rect 25501 6239 25559 6245
rect 25501 6236 25513 6239
rect 25372 6208 25513 6236
rect 25372 6196 25378 6208
rect 25501 6205 25513 6208
rect 25547 6205 25559 6239
rect 25501 6199 25559 6205
rect 25590 6196 25596 6248
rect 25648 6196 25654 6248
rect 25682 6196 25688 6248
rect 25740 6196 25746 6248
rect 25774 6196 25780 6248
rect 25832 6196 25838 6248
rect 26436 6245 26464 6276
rect 26145 6239 26203 6245
rect 26145 6205 26157 6239
rect 26191 6205 26203 6239
rect 26145 6199 26203 6205
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 25961 6171 26019 6177
rect 25961 6168 25973 6171
rect 25056 6140 25973 6168
rect 24213 6131 24271 6137
rect 25961 6137 25973 6140
rect 26007 6137 26019 6171
rect 25961 6131 26019 6137
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22520 6072 22661 6100
rect 22520 6060 22526 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 23845 6103 23903 6109
rect 23845 6069 23857 6103
rect 23891 6069 23903 6103
rect 24228 6100 24256 6131
rect 25130 6100 25136 6112
rect 24228 6072 25136 6100
rect 23845 6063 23903 6069
rect 25130 6060 25136 6072
rect 25188 6060 25194 6112
rect 25314 6060 25320 6112
rect 25372 6060 25378 6112
rect 25590 6060 25596 6112
rect 25648 6100 25654 6112
rect 26160 6100 26188 6199
rect 26694 6196 26700 6248
rect 26752 6196 26758 6248
rect 27154 6196 27160 6248
rect 27212 6196 27218 6248
rect 27338 6196 27344 6248
rect 27396 6236 27402 6248
rect 27448 6245 27476 6344
rect 28644 6304 28672 6400
rect 27540 6276 28396 6304
rect 28644 6276 28856 6304
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 27396 6208 27445 6236
rect 27396 6196 27402 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 27433 6199 27491 6205
rect 27172 6168 27200 6196
rect 27540 6168 27568 6276
rect 28074 6196 28080 6248
rect 28132 6196 28138 6248
rect 28368 6180 28396 6276
rect 28629 6239 28687 6245
rect 28629 6205 28641 6239
rect 28675 6236 28687 6239
rect 28718 6236 28724 6248
rect 28675 6208 28724 6236
rect 28675 6205 28687 6208
rect 28629 6199 28687 6205
rect 27172 6140 27568 6168
rect 27614 6128 27620 6180
rect 27672 6168 27678 6180
rect 27982 6168 27988 6180
rect 27672 6140 27988 6168
rect 27672 6128 27678 6140
rect 27982 6128 27988 6140
rect 28040 6128 28046 6180
rect 28350 6128 28356 6180
rect 28408 6128 28414 6180
rect 28644 6168 28672 6199
rect 28718 6196 28724 6208
rect 28776 6196 28782 6248
rect 28828 6245 28856 6276
rect 28813 6239 28871 6245
rect 28813 6205 28825 6239
rect 28859 6236 28871 6239
rect 29362 6236 29368 6248
rect 28859 6208 29368 6236
rect 28859 6205 28871 6208
rect 28813 6199 28871 6205
rect 29362 6196 29368 6208
rect 29420 6196 29426 6248
rect 28644 6140 29684 6168
rect 29656 6112 29684 6140
rect 25648 6072 26188 6100
rect 25648 6060 25654 6072
rect 26234 6060 26240 6112
rect 26292 6100 26298 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 26292 6072 26341 6100
rect 26292 6060 26298 6072
rect 26329 6069 26341 6072
rect 26375 6100 26387 6103
rect 26602 6100 26608 6112
rect 26375 6072 26608 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 26602 6060 26608 6072
rect 26660 6060 26666 6112
rect 26970 6060 26976 6112
rect 27028 6100 27034 6112
rect 28721 6103 28779 6109
rect 28721 6100 28733 6103
rect 27028 6072 28733 6100
rect 27028 6060 27034 6072
rect 28721 6069 28733 6072
rect 28767 6069 28779 6103
rect 28721 6063 28779 6069
rect 28994 6060 29000 6112
rect 29052 6100 29058 6112
rect 29089 6103 29147 6109
rect 29089 6100 29101 6103
rect 29052 6072 29101 6100
rect 29052 6060 29058 6072
rect 29089 6069 29101 6072
rect 29135 6069 29147 6103
rect 29089 6063 29147 6069
rect 29638 6060 29644 6112
rect 29696 6060 29702 6112
rect 552 6010 31808 6032
rect 552 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 15946 6010
rect 15998 5958 16010 6010
rect 16062 5958 16074 6010
rect 16126 5958 16138 6010
rect 16190 5958 16202 6010
rect 16254 5958 23720 6010
rect 23772 5958 23784 6010
rect 23836 5958 23848 6010
rect 23900 5958 23912 6010
rect 23964 5958 23976 6010
rect 24028 5958 31494 6010
rect 31546 5958 31558 6010
rect 31610 5958 31622 6010
rect 31674 5958 31686 6010
rect 31738 5958 31750 6010
rect 31802 5958 31808 6010
rect 552 5936 31808 5958
rect 1486 5856 1492 5908
rect 1544 5856 1550 5908
rect 1946 5896 1952 5908
rect 1780 5868 1952 5896
rect 750 5788 756 5840
rect 808 5828 814 5840
rect 1121 5831 1179 5837
rect 808 5800 1072 5828
rect 808 5788 814 5800
rect 937 5763 995 5769
rect 937 5729 949 5763
rect 983 5729 995 5763
rect 937 5723 995 5729
rect 952 5556 980 5723
rect 1044 5692 1072 5800
rect 1121 5797 1133 5831
rect 1167 5828 1179 5831
rect 1780 5828 1808 5868
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2866 5896 2872 5908
rect 2148 5868 2872 5896
rect 1167 5800 1808 5828
rect 1167 5797 1179 5800
rect 1121 5791 1179 5797
rect 1854 5788 1860 5840
rect 1912 5788 1918 5840
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5729 1271 5763
rect 1213 5723 1271 5729
rect 1305 5763 1363 5769
rect 1305 5729 1317 5763
rect 1351 5760 1363 5763
rect 1762 5760 1768 5772
rect 1351 5732 1768 5760
rect 1351 5729 1363 5732
rect 1305 5723 1363 5729
rect 1228 5692 1256 5723
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 1964 5769 1992 5856
rect 2148 5769 2176 5868
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 4019 5899 4077 5905
rect 4019 5896 4031 5899
rect 3844 5868 4031 5896
rect 3844 5856 3850 5868
rect 4019 5865 4031 5868
rect 4065 5865 4077 5899
rect 4019 5859 4077 5865
rect 4798 5856 4804 5908
rect 4856 5856 4862 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5224 5868 5365 5896
rect 5224 5856 5230 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6181 5899 6239 5905
rect 6181 5896 6193 5899
rect 6052 5868 6193 5896
rect 6052 5856 6058 5868
rect 6181 5865 6193 5868
rect 6227 5865 6239 5899
rect 6181 5859 6239 5865
rect 6270 5856 6276 5908
rect 6328 5856 6334 5908
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 4816 5828 4844 5856
rect 6656 5828 6684 5859
rect 6914 5856 6920 5908
rect 6972 5856 6978 5908
rect 7101 5899 7159 5905
rect 7101 5865 7113 5899
rect 7147 5896 7159 5899
rect 7374 5896 7380 5908
rect 7147 5868 7380 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 7708 5868 7757 5896
rect 7708 5856 7714 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 7745 5859 7803 5865
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9214 5896 9220 5908
rect 8812 5868 9220 5896
rect 8812 5856 8818 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 9355 5868 12817 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 13630 5856 13636 5908
rect 13688 5856 13694 5908
rect 14001 5899 14059 5905
rect 14001 5865 14013 5899
rect 14047 5896 14059 5899
rect 14047 5868 14872 5896
rect 14047 5865 14059 5868
rect 14001 5859 14059 5865
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 2133 5723 2191 5729
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2682 5760 2688 5772
rect 2271 5732 2688 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 1044 5664 1256 5692
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2240 5692 2268 5723
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3620 5760 3648 5814
rect 4816 5800 6684 5828
rect 4062 5760 4068 5772
rect 3620 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4614 5760 4620 5772
rect 4304 5732 4620 5760
rect 4304 5720 4310 5732
rect 4614 5720 4620 5732
rect 4672 5760 4678 5772
rect 4709 5763 4767 5769
rect 4709 5760 4721 5763
rect 4672 5732 4721 5760
rect 4672 5720 4678 5732
rect 4709 5729 4721 5732
rect 4755 5729 4767 5763
rect 4709 5723 4767 5729
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5994 5760 6000 5772
rect 5316 5732 6000 5760
rect 5316 5720 5322 5732
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6178 5760 6184 5772
rect 6104 5732 6184 5760
rect 2096 5664 2268 5692
rect 2593 5695 2651 5701
rect 2096 5652 2102 5664
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2774 5692 2780 5704
rect 2639 5664 2780 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 3936 5664 5549 5692
rect 3936 5652 3942 5664
rect 5537 5661 5549 5664
rect 5583 5692 5595 5695
rect 6104 5692 6132 5732
rect 6178 5720 6184 5732
rect 6236 5760 6242 5772
rect 6932 5760 6960 5856
rect 8588 5828 8616 5856
rect 7305 5800 8616 5828
rect 8665 5831 8723 5837
rect 7006 5760 7012 5772
rect 6236 5732 6500 5760
rect 6932 5732 7012 5760
rect 6236 5720 6242 5732
rect 5583 5664 6132 5692
rect 6365 5695 6423 5701
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6472 5692 6500 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7305 5701 7333 5800
rect 8665 5797 8677 5831
rect 8711 5828 8723 5831
rect 9398 5828 9404 5840
rect 8711 5800 9404 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 9784 5800 10548 5828
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8754 5760 8760 5772
rect 7883 5732 8760 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9784 5769 9812 5800
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 10226 5720 10232 5772
rect 10284 5720 10290 5772
rect 10318 5720 10324 5772
rect 10376 5720 10382 5772
rect 10410 5720 10416 5772
rect 10468 5720 10474 5772
rect 10520 5760 10548 5800
rect 10686 5788 10692 5840
rect 10744 5828 10750 5840
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 10744 5800 11253 5828
rect 10744 5788 10750 5800
rect 11241 5797 11253 5800
rect 11287 5797 11299 5831
rect 12894 5828 12900 5840
rect 12466 5800 12900 5828
rect 11241 5791 11299 5797
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 13648 5828 13676 5856
rect 14277 5831 14335 5837
rect 14277 5828 14289 5831
rect 13648 5800 14289 5828
rect 14277 5797 14289 5800
rect 14323 5797 14335 5831
rect 14277 5791 14335 5797
rect 10870 5760 10876 5772
rect 10520 5732 10876 5760
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6472 5664 7297 5692
rect 6365 5655 6423 5661
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 1118 5584 1124 5636
rect 1176 5624 1182 5636
rect 1581 5627 1639 5633
rect 1581 5624 1593 5627
rect 1176 5596 1593 5624
rect 1176 5584 1182 5596
rect 1581 5593 1593 5596
rect 1627 5593 1639 5627
rect 1581 5587 1639 5593
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 5813 5627 5871 5633
rect 5813 5624 5825 5627
rect 5040 5596 5825 5624
rect 5040 5584 5046 5596
rect 5813 5593 5825 5596
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 6380 5624 6408 5655
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7524 5664 7573 5692
rect 7524 5652 7530 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 7561 5655 7619 5661
rect 8404 5664 9413 5692
rect 8404 5633 8432 5664
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10244 5692 10272 5720
rect 10183 5664 10272 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10980 5636 11008 5723
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 14185 5763 14243 5769
rect 13044 5732 13952 5760
rect 13044 5720 13050 5732
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 11388 5664 13369 5692
rect 11388 5652 11394 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 13817 5695 13875 5701
rect 13817 5661 13829 5695
rect 13863 5661 13875 5695
rect 13924 5692 13952 5732
rect 14185 5729 14197 5763
rect 14231 5760 14243 5763
rect 14366 5760 14372 5772
rect 14231 5732 14372 5760
rect 14231 5729 14243 5732
rect 14185 5723 14243 5729
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 14552 5763 14610 5769
rect 14552 5760 14564 5763
rect 14516 5732 14564 5760
rect 14516 5720 14522 5732
rect 14552 5729 14564 5732
rect 14598 5729 14610 5763
rect 14552 5723 14610 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 14660 5692 14688 5723
rect 14734 5720 14740 5772
rect 14792 5720 14798 5772
rect 14844 5760 14872 5868
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18230 5896 18236 5908
rect 18187 5868 18236 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 18524 5868 19625 5896
rect 14936 5828 14964 5856
rect 14936 5800 15516 5828
rect 15488 5769 15516 5800
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 17865 5831 17923 5837
rect 15896 5800 17540 5828
rect 15896 5788 15902 5800
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 14844 5732 14933 5760
rect 14921 5729 14933 5732
rect 14967 5760 14979 5763
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 14967 5732 15025 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5729 15531 5763
rect 15473 5723 15531 5729
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5760 17003 5763
rect 17034 5760 17040 5772
rect 16991 5732 17040 5760
rect 16991 5729 17003 5732
rect 16945 5723 17003 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 16114 5692 16120 5704
rect 13924 5664 14595 5692
rect 14660 5664 16120 5692
rect 13817 5655 13875 5661
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 6144 5596 8401 5624
rect 6144 5584 6150 5596
rect 7760 5568 7788 5596
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 9953 5627 10011 5633
rect 9953 5593 9965 5627
rect 9999 5624 10011 5627
rect 9999 5596 10916 5624
rect 9999 5593 10011 5596
rect 9953 5587 10011 5593
rect 3786 5556 3792 5568
rect 952 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4890 5516 4896 5568
rect 4948 5516 4954 5568
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7984 5528 8217 5556
rect 7984 5516 7990 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 8849 5559 8907 5565
rect 8849 5556 8861 5559
rect 8628 5528 8861 5556
rect 8628 5516 8634 5528
rect 8849 5525 8861 5528
rect 8895 5525 8907 5559
rect 8849 5519 8907 5525
rect 10778 5516 10784 5568
rect 10836 5516 10842 5568
rect 10888 5556 10916 5596
rect 10962 5584 10968 5636
rect 11020 5584 11026 5636
rect 12802 5624 12808 5636
rect 12406 5596 12808 5624
rect 12406 5556 12434 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 10888 5528 12434 5556
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 13464 5556 13492 5652
rect 13832 5624 13860 5655
rect 14567 5624 14595 5664
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 16356 5664 16681 5692
rect 16356 5652 16362 5664
rect 16669 5661 16681 5664
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 17512 5624 17540 5800
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 17911 5800 18337 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18325 5791 18383 5797
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17604 5692 17632 5723
rect 17770 5720 17776 5772
rect 17828 5720 17834 5772
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18012 5732 18184 5760
rect 18012 5720 18018 5732
rect 18046 5692 18052 5704
rect 17604 5664 18052 5692
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18156 5692 18184 5732
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 18288 5732 18429 5760
rect 18288 5720 18294 5732
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 18524 5692 18552 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 18874 5788 18880 5840
rect 18932 5788 18938 5840
rect 19628 5828 19656 5859
rect 19794 5856 19800 5908
rect 19852 5896 19858 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 19852 5868 20177 5896
rect 19852 5856 19858 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 21174 5896 21180 5908
rect 20165 5859 20223 5865
rect 20456 5868 21180 5896
rect 19978 5828 19984 5840
rect 19628 5800 19984 5828
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20456 5837 20484 5868
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 22370 5856 22376 5908
rect 22428 5856 22434 5908
rect 22922 5856 22928 5908
rect 22980 5896 22986 5908
rect 23198 5896 23204 5908
rect 22980 5868 23204 5896
rect 22980 5856 22986 5868
rect 23198 5856 23204 5868
rect 23256 5856 23262 5908
rect 24486 5896 24492 5908
rect 24228 5868 24492 5896
rect 20441 5831 20499 5837
rect 20441 5797 20453 5831
rect 20487 5797 20499 5831
rect 20441 5791 20499 5797
rect 20530 5788 20536 5840
rect 20588 5788 20594 5840
rect 22388 5828 22416 5856
rect 23845 5831 23903 5837
rect 23845 5828 23857 5831
rect 21376 5800 21772 5828
rect 18156 5664 18552 5692
rect 18892 5692 18920 5788
rect 19518 5720 19524 5772
rect 19576 5769 19582 5772
rect 19576 5763 19612 5769
rect 19600 5729 19612 5763
rect 19576 5723 19612 5729
rect 19576 5720 19582 5723
rect 20070 5720 20076 5772
rect 20128 5720 20134 5772
rect 20254 5720 20260 5772
rect 20312 5769 20318 5772
rect 20312 5763 20361 5769
rect 20312 5729 20315 5763
rect 20349 5729 20361 5763
rect 20312 5723 20361 5729
rect 20312 5720 20318 5723
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 20716 5763 20774 5769
rect 20716 5760 20728 5763
rect 20680 5732 20728 5760
rect 20680 5720 20686 5732
rect 20716 5729 20728 5732
rect 20762 5729 20774 5763
rect 20716 5723 20774 5729
rect 20809 5763 20867 5769
rect 20809 5729 20821 5763
rect 20855 5760 20867 5763
rect 20898 5760 20904 5772
rect 20855 5732 20904 5760
rect 20855 5729 20867 5732
rect 20809 5723 20867 5729
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21376 5769 21404 5800
rect 21744 5772 21772 5800
rect 22204 5800 23857 5828
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5729 21419 5763
rect 21361 5723 21419 5729
rect 21545 5763 21603 5769
rect 21545 5729 21557 5763
rect 21591 5729 21603 5763
rect 21545 5723 21603 5729
rect 19702 5692 19708 5704
rect 18892 5664 19708 5692
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21560 5692 21588 5723
rect 21634 5720 21640 5772
rect 21692 5720 21698 5772
rect 21726 5720 21732 5772
rect 21784 5720 21790 5772
rect 21818 5720 21824 5772
rect 21876 5720 21882 5772
rect 22204 5769 22232 5800
rect 23845 5797 23857 5800
rect 23891 5828 23903 5831
rect 24118 5828 24124 5840
rect 23891 5800 24124 5828
rect 23891 5797 23903 5800
rect 23845 5791 23903 5797
rect 24118 5788 24124 5800
rect 24176 5788 24182 5840
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 22373 5763 22431 5769
rect 22373 5729 22385 5763
rect 22419 5760 22431 5763
rect 22554 5760 22560 5772
rect 22419 5732 22560 5760
rect 22419 5729 22431 5732
rect 22373 5723 22431 5729
rect 22554 5720 22560 5732
rect 22612 5760 22618 5772
rect 22612 5732 22784 5760
rect 22612 5720 22618 5732
rect 21836 5692 21864 5720
rect 22756 5692 22784 5732
rect 22830 5720 22836 5772
rect 22888 5760 22894 5772
rect 23385 5763 23443 5769
rect 23385 5760 23397 5763
rect 22888 5732 23397 5760
rect 22888 5720 22894 5732
rect 23385 5729 23397 5732
rect 23431 5729 23443 5763
rect 23385 5723 23443 5729
rect 23474 5720 23480 5772
rect 23532 5720 23538 5772
rect 23566 5720 23572 5772
rect 23624 5760 23630 5772
rect 24228 5769 24256 5868
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 25130 5856 25136 5908
rect 25188 5856 25194 5908
rect 25222 5856 25228 5908
rect 25280 5896 25286 5908
rect 25869 5899 25927 5905
rect 25280 5868 25728 5896
rect 25280 5856 25286 5868
rect 25148 5828 25176 5856
rect 25317 5831 25375 5837
rect 25317 5828 25329 5831
rect 25148 5800 25329 5828
rect 25317 5797 25329 5800
rect 25363 5797 25375 5831
rect 25317 5791 25375 5797
rect 24029 5763 24087 5769
rect 24029 5760 24041 5763
rect 23624 5732 24041 5760
rect 23624 5720 23630 5732
rect 24029 5729 24041 5732
rect 24075 5729 24087 5763
rect 24029 5723 24087 5729
rect 24213 5763 24271 5769
rect 24213 5729 24225 5763
rect 24259 5729 24271 5763
rect 24213 5723 24271 5729
rect 24397 5763 24455 5769
rect 24397 5729 24409 5763
rect 24443 5760 24455 5763
rect 24443 5732 24808 5760
rect 24443 5729 24455 5732
rect 24397 5723 24455 5729
rect 23198 5692 23204 5704
rect 21140 5664 21864 5692
rect 22066 5664 22692 5692
rect 22756 5664 23204 5692
rect 21140 5652 21146 5664
rect 18966 5624 18972 5636
rect 13832 5596 14504 5624
rect 14567 5596 16896 5624
rect 17512 5596 18972 5624
rect 12759 5528 13492 5556
rect 13817 5559 13875 5565
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 13817 5525 13829 5559
rect 13863 5556 13875 5559
rect 14274 5556 14280 5568
rect 13863 5528 14280 5556
rect 13863 5525 13875 5528
rect 13817 5519 13875 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14476 5556 14504 5596
rect 14550 5556 14556 5568
rect 14476 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 15010 5516 15016 5568
rect 15068 5556 15074 5568
rect 15657 5559 15715 5565
rect 15657 5556 15669 5559
rect 15068 5528 15669 5556
rect 15068 5516 15074 5528
rect 15657 5525 15669 5528
rect 15703 5525 15715 5559
rect 16868 5556 16896 5596
rect 18966 5584 18972 5596
rect 19024 5584 19030 5636
rect 19981 5627 20039 5633
rect 19306 5596 19564 5624
rect 19306 5556 19334 5596
rect 16868 5528 19334 5556
rect 15657 5519 15715 5525
rect 19426 5516 19432 5568
rect 19484 5516 19490 5568
rect 19536 5556 19564 5596
rect 19981 5593 19993 5627
rect 20027 5624 20039 5627
rect 21910 5624 21916 5636
rect 20027 5596 21916 5624
rect 20027 5593 20039 5596
rect 19981 5587 20039 5593
rect 21910 5584 21916 5596
rect 21968 5584 21974 5636
rect 20254 5556 20260 5568
rect 19536 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 22066 5556 22094 5664
rect 22278 5584 22284 5636
rect 22336 5624 22342 5636
rect 22557 5627 22615 5633
rect 22557 5624 22569 5627
rect 22336 5596 22569 5624
rect 22336 5584 22342 5596
rect 22557 5593 22569 5596
rect 22603 5593 22615 5627
rect 22664 5624 22692 5664
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 23290 5652 23296 5704
rect 23348 5652 23354 5704
rect 23492 5692 23520 5720
rect 24302 5692 24308 5704
rect 23492 5664 24308 5692
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24780 5692 24808 5732
rect 24854 5720 24860 5772
rect 24912 5720 24918 5772
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5729 25099 5763
rect 25041 5723 25099 5729
rect 25134 5763 25192 5769
rect 25134 5729 25146 5763
rect 25180 5760 25192 5763
rect 25222 5760 25228 5772
rect 25180 5732 25228 5760
rect 25180 5729 25192 5732
rect 25134 5723 25192 5729
rect 24946 5692 24952 5704
rect 24780 5664 24952 5692
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 25056 5624 25084 5723
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 25590 5769 25596 5772
rect 25409 5763 25467 5769
rect 25409 5729 25421 5763
rect 25455 5729 25467 5763
rect 25409 5723 25467 5729
rect 25547 5763 25596 5769
rect 25547 5729 25559 5763
rect 25593 5729 25596 5763
rect 25547 5723 25596 5729
rect 25424 5692 25452 5723
rect 25590 5720 25596 5723
rect 25648 5720 25654 5772
rect 25700 5692 25728 5868
rect 25869 5865 25881 5899
rect 25915 5896 25927 5899
rect 26234 5896 26240 5908
rect 25915 5868 26240 5896
rect 25915 5865 25927 5868
rect 25869 5859 25927 5865
rect 26234 5856 26240 5868
rect 26292 5856 26298 5908
rect 26418 5856 26424 5908
rect 26476 5856 26482 5908
rect 28537 5899 28595 5905
rect 28537 5865 28549 5899
rect 28583 5896 28595 5899
rect 28810 5896 28816 5908
rect 28583 5868 28816 5896
rect 28583 5865 28595 5868
rect 28537 5859 28595 5865
rect 26436 5828 26464 5856
rect 28074 5828 28080 5840
rect 26436 5800 26832 5828
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5750 25835 5763
rect 25958 5750 25964 5772
rect 25823 5729 25964 5750
rect 25777 5723 25964 5729
rect 25792 5722 25964 5723
rect 25958 5720 25964 5722
rect 26016 5720 26022 5772
rect 26053 5763 26111 5769
rect 26053 5729 26065 5763
rect 26099 5729 26111 5763
rect 26053 5723 26111 5729
rect 26068 5692 26096 5723
rect 26142 5720 26148 5772
rect 26200 5760 26206 5772
rect 26804 5769 26832 5800
rect 28000 5800 28080 5828
rect 26605 5763 26663 5769
rect 26605 5760 26617 5763
rect 26200 5732 26617 5760
rect 26200 5720 26206 5732
rect 26605 5729 26617 5732
rect 26651 5729 26663 5763
rect 26605 5723 26663 5729
rect 26789 5763 26847 5769
rect 26789 5729 26801 5763
rect 26835 5729 26847 5763
rect 26789 5723 26847 5729
rect 26970 5720 26976 5772
rect 27028 5760 27034 5772
rect 28000 5769 28028 5800
rect 28074 5788 28080 5800
rect 28132 5828 28138 5840
rect 28552 5828 28580 5859
rect 28810 5856 28816 5868
rect 28868 5896 28874 5908
rect 28997 5899 29055 5905
rect 28997 5896 29009 5899
rect 28868 5868 29009 5896
rect 28868 5856 28874 5868
rect 28997 5865 29009 5868
rect 29043 5865 29055 5899
rect 28997 5859 29055 5865
rect 29362 5856 29368 5908
rect 29420 5856 29426 5908
rect 28132 5800 28580 5828
rect 28132 5788 28138 5800
rect 27157 5763 27215 5769
rect 27157 5760 27169 5763
rect 27028 5732 27169 5760
rect 27028 5720 27034 5732
rect 27157 5729 27169 5732
rect 27203 5729 27215 5763
rect 27157 5723 27215 5729
rect 27985 5763 28043 5769
rect 27985 5729 27997 5763
rect 28031 5729 28043 5763
rect 27985 5723 28043 5729
rect 28442 5720 28448 5772
rect 28500 5760 28506 5772
rect 29380 5760 29408 5856
rect 29457 5763 29515 5769
rect 29457 5760 29469 5763
rect 28500 5732 29316 5760
rect 29380 5732 29469 5760
rect 28500 5720 28506 5732
rect 25424 5664 25636 5692
rect 25700 5664 26096 5692
rect 22664 5596 24624 5624
rect 22557 5587 22615 5593
rect 20588 5528 22094 5556
rect 22189 5559 22247 5565
rect 20588 5516 20594 5528
rect 22189 5525 22201 5559
rect 22235 5556 22247 5559
rect 22830 5556 22836 5568
rect 22235 5528 22836 5556
rect 22235 5525 22247 5528
rect 22189 5519 22247 5525
rect 22830 5516 22836 5528
rect 22888 5556 22894 5568
rect 22925 5559 22983 5565
rect 22925 5556 22937 5559
rect 22888 5528 22937 5556
rect 22888 5516 22894 5528
rect 22925 5525 22937 5528
rect 22971 5525 22983 5559
rect 22925 5519 22983 5525
rect 23106 5516 23112 5568
rect 23164 5516 23170 5568
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 23753 5559 23811 5565
rect 23753 5556 23765 5559
rect 23624 5528 23765 5556
rect 23624 5516 23630 5528
rect 23753 5525 23765 5528
rect 23799 5525 23811 5559
rect 23753 5519 23811 5525
rect 24486 5516 24492 5568
rect 24544 5516 24550 5568
rect 24596 5556 24624 5596
rect 25056 5596 25544 5624
rect 25056 5568 25084 5596
rect 25516 5568 25544 5596
rect 24719 5559 24777 5565
rect 24719 5556 24731 5559
rect 24596 5528 24731 5556
rect 24719 5525 24731 5528
rect 24765 5525 24777 5559
rect 24719 5519 24777 5525
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 25498 5516 25504 5568
rect 25556 5516 25562 5568
rect 25608 5556 25636 5664
rect 26510 5652 26516 5704
rect 26568 5692 26574 5704
rect 26881 5695 26939 5701
rect 26881 5692 26893 5695
rect 26568 5664 26893 5692
rect 26568 5652 26574 5664
rect 26881 5661 26893 5664
rect 26927 5661 26939 5695
rect 26881 5655 26939 5661
rect 27062 5652 27068 5704
rect 27120 5692 27126 5704
rect 27525 5695 27583 5701
rect 27525 5692 27537 5695
rect 27120 5664 27537 5692
rect 27120 5652 27126 5664
rect 27525 5661 27537 5664
rect 27571 5661 27583 5695
rect 28994 5692 29000 5704
rect 27525 5655 27583 5661
rect 28184 5664 29000 5692
rect 25685 5627 25743 5633
rect 25685 5593 25697 5627
rect 25731 5624 25743 5627
rect 26602 5624 26608 5636
rect 25731 5596 26608 5624
rect 25731 5593 25743 5596
rect 25685 5587 25743 5593
rect 26602 5584 26608 5596
rect 26660 5584 26666 5636
rect 26694 5584 26700 5636
rect 26752 5624 26758 5636
rect 28184 5633 28212 5664
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 28169 5627 28227 5633
rect 28169 5624 28181 5627
rect 26752 5596 28181 5624
rect 26752 5584 26758 5596
rect 28169 5593 28181 5596
rect 28215 5593 28227 5627
rect 28169 5587 28227 5593
rect 28721 5627 28779 5633
rect 28721 5593 28733 5627
rect 28767 5624 28779 5627
rect 29086 5624 29092 5636
rect 28767 5596 29092 5624
rect 28767 5593 28779 5596
rect 28721 5587 28779 5593
rect 29086 5584 29092 5596
rect 29144 5584 29150 5636
rect 29288 5624 29316 5732
rect 29457 5729 29469 5732
rect 29503 5729 29515 5763
rect 29457 5723 29515 5729
rect 29365 5627 29423 5633
rect 29365 5624 29377 5627
rect 29288 5596 29377 5624
rect 29365 5593 29377 5596
rect 29411 5593 29423 5627
rect 29365 5587 29423 5593
rect 25958 5556 25964 5568
rect 25608 5528 25964 5556
rect 25958 5516 25964 5528
rect 26016 5516 26022 5568
rect 26050 5516 26056 5568
rect 26108 5556 26114 5568
rect 26237 5559 26295 5565
rect 26237 5556 26249 5559
rect 26108 5528 26249 5556
rect 26108 5516 26114 5528
rect 26237 5525 26249 5528
rect 26283 5525 26295 5559
rect 26237 5519 26295 5525
rect 26421 5559 26479 5565
rect 26421 5525 26433 5559
rect 26467 5556 26479 5559
rect 26510 5556 26516 5568
rect 26467 5528 26516 5556
rect 26467 5525 26479 5528
rect 26421 5519 26479 5525
rect 26510 5516 26516 5528
rect 26568 5516 26574 5568
rect 28442 5516 28448 5568
rect 28500 5556 28506 5568
rect 28537 5559 28595 5565
rect 28537 5556 28549 5559
rect 28500 5528 28549 5556
rect 28500 5516 28506 5528
rect 28537 5525 28549 5528
rect 28583 5525 28595 5559
rect 28537 5519 28595 5525
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 28813 5559 28871 5565
rect 28813 5556 28825 5559
rect 28684 5528 28825 5556
rect 28684 5516 28690 5528
rect 28813 5525 28825 5528
rect 28859 5525 28871 5559
rect 28813 5519 28871 5525
rect 28997 5559 29055 5565
rect 28997 5525 29009 5559
rect 29043 5556 29055 5559
rect 29472 5556 29500 5723
rect 29638 5720 29644 5772
rect 29696 5720 29702 5772
rect 29043 5528 29500 5556
rect 29043 5525 29055 5528
rect 28997 5519 29055 5525
rect 29546 5516 29552 5568
rect 29604 5516 29610 5568
rect 552 5466 31648 5488
rect 552 5414 4285 5466
rect 4337 5414 4349 5466
rect 4401 5414 4413 5466
rect 4465 5414 4477 5466
rect 4529 5414 4541 5466
rect 4593 5414 12059 5466
rect 12111 5414 12123 5466
rect 12175 5414 12187 5466
rect 12239 5414 12251 5466
rect 12303 5414 12315 5466
rect 12367 5414 19833 5466
rect 19885 5414 19897 5466
rect 19949 5414 19961 5466
rect 20013 5414 20025 5466
rect 20077 5414 20089 5466
rect 20141 5414 27607 5466
rect 27659 5414 27671 5466
rect 27723 5414 27735 5466
rect 27787 5414 27799 5466
rect 27851 5414 27863 5466
rect 27915 5414 31648 5466
rect 552 5392 31648 5414
rect 4798 5352 4804 5364
rect 2746 5324 4804 5352
rect 842 5176 848 5228
rect 900 5176 906 5228
rect 2314 5216 2320 5228
rect 2240 5188 2320 5216
rect 2240 5134 2268 5188
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2746 5148 2774 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6822 5352 6828 5364
rect 6227 5324 6828 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7558 5352 7564 5364
rect 6932 5324 7564 5352
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 6457 5287 6515 5293
rect 2924 5256 4476 5284
rect 2924 5244 2930 5256
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4448 5225 4476 5256
rect 6457 5253 6469 5287
rect 6503 5284 6515 5287
rect 6932 5284 6960 5324
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 9490 5352 9496 5364
rect 7892 5324 9496 5352
rect 7892 5312 7898 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10318 5312 10324 5364
rect 10376 5312 10382 5364
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 11866 5355 11924 5361
rect 11866 5352 11878 5355
rect 10735 5324 11878 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 11866 5321 11878 5324
rect 11912 5321 11924 5355
rect 11866 5315 11924 5321
rect 13955 5355 14013 5361
rect 13955 5321 13967 5355
rect 14001 5352 14013 5355
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 14001 5324 16313 5352
rect 14001 5321 14013 5324
rect 13955 5315 14013 5321
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17681 5355 17739 5361
rect 17681 5352 17693 5355
rect 16816 5324 17693 5352
rect 16816 5312 16822 5324
rect 17681 5321 17693 5324
rect 17727 5352 17739 5355
rect 17727 5324 19380 5352
rect 17727 5321 17739 5324
rect 17681 5315 17739 5321
rect 6503 5256 6960 5284
rect 6503 5253 6515 5256
rect 6457 5247 6515 5253
rect 10962 5244 10968 5296
rect 11020 5284 11026 5296
rect 11020 5256 11652 5284
rect 11020 5244 11026 5256
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4798 5216 4804 5228
rect 4479 5188 4804 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 11425 5219 11483 5225
rect 9272 5188 10088 5216
rect 9272 5176 9278 5188
rect 2464 5120 2774 5148
rect 3053 5151 3111 5157
rect 2464 5108 2470 5120
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3697 5151 3755 5157
rect 3099 5120 3280 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 1118 5040 1124 5092
rect 1176 5040 1182 5092
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2593 5015 2651 5021
rect 2593 5012 2605 5015
rect 2464 4984 2605 5012
rect 2464 4972 2470 4984
rect 2593 4981 2605 4984
rect 2639 4981 2651 5015
rect 2593 4975 2651 4981
rect 2866 4972 2872 5024
rect 2924 4972 2930 5024
rect 3252 5021 3280 5120
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4172 5148 4200 5176
rect 3743 5120 4200 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 8205 5151 8263 5157
rect 6052 5120 6592 5148
rect 6052 5108 6058 5120
rect 4706 5040 4712 5092
rect 4764 5040 4770 5092
rect 6178 5080 6184 5092
rect 5934 5052 6184 5080
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 4981 3295 5015
rect 3237 4975 3295 4981
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 3384 4984 3617 5012
rect 3384 4972 3390 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 3605 4975 3663 4981
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 6012 5012 6040 5052
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 4120 4984 6040 5012
rect 6564 5012 6592 5120
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8251 5120 8585 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 7190 5040 7196 5092
rect 7248 5040 7254 5092
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7892 5052 7941 5080
rect 7892 5040 7898 5052
rect 7929 5049 7941 5052
rect 7975 5049 7987 5083
rect 7929 5043 7987 5049
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8220 5080 8248 5111
rect 8076 5052 8248 5080
rect 8076 5040 8082 5052
rect 8846 5040 8852 5092
rect 8904 5040 8910 5092
rect 10060 5080 10088 5188
rect 10433 5188 11192 5216
rect 10318 5080 10324 5092
rect 10060 5066 10324 5080
rect 10074 5052 10324 5066
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 10433 5012 10461 5188
rect 11164 5157 11192 5188
rect 11425 5185 11437 5219
rect 11471 5216 11483 5219
rect 11514 5216 11520 5228
rect 11471 5188 11520 5216
rect 11471 5185 11483 5188
rect 11425 5179 11483 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11624 5225 11652 5256
rect 13354 5244 13360 5296
rect 13412 5244 13418 5296
rect 14182 5244 14188 5296
rect 14240 5244 14246 5296
rect 14642 5284 14648 5296
rect 14476 5256 14648 5284
rect 11609 5219 11667 5225
rect 11609 5185 11621 5219
rect 11655 5216 11667 5219
rect 12526 5216 12532 5228
rect 11655 5188 12532 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 11149 5151 11207 5157
rect 10551 5120 10824 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10796 5021 10824 5120
rect 11149 5117 11161 5151
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 11164 5080 11192 5111
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 12952 5120 13018 5148
rect 12952 5108 12958 5120
rect 11790 5080 11796 5092
rect 11164 5052 11796 5080
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 6564 4984 10461 5012
rect 10781 5015 10839 5021
rect 4120 4972 4126 4984
rect 10781 4981 10793 5015
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11241 5015 11299 5021
rect 11241 5012 11253 5015
rect 11204 4984 11253 5012
rect 11204 4972 11210 4984
rect 11241 4981 11253 4984
rect 11287 5012 11299 5015
rect 13372 5012 13400 5244
rect 14476 5225 14504 5256
rect 14642 5244 14648 5256
rect 14700 5284 14706 5296
rect 15841 5287 15899 5293
rect 15841 5284 15853 5287
rect 14700 5256 15853 5284
rect 14700 5244 14706 5256
rect 15841 5253 15853 5256
rect 15887 5284 15899 5287
rect 16114 5284 16120 5296
rect 15887 5256 16120 5284
rect 15887 5253 15899 5256
rect 15841 5247 15899 5253
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 16850 5244 16856 5296
rect 16908 5284 16914 5296
rect 19245 5287 19303 5293
rect 19245 5284 19257 5287
rect 16908 5256 17816 5284
rect 16908 5244 16914 5256
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14461 5219 14519 5225
rect 13679 5188 14412 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13832 5157 13860 5188
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 13740 5080 13768 5111
rect 14090 5108 14096 5160
rect 14148 5108 14154 5160
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 14384 5148 14412 5188
rect 14461 5185 14473 5219
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14568 5188 15056 5216
rect 14568 5148 14596 5188
rect 14384 5120 14596 5148
rect 14631 5151 14689 5157
rect 14631 5117 14643 5151
rect 14677 5148 14689 5151
rect 14918 5148 14924 5160
rect 14677 5120 14924 5148
rect 14677 5117 14689 5120
rect 14631 5111 14689 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15028 5148 15056 5188
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 16945 5219 17003 5225
rect 15344 5188 16344 5216
rect 15344 5176 15350 5188
rect 15746 5148 15752 5160
rect 15028 5120 15752 5148
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15856 5120 16037 5148
rect 14936 5080 14964 5108
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 13740 5052 14044 5080
rect 14936 5052 15485 5080
rect 14016 5024 14044 5052
rect 15473 5049 15485 5052
rect 15519 5049 15531 5083
rect 15473 5043 15531 5049
rect 11287 4984 13400 5012
rect 11287 4981 11299 4984
rect 11241 4975 11299 4981
rect 13998 4972 14004 5024
rect 14056 4972 14062 5024
rect 14921 5015 14979 5021
rect 14921 4981 14933 5015
rect 14967 5012 14979 5015
rect 15378 5012 15384 5024
rect 14967 4984 15384 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15378 4972 15384 4984
rect 15436 5012 15442 5024
rect 15856 5012 15884 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16206 5148 16212 5160
rect 16163 5120 16212 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16316 5089 16344 5188
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17126 5216 17132 5228
rect 16991 5188 17132 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17126 5176 17132 5188
rect 17184 5216 17190 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17184 5188 17325 5216
rect 17184 5176 17190 5188
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17034 5148 17040 5160
rect 16899 5120 17040 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 17788 5157 17816 5256
rect 18340 5256 19257 5284
rect 18046 5176 18052 5228
rect 18104 5176 18110 5228
rect 18340 5225 18368 5256
rect 19245 5253 19257 5256
rect 19291 5253 19303 5287
rect 19245 5247 19303 5253
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 18414 5176 18420 5228
rect 18472 5176 18478 5228
rect 17773 5151 17831 5157
rect 17773 5117 17785 5151
rect 17819 5148 17831 5151
rect 17819 5120 18092 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 16301 5083 16359 5089
rect 15948 5052 16252 5080
rect 15948 5021 15976 5052
rect 15436 4984 15884 5012
rect 15933 5015 15991 5021
rect 15436 4972 15442 4984
rect 15933 4981 15945 5015
rect 15979 4981 15991 5015
rect 16224 5012 16252 5052
rect 16301 5049 16313 5083
rect 16347 5080 16359 5083
rect 18064 5080 18092 5120
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18432 5148 18460 5176
rect 18279 5120 18460 5148
rect 19352 5148 19380 5324
rect 19610 5312 19616 5364
rect 19668 5312 19674 5364
rect 20993 5355 21051 5361
rect 20993 5321 21005 5355
rect 21039 5352 21051 5355
rect 21726 5352 21732 5364
rect 21039 5324 21732 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 22278 5312 22284 5364
rect 22336 5312 22342 5364
rect 22741 5355 22799 5361
rect 22741 5321 22753 5355
rect 22787 5352 22799 5355
rect 23569 5355 23627 5361
rect 22787 5324 22968 5352
rect 22787 5321 22799 5324
rect 22741 5315 22799 5321
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 19760 5256 20852 5284
rect 19760 5244 19766 5256
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 20824 5225 20852 5256
rect 21082 5244 21088 5296
rect 21140 5244 21146 5296
rect 21634 5244 21640 5296
rect 21692 5244 21698 5296
rect 20809 5219 20867 5225
rect 19484 5188 19840 5216
rect 19484 5176 19490 5188
rect 19521 5151 19579 5157
rect 19352 5120 19472 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 19334 5080 19340 5092
rect 16347 5052 17908 5080
rect 18064 5052 19340 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16482 5012 16488 5024
rect 16224 4984 16488 5012
rect 15933 4975 15991 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 17218 4972 17224 5024
rect 17276 4972 17282 5024
rect 17880 5021 17908 5052
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 17865 5015 17923 5021
rect 17865 4981 17877 5015
rect 17911 4981 17923 5015
rect 17865 4975 17923 4981
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 19444 5012 19472 5120
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 19702 5148 19708 5160
rect 19567 5120 19708 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 19812 5157 19840 5188
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21100 5216 21128 5244
rect 20855 5188 21128 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 19797 5151 19855 5157
rect 19797 5117 19809 5151
rect 19843 5117 19855 5151
rect 19797 5111 19855 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5148 21143 5151
rect 21652 5148 21680 5244
rect 21913 5219 21971 5225
rect 21913 5185 21925 5219
rect 21959 5216 21971 5219
rect 22094 5216 22100 5228
rect 21959 5188 22100 5216
rect 21959 5185 21971 5188
rect 21913 5179 21971 5185
rect 22094 5176 22100 5188
rect 22152 5176 22158 5228
rect 22296 5216 22324 5312
rect 22940 5216 22968 5324
rect 23569 5321 23581 5355
rect 23615 5352 23627 5355
rect 24210 5352 24216 5364
rect 23615 5324 24216 5352
rect 23615 5321 23627 5324
rect 23569 5315 23627 5321
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 24946 5312 24952 5364
rect 25004 5312 25010 5364
rect 25317 5355 25375 5361
rect 25317 5321 25329 5355
rect 25363 5352 25375 5355
rect 25774 5352 25780 5364
rect 25363 5324 25780 5352
rect 25363 5321 25375 5324
rect 25317 5315 25375 5321
rect 25774 5312 25780 5324
rect 25832 5312 25838 5364
rect 25958 5312 25964 5364
rect 26016 5352 26022 5364
rect 26510 5352 26516 5364
rect 26016 5324 26516 5352
rect 26016 5312 26022 5324
rect 26510 5312 26516 5324
rect 26568 5312 26574 5364
rect 26694 5312 26700 5364
rect 26752 5352 26758 5364
rect 27249 5355 27307 5361
rect 27249 5352 27261 5355
rect 26752 5324 27261 5352
rect 26752 5312 26758 5324
rect 27249 5321 27261 5324
rect 27295 5321 27307 5355
rect 28626 5352 28632 5364
rect 27249 5315 27307 5321
rect 27356 5324 28632 5352
rect 23014 5244 23020 5296
rect 23072 5284 23078 5296
rect 23845 5287 23903 5293
rect 23845 5284 23857 5287
rect 23072 5256 23857 5284
rect 23072 5244 23078 5256
rect 23845 5253 23857 5256
rect 23891 5253 23903 5287
rect 24394 5284 24400 5296
rect 23845 5247 23903 5253
rect 23952 5256 24400 5284
rect 23290 5216 23296 5228
rect 22296 5188 22692 5216
rect 22940 5188 23296 5216
rect 21821 5151 21879 5157
rect 21821 5148 21833 5151
rect 21131 5120 21680 5148
rect 21744 5120 21833 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 20254 5040 20260 5092
rect 20312 5080 20318 5092
rect 21177 5083 21235 5089
rect 21177 5080 21189 5083
rect 20312 5052 21189 5080
rect 20312 5040 20318 5052
rect 21177 5049 21189 5052
rect 21223 5049 21235 5083
rect 21177 5043 21235 5049
rect 21744 5024 21772 5120
rect 21821 5117 21833 5120
rect 21867 5117 21879 5151
rect 22189 5151 22247 5157
rect 22189 5148 22201 5151
rect 21821 5111 21879 5117
rect 22066 5120 22201 5148
rect 22066 5080 22094 5120
rect 22189 5117 22201 5120
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 22370 5108 22376 5160
rect 22428 5148 22434 5160
rect 22664 5157 22692 5188
rect 23290 5176 23296 5188
rect 23348 5216 23354 5228
rect 23952 5216 23980 5256
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 24762 5244 24768 5296
rect 24820 5244 24826 5296
rect 24964 5284 24992 5312
rect 25501 5287 25559 5293
rect 25501 5284 25513 5287
rect 24964 5256 25513 5284
rect 25501 5253 25513 5256
rect 25547 5253 25559 5287
rect 25501 5247 25559 5253
rect 24857 5219 24915 5225
rect 23348 5188 23980 5216
rect 24136 5188 24808 5216
rect 23348 5176 23354 5188
rect 22649 5151 22707 5157
rect 22428 5120 22600 5148
rect 22428 5108 22434 5120
rect 21836 5052 22094 5080
rect 21836 5024 21864 5052
rect 20438 5012 20444 5024
rect 19300 4984 20444 5012
rect 19300 4972 19306 4984
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 20530 4972 20536 5024
rect 20588 4972 20594 5024
rect 21726 4972 21732 5024
rect 21784 4972 21790 5024
rect 21818 4972 21824 5024
rect 21876 4972 21882 5024
rect 22462 4972 22468 5024
rect 22520 4972 22526 5024
rect 22572 5012 22600 5120
rect 22649 5117 22661 5151
rect 22695 5117 22707 5151
rect 22649 5111 22707 5117
rect 22830 5108 22836 5160
rect 22888 5108 22894 5160
rect 22922 5108 22928 5160
rect 22980 5148 22986 5160
rect 23860 5157 24072 5158
rect 24136 5157 24164 5188
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 22980 5120 23029 5148
rect 22980 5108 22986 5120
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 23017 5111 23075 5117
rect 23109 5151 23167 5157
rect 23109 5117 23121 5151
rect 23155 5148 23167 5151
rect 23860 5151 24087 5157
rect 23860 5148 24041 5151
rect 23155 5130 24041 5148
rect 23155 5120 23888 5130
rect 23155 5117 23167 5120
rect 23109 5111 23167 5117
rect 24029 5117 24041 5130
rect 24075 5117 24087 5151
rect 24029 5111 24087 5117
rect 24121 5151 24179 5157
rect 24121 5117 24133 5151
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 22848 5080 22876 5108
rect 23124 5080 23152 5111
rect 22848 5052 23152 5080
rect 23198 5040 23204 5092
rect 23256 5080 23262 5092
rect 23293 5083 23351 5089
rect 23293 5080 23305 5083
rect 23256 5052 23305 5080
rect 23256 5040 23262 5052
rect 23293 5049 23305 5052
rect 23339 5049 23351 5083
rect 23293 5043 23351 5049
rect 23382 5040 23388 5092
rect 23440 5080 23446 5092
rect 23477 5083 23535 5089
rect 23477 5080 23489 5083
rect 23440 5052 23489 5080
rect 23440 5040 23446 5052
rect 23477 5049 23489 5052
rect 23523 5049 23535 5083
rect 23477 5043 23535 5049
rect 23842 5040 23848 5092
rect 23900 5040 23906 5092
rect 24394 5040 24400 5092
rect 24452 5040 24458 5092
rect 24780 5080 24808 5188
rect 24857 5185 24869 5219
rect 24903 5216 24915 5219
rect 25593 5219 25651 5225
rect 25593 5216 25605 5219
rect 24903 5188 25605 5216
rect 24903 5185 24915 5188
rect 24857 5179 24915 5185
rect 25593 5185 25605 5188
rect 25639 5185 25651 5219
rect 25792 5216 25820 5312
rect 27356 5216 27384 5324
rect 28626 5312 28632 5324
rect 28684 5312 28690 5364
rect 25792 5188 26832 5216
rect 25593 5179 25651 5185
rect 25406 5108 25412 5160
rect 25464 5108 25470 5160
rect 25685 5151 25743 5157
rect 25685 5117 25697 5151
rect 25731 5148 25743 5151
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 25731 5120 26433 5148
rect 25731 5117 25743 5120
rect 25685 5111 25743 5117
rect 26421 5117 26433 5120
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 26602 5108 26608 5160
rect 26660 5108 26666 5160
rect 26804 5157 26832 5188
rect 26896 5188 27384 5216
rect 27985 5219 28043 5225
rect 26896 5157 26924 5188
rect 27985 5185 27997 5219
rect 28031 5216 28043 5219
rect 28074 5216 28080 5228
rect 28031 5188 28080 5216
rect 28031 5185 28043 5188
rect 27985 5179 28043 5185
rect 26789 5151 26847 5157
rect 26789 5117 26801 5151
rect 26835 5117 26847 5151
rect 26789 5111 26847 5117
rect 26881 5151 26939 5157
rect 26881 5117 26893 5151
rect 26927 5117 26939 5151
rect 27801 5151 27859 5157
rect 27801 5148 27813 5151
rect 26881 5111 26939 5117
rect 26988 5120 27813 5148
rect 25424 5080 25452 5108
rect 25869 5083 25927 5089
rect 25869 5080 25881 5083
rect 24780 5052 25360 5080
rect 25424 5052 25881 5080
rect 23934 5012 23940 5024
rect 22572 4984 23940 5012
rect 23934 4972 23940 4984
rect 23992 4972 23998 5024
rect 24412 5012 24440 5040
rect 24949 5015 25007 5021
rect 24949 5012 24961 5015
rect 24412 4984 24961 5012
rect 24949 4981 24961 4984
rect 24995 4981 25007 5015
rect 25332 5012 25360 5052
rect 25869 5049 25881 5052
rect 25915 5049 25927 5083
rect 25869 5043 25927 5049
rect 25958 5040 25964 5092
rect 26016 5080 26022 5092
rect 26694 5080 26700 5092
rect 26016 5052 26700 5080
rect 26016 5040 26022 5052
rect 26694 5040 26700 5052
rect 26752 5040 26758 5092
rect 26988 5024 27016 5120
rect 27801 5117 27813 5120
rect 27847 5117 27859 5151
rect 27801 5111 27859 5117
rect 27249 5083 27307 5089
rect 27249 5049 27261 5083
rect 27295 5080 27307 5083
rect 27338 5080 27344 5092
rect 27295 5052 27344 5080
rect 27295 5049 27307 5052
rect 27249 5043 27307 5049
rect 27338 5040 27344 5052
rect 27396 5040 27402 5092
rect 27433 5083 27491 5089
rect 27433 5049 27445 5083
rect 27479 5080 27491 5083
rect 28000 5080 28028 5179
rect 28074 5176 28080 5188
rect 28132 5176 28138 5228
rect 28276 5188 29592 5216
rect 28276 5157 28304 5188
rect 29564 5160 29592 5188
rect 28261 5151 28319 5157
rect 28261 5117 28273 5151
rect 28307 5117 28319 5151
rect 28261 5111 28319 5117
rect 28350 5108 28356 5160
rect 28408 5148 28414 5160
rect 28445 5151 28503 5157
rect 28445 5148 28457 5151
rect 28408 5120 28457 5148
rect 28408 5108 28414 5120
rect 28445 5117 28457 5120
rect 28491 5148 28503 5151
rect 28491 5120 28994 5148
rect 28491 5117 28503 5120
rect 28445 5111 28503 5117
rect 27479 5052 28028 5080
rect 27479 5049 27491 5052
rect 27433 5043 27491 5049
rect 28074 5040 28080 5092
rect 28132 5040 28138 5092
rect 28966 5080 28994 5120
rect 29086 5108 29092 5160
rect 29144 5148 29150 5160
rect 29457 5151 29515 5157
rect 29457 5148 29469 5151
rect 29144 5120 29469 5148
rect 29144 5108 29150 5120
rect 29457 5117 29469 5120
rect 29503 5117 29515 5151
rect 29457 5111 29515 5117
rect 29546 5108 29552 5160
rect 29604 5108 29610 5160
rect 29181 5083 29239 5089
rect 29181 5080 29193 5083
rect 28966 5052 29193 5080
rect 29181 5049 29193 5052
rect 29227 5049 29239 5083
rect 29181 5043 29239 5049
rect 29365 5083 29423 5089
rect 29365 5049 29377 5083
rect 29411 5080 29423 5083
rect 29564 5080 29592 5108
rect 29411 5052 29592 5080
rect 29411 5049 29423 5052
rect 29365 5043 29423 5049
rect 26970 5012 26976 5024
rect 25332 4984 26976 5012
rect 24949 4975 25007 4981
rect 26970 4972 26976 4984
rect 27028 4972 27034 5024
rect 27065 5015 27123 5021
rect 27065 4981 27077 5015
rect 27111 5012 27123 5015
rect 27154 5012 27160 5024
rect 27111 4984 27160 5012
rect 27111 4981 27123 4984
rect 27065 4975 27123 4981
rect 27154 4972 27160 4984
rect 27212 4972 27218 5024
rect 27614 4972 27620 5024
rect 27672 4972 27678 5024
rect 28258 4972 28264 5024
rect 28316 5012 28322 5024
rect 28997 5015 29055 5021
rect 28997 5012 29009 5015
rect 28316 4984 29009 5012
rect 28316 4972 28322 4984
rect 28997 4981 29009 4984
rect 29043 4981 29055 5015
rect 28997 4975 29055 4981
rect 29638 4972 29644 5024
rect 29696 4972 29702 5024
rect 552 4922 31808 4944
rect 552 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 15946 4922
rect 15998 4870 16010 4922
rect 16062 4870 16074 4922
rect 16126 4870 16138 4922
rect 16190 4870 16202 4922
rect 16254 4870 23720 4922
rect 23772 4870 23784 4922
rect 23836 4870 23848 4922
rect 23900 4870 23912 4922
rect 23964 4870 23976 4922
rect 24028 4870 31494 4922
rect 31546 4870 31558 4922
rect 31610 4870 31622 4922
rect 31674 4870 31686 4922
rect 31738 4870 31750 4922
rect 31802 4870 31808 4922
rect 552 4848 31808 4870
rect 1026 4768 1032 4820
rect 1084 4768 1090 4820
rect 1121 4811 1179 4817
rect 1121 4777 1133 4811
rect 1167 4808 1179 4811
rect 1210 4808 1216 4820
rect 1167 4780 1216 4808
rect 1167 4777 1179 4780
rect 1121 4771 1179 4777
rect 1210 4768 1216 4780
rect 1268 4768 1274 4820
rect 1670 4768 1676 4820
rect 1728 4768 1734 4820
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2590 4808 2596 4820
rect 2087 4780 2596 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2866 4768 2872 4820
rect 2924 4768 2930 4820
rect 4249 4811 4307 4817
rect 4249 4777 4261 4811
rect 4295 4808 4307 4811
rect 4614 4808 4620 4820
rect 4295 4780 4620 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 937 4675 995 4681
rect 937 4641 949 4675
rect 983 4672 995 4675
rect 1044 4672 1072 4768
rect 983 4644 1072 4672
rect 1397 4675 1455 4681
rect 983 4641 995 4644
rect 937 4635 995 4641
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1688 4672 1716 4768
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 2682 4740 2688 4752
rect 2188 4712 2688 4740
rect 2188 4700 2194 4712
rect 2406 4672 2412 4684
rect 1443 4644 1716 4672
rect 2148 4644 2412 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2148 4613 2176 4644
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 2516 4681 2544 4712
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 2884 4740 2912 4768
rect 4062 4740 4068 4752
rect 2823 4712 2912 4740
rect 4002 4712 4068 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4908 4672 4936 4771
rect 5258 4768 5264 4820
rect 5316 4768 5322 4820
rect 7466 4808 7472 4820
rect 6104 4780 7472 4808
rect 5994 4740 6000 4752
rect 4663 4644 4936 4672
rect 5276 4712 6000 4740
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2363 4576 2636 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 934 4496 940 4548
rect 992 4496 998 4548
rect 1026 4496 1032 4548
rect 1084 4536 1090 4548
rect 1673 4539 1731 4545
rect 1673 4536 1685 4539
rect 1084 4508 1685 4536
rect 1084 4496 1090 4508
rect 1673 4505 1685 4508
rect 1719 4505 1731 4539
rect 1673 4499 1731 4505
rect 952 4468 980 4496
rect 2608 4480 2636 4576
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 5276 4604 5304 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4672 5411 4675
rect 5810 4672 5816 4684
rect 5399 4644 5816 4672
rect 5399 4641 5411 4644
rect 5353 4635 5411 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 3384 4576 5304 4604
rect 5537 4607 5595 4613
rect 3384 4564 3390 4576
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 6104 4604 6132 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7616 4780 8125 4808
rect 7616 4768 7622 4780
rect 8113 4777 8125 4780
rect 8159 4808 8171 4811
rect 8938 4808 8944 4820
rect 8159 4780 8944 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 10962 4768 10968 4820
rect 11020 4768 11026 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 11940 4780 13308 4808
rect 11940 4768 11946 4780
rect 6181 4743 6239 4749
rect 6181 4709 6193 4743
rect 6227 4740 6239 4743
rect 6546 4740 6552 4752
rect 6227 4712 6552 4740
rect 6227 4709 6239 4712
rect 6181 4703 6239 4709
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 7190 4700 7196 4752
rect 7248 4700 7254 4752
rect 9214 4700 9220 4752
rect 9272 4700 9278 4752
rect 10980 4740 11008 4768
rect 10152 4712 11284 4740
rect 10152 4681 10180 4712
rect 11256 4684 11284 4712
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 10410 4632 10416 4684
rect 10468 4632 10474 4684
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10778 4672 10784 4684
rect 10551 4644 10784 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 12618 4632 12624 4684
rect 12676 4632 12682 4684
rect 13280 4681 13308 4780
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 14148 4780 14565 4808
rect 14148 4768 14154 4780
rect 14553 4777 14565 4780
rect 14599 4777 14611 4811
rect 14553 4771 14611 4777
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14792 4780 15025 4808
rect 14792 4768 14798 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15194 4808 15200 4820
rect 15013 4771 15071 4777
rect 15120 4780 15200 4808
rect 13906 4700 13912 4752
rect 13964 4700 13970 4752
rect 15120 4740 15148 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 15286 4768 15292 4820
rect 15344 4768 15350 4820
rect 15378 4768 15384 4820
rect 15436 4768 15442 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15528 4780 15608 4808
rect 15528 4768 15534 4780
rect 14936 4712 15148 4740
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 14458 4632 14464 4684
rect 14516 4632 14522 4684
rect 14642 4632 14648 4684
rect 14700 4632 14706 4684
rect 14936 4681 14964 4712
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4641 14795 4675
rect 14737 4635 14795 4641
rect 14921 4675 14979 4681
rect 14921 4641 14933 4675
rect 14967 4641 14979 4675
rect 14921 4635 14979 4641
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 15304 4672 15332 4768
rect 15396 4740 15424 4768
rect 15396 4712 15516 4740
rect 15243 4644 15332 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 5583 4576 6132 4604
rect 6365 4607 6423 4613
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 6380 4536 6408 4567
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 9861 4607 9919 4613
rect 7064 4576 8800 4604
rect 7064 4564 7070 4576
rect 8772 4548 8800 4576
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 9907 4576 10272 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 3936 4508 6408 4536
rect 3936 4496 3942 4508
rect 8754 4496 8760 4548
rect 8812 4496 8818 4548
rect 10244 4545 10272 4576
rect 11164 4576 11529 4604
rect 11164 4545 11192 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4573 13967 4607
rect 13909 4567 13967 4573
rect 10229 4539 10287 4545
rect 10229 4505 10241 4539
rect 10275 4505 10287 4539
rect 10229 4499 10287 4505
rect 11149 4539 11207 4545
rect 11149 4505 11161 4539
rect 11195 4505 11207 4539
rect 11149 4499 11207 4505
rect 12986 4496 12992 4548
rect 13044 4496 13050 4548
rect 13078 4496 13084 4548
rect 13136 4496 13142 4548
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 13228 4508 13461 4536
rect 13228 4496 13234 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 1213 4471 1271 4477
rect 1213 4468 1225 4471
rect 952 4440 1225 4468
rect 1213 4437 1225 4440
rect 1259 4437 1271 4471
rect 1213 4431 1271 4437
rect 2590 4428 2596 4480
rect 2648 4428 2654 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4801 4471 4859 4477
rect 4801 4468 4813 4471
rect 4672 4440 4813 4468
rect 4672 4428 4678 4440
rect 4801 4437 4813 4440
rect 4847 4437 4859 4471
rect 4801 4431 4859 4437
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6178 4468 6184 4480
rect 6135 4440 6184 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6178 4428 6184 4440
rect 6236 4468 6242 4480
rect 7006 4468 7012 4480
rect 6236 4440 7012 4468
rect 6236 4428 6242 4440
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 8389 4471 8447 4477
rect 8389 4437 8401 4471
rect 8435 4468 8447 4471
rect 9398 4468 9404 4480
rect 8435 4440 9404 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 13924 4468 13952 4567
rect 13998 4564 14004 4616
rect 14056 4564 14062 4616
rect 14476 4604 14504 4632
rect 14752 4604 14780 4635
rect 15378 4632 15384 4684
rect 15436 4632 15442 4684
rect 15488 4681 15516 4712
rect 15580 4681 15608 4780
rect 15746 4768 15752 4820
rect 15804 4768 15810 4820
rect 16758 4768 16764 4820
rect 16816 4768 16822 4820
rect 16850 4768 16856 4820
rect 16908 4768 16914 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 17589 4811 17647 4817
rect 17589 4777 17601 4811
rect 17635 4808 17647 4811
rect 17770 4808 17776 4820
rect 17635 4780 17776 4808
rect 17635 4777 17647 4780
rect 17589 4771 17647 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 18138 4768 18144 4820
rect 18196 4768 18202 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 21818 4808 21824 4820
rect 18380 4780 21824 4808
rect 18380 4768 18386 4780
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 21910 4768 21916 4820
rect 21968 4768 21974 4820
rect 23014 4808 23020 4820
rect 22388 4780 23020 4808
rect 15473 4675 15531 4681
rect 15473 4641 15485 4675
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4641 16359 4675
rect 16776 4672 16804 4768
rect 16868 4740 16896 4768
rect 17037 4743 17095 4749
rect 17037 4740 17049 4743
rect 16868 4712 17049 4740
rect 17037 4709 17049 4712
rect 17083 4709 17095 4743
rect 17037 4703 17095 4709
rect 17144 4681 17172 4768
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 18064 4740 18092 4768
rect 18233 4743 18291 4749
rect 18233 4740 18245 4743
rect 17276 4712 17816 4740
rect 18064 4712 18245 4740
rect 17276 4700 17282 4712
rect 17788 4681 17816 4712
rect 18233 4709 18245 4712
rect 18279 4709 18291 4743
rect 20625 4743 20683 4749
rect 20625 4740 20637 4743
rect 18233 4703 18291 4709
rect 19076 4712 20637 4740
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 16776 4644 16865 4672
rect 16301 4635 16359 4641
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4641 17187 4675
rect 17129 4635 17187 4641
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 18509 4675 18567 4681
rect 17819 4644 18000 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 14476 4576 14780 4604
rect 14752 4536 14780 4576
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15102 4604 15108 4616
rect 14875 4576 15108 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15102 4564 15108 4576
rect 15160 4604 15166 4616
rect 16132 4604 16160 4635
rect 15160 4576 16160 4604
rect 15160 4564 15166 4576
rect 16206 4564 16212 4616
rect 16264 4564 16270 4616
rect 15562 4536 15568 4548
rect 14752 4508 15568 4536
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 15654 4496 15660 4548
rect 15712 4536 15718 4548
rect 16316 4536 16344 4635
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 17972 4604 18000 4644
rect 18509 4641 18521 4675
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 17972 4576 18245 4604
rect 17865 4567 17923 4573
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 15712 4508 16344 4536
rect 17880 4536 17908 4567
rect 18138 4536 18144 4548
rect 17880 4508 18144 4536
rect 15712 4496 15718 4508
rect 18138 4496 18144 4508
rect 18196 4536 18202 4548
rect 18524 4536 18552 4635
rect 18196 4508 18552 4536
rect 18196 4496 18202 4508
rect 16574 4468 16580 4480
rect 13924 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 16666 4428 16672 4480
rect 16724 4428 16730 4480
rect 17034 4428 17040 4480
rect 17092 4468 17098 4480
rect 17221 4471 17279 4477
rect 17221 4468 17233 4471
rect 17092 4440 17233 4468
rect 17092 4428 17098 4440
rect 17221 4437 17233 4440
rect 17267 4437 17279 4471
rect 17221 4431 17279 4437
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 17828 4440 18429 4468
rect 17828 4428 17834 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 19076 4468 19104 4712
rect 19242 4632 19248 4684
rect 19300 4632 19306 4684
rect 19334 4632 19340 4684
rect 19392 4672 19398 4684
rect 19904 4681 19932 4712
rect 20625 4709 20637 4712
rect 20671 4709 20683 4743
rect 21174 4740 21180 4752
rect 20625 4703 20683 4709
rect 20732 4712 21180 4740
rect 20438 4681 20444 4684
rect 19429 4675 19487 4681
rect 19429 4672 19441 4675
rect 19392 4644 19441 4672
rect 19392 4632 19398 4644
rect 19429 4641 19441 4644
rect 19475 4672 19487 4675
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19475 4644 19533 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 20436 4672 20444 4681
rect 20399 4644 20444 4672
rect 19889 4635 19947 4641
rect 20436 4635 20444 4644
rect 20438 4632 20444 4635
rect 20496 4632 20502 4684
rect 20533 4675 20591 4681
rect 20533 4641 20545 4675
rect 20579 4672 20591 4675
rect 20732 4672 20760 4712
rect 21174 4700 21180 4712
rect 21232 4700 21238 4752
rect 21726 4700 21732 4752
rect 21784 4700 21790 4752
rect 20579 4644 20760 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20806 4632 20812 4684
rect 20864 4632 20870 4684
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 21637 4675 21695 4681
rect 20956 4644 21588 4672
rect 20956 4632 20962 4644
rect 19610 4564 19616 4616
rect 19668 4564 19674 4616
rect 19981 4607 20039 4613
rect 19981 4573 19993 4607
rect 20027 4604 20039 4607
rect 20823 4604 20851 4632
rect 21560 4604 21588 4644
rect 21637 4641 21649 4675
rect 21683 4672 21695 4675
rect 21836 4672 21864 4768
rect 21683 4644 21864 4672
rect 21683 4641 21695 4644
rect 21637 4635 21695 4641
rect 20027 4576 20760 4604
rect 20823 4576 21404 4604
rect 21560 4576 21864 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 19150 4496 19156 4548
rect 19208 4536 19214 4548
rect 20257 4539 20315 4545
rect 20257 4536 20269 4539
rect 19208 4508 20269 4536
rect 19208 4496 19214 4508
rect 20257 4505 20269 4508
rect 20303 4505 20315 4539
rect 20257 4499 20315 4505
rect 19337 4471 19395 4477
rect 19337 4468 19349 4471
rect 18840 4440 19349 4468
rect 18840 4428 18846 4440
rect 19337 4437 19349 4440
rect 19383 4437 19395 4471
rect 19337 4431 19395 4437
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 20165 4471 20223 4477
rect 20165 4468 20177 4471
rect 19484 4440 20177 4468
rect 19484 4428 19490 4440
rect 20165 4437 20177 4440
rect 20211 4437 20223 4471
rect 20732 4468 20760 4576
rect 21376 4548 21404 4576
rect 21836 4548 21864 4576
rect 21358 4496 21364 4548
rect 21416 4496 21422 4548
rect 21818 4496 21824 4548
rect 21876 4496 21882 4548
rect 21928 4536 21956 4768
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4672 22155 4675
rect 22278 4672 22284 4684
rect 22143 4644 22284 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22278 4632 22284 4644
rect 22336 4632 22342 4684
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22388 4604 22416 4780
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 23106 4768 23112 4820
rect 23164 4768 23170 4820
rect 23566 4768 23572 4820
rect 23624 4768 23630 4820
rect 24210 4768 24216 4820
rect 24268 4768 24274 4820
rect 24394 4768 24400 4820
rect 24452 4808 24458 4820
rect 25130 4808 25136 4820
rect 24452 4780 25136 4808
rect 24452 4768 24458 4780
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 25774 4808 25780 4820
rect 25608 4780 25780 4808
rect 22554 4700 22560 4752
rect 22612 4740 22618 4752
rect 23124 4740 23152 4768
rect 22612 4712 22968 4740
rect 23124 4712 23336 4740
rect 22612 4700 22618 4712
rect 22940 4684 22968 4712
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4672 22523 4675
rect 22649 4675 22707 4681
rect 22511 4644 22600 4672
rect 22511 4641 22523 4644
rect 22465 4635 22523 4641
rect 22051 4576 22416 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22572 4536 22600 4644
rect 22649 4641 22661 4675
rect 22695 4672 22707 4675
rect 22830 4672 22836 4684
rect 22695 4644 22836 4672
rect 22695 4641 22707 4644
rect 22649 4635 22707 4641
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 22922 4632 22928 4684
rect 22980 4632 22986 4684
rect 23308 4681 23336 4712
rect 23109 4675 23167 4681
rect 23109 4641 23121 4675
rect 23155 4641 23167 4675
rect 23109 4635 23167 4641
rect 23201 4675 23259 4681
rect 23201 4641 23213 4675
rect 23247 4641 23259 4675
rect 23201 4635 23259 4641
rect 23293 4675 23351 4681
rect 23293 4641 23305 4675
rect 23339 4641 23351 4675
rect 23584 4672 23612 4768
rect 25222 4700 25228 4752
rect 25280 4740 25286 4752
rect 25608 4740 25636 4780
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26326 4768 26332 4820
rect 26384 4808 26390 4820
rect 26384 4780 27752 4808
rect 26384 4768 26390 4780
rect 26421 4743 26479 4749
rect 26421 4740 26433 4743
rect 25280 4712 25636 4740
rect 25280 4700 25286 4712
rect 23661 4675 23719 4681
rect 23661 4672 23673 4675
rect 23293 4635 23351 4641
rect 23400 4644 23673 4672
rect 21928 4508 22600 4536
rect 23124 4536 23152 4635
rect 23216 4604 23244 4635
rect 23400 4604 23428 4644
rect 23661 4641 23673 4644
rect 23707 4641 23719 4675
rect 23661 4635 23719 4641
rect 23937 4675 23995 4681
rect 23937 4641 23949 4675
rect 23983 4641 23995 4675
rect 23937 4635 23995 4641
rect 24029 4675 24087 4681
rect 24029 4641 24041 4675
rect 24075 4672 24087 4675
rect 24486 4672 24492 4684
rect 24075 4644 24492 4672
rect 24075 4641 24087 4644
rect 24029 4635 24087 4641
rect 23216 4576 23428 4604
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23952 4604 23980 4635
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 24949 4675 25007 4681
rect 24949 4641 24961 4675
rect 24995 4672 25007 4675
rect 25130 4672 25136 4684
rect 24995 4644 25136 4672
rect 24995 4641 25007 4644
rect 24949 4635 25007 4641
rect 25130 4632 25136 4644
rect 25188 4672 25194 4684
rect 25608 4681 25636 4712
rect 25700 4712 26433 4740
rect 25700 4684 25728 4712
rect 26421 4709 26433 4712
rect 26467 4740 26479 4743
rect 26510 4740 26516 4752
rect 26467 4712 26516 4740
rect 26467 4709 26479 4712
rect 26421 4703 26479 4709
rect 26510 4700 26516 4712
rect 26568 4700 26574 4752
rect 26637 4743 26695 4749
rect 26637 4709 26649 4743
rect 26683 4740 26695 4743
rect 26878 4740 26884 4752
rect 26683 4712 26884 4740
rect 26683 4709 26695 4712
rect 26637 4703 26695 4709
rect 26878 4700 26884 4712
rect 26936 4700 26942 4752
rect 27724 4749 27752 4780
rect 27709 4743 27767 4749
rect 27172 4712 27660 4740
rect 25593 4675 25651 4681
rect 25188 4644 25452 4672
rect 25188 4632 25194 4644
rect 23615 4576 23980 4604
rect 25041 4607 25099 4613
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 25041 4573 25053 4607
rect 25087 4604 25099 4607
rect 25314 4604 25320 4616
rect 25087 4576 25320 4604
rect 25087 4573 25099 4576
rect 25041 4567 25099 4573
rect 25314 4564 25320 4576
rect 25372 4564 25378 4616
rect 25424 4604 25452 4644
rect 25593 4641 25605 4675
rect 25639 4641 25651 4675
rect 25593 4635 25651 4641
rect 25682 4632 25688 4684
rect 25740 4632 25746 4684
rect 25869 4675 25927 4681
rect 25869 4641 25881 4675
rect 25915 4641 25927 4675
rect 25869 4635 25927 4641
rect 25961 4675 26019 4681
rect 25961 4641 25973 4675
rect 26007 4672 26019 4675
rect 26326 4672 26332 4684
rect 26007 4644 26332 4672
rect 26007 4641 26019 4644
rect 25961 4635 26019 4641
rect 25884 4604 25912 4635
rect 26326 4632 26332 4644
rect 26384 4632 26390 4684
rect 26786 4632 26792 4684
rect 26844 4672 26850 4684
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 26844 4644 27077 4672
rect 26844 4632 26850 4644
rect 27065 4641 27077 4644
rect 27111 4641 27123 4675
rect 27065 4635 27123 4641
rect 26804 4604 26832 4632
rect 27172 4613 27200 4712
rect 27525 4675 27583 4681
rect 27525 4672 27537 4675
rect 27264 4644 27537 4672
rect 25424 4576 26832 4604
rect 27157 4607 27215 4613
rect 27157 4573 27169 4607
rect 27203 4573 27215 4607
rect 27157 4567 27215 4573
rect 23198 4536 23204 4548
rect 23124 4508 23204 4536
rect 21928 4468 21956 4508
rect 20732 4440 21956 4468
rect 22572 4468 22600 4508
rect 23198 4496 23204 4508
rect 23256 4496 23262 4548
rect 23308 4508 25544 4536
rect 23308 4468 23336 4508
rect 25516 4480 25544 4508
rect 25590 4496 25596 4548
rect 25648 4536 25654 4548
rect 26326 4536 26332 4548
rect 25648 4508 26332 4536
rect 25648 4496 25654 4508
rect 26326 4496 26332 4508
rect 26384 4496 26390 4548
rect 26510 4496 26516 4548
rect 26568 4536 26574 4548
rect 26789 4539 26847 4545
rect 26789 4536 26801 4539
rect 26568 4508 26801 4536
rect 26568 4496 26574 4508
rect 26789 4505 26801 4508
rect 26835 4536 26847 4539
rect 27264 4536 27292 4644
rect 27525 4641 27537 4644
rect 27571 4641 27583 4675
rect 27632 4672 27660 4712
rect 27709 4709 27721 4743
rect 27755 4709 27767 4743
rect 27709 4703 27767 4709
rect 27893 4743 27951 4749
rect 27893 4709 27905 4743
rect 27939 4709 27951 4743
rect 27893 4703 27951 4709
rect 27908 4672 27936 4703
rect 27632 4644 27936 4672
rect 27525 4635 27583 4641
rect 26835 4508 27292 4536
rect 27433 4539 27491 4545
rect 26835 4505 26847 4508
rect 26789 4499 26847 4505
rect 27433 4505 27445 4539
rect 27479 4536 27491 4539
rect 27522 4536 27528 4548
rect 27479 4508 27528 4536
rect 27479 4505 27491 4508
rect 27433 4499 27491 4505
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 22572 4440 23336 4468
rect 20165 4431 20223 4437
rect 23382 4428 23388 4480
rect 23440 4468 23446 4480
rect 23753 4471 23811 4477
rect 23753 4468 23765 4471
rect 23440 4440 23765 4468
rect 23440 4428 23446 4440
rect 23753 4437 23765 4440
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 23842 4428 23848 4480
rect 23900 4468 23906 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 23900 4440 24685 4468
rect 23900 4428 23906 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 25406 4428 25412 4480
rect 25464 4428 25470 4480
rect 25498 4428 25504 4480
rect 25556 4428 25562 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 26605 4471 26663 4477
rect 26605 4468 26617 4471
rect 26292 4440 26617 4468
rect 26292 4428 26298 4440
rect 26605 4437 26617 4440
rect 26651 4437 26663 4471
rect 26605 4431 26663 4437
rect 26694 4428 26700 4480
rect 26752 4468 26758 4480
rect 26970 4468 26976 4480
rect 26752 4440 26976 4468
rect 26752 4428 26758 4440
rect 26970 4428 26976 4440
rect 27028 4468 27034 4480
rect 29638 4468 29644 4480
rect 27028 4440 29644 4468
rect 27028 4428 27034 4440
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 552 4378 31648 4400
rect 552 4326 4285 4378
rect 4337 4326 4349 4378
rect 4401 4326 4413 4378
rect 4465 4326 4477 4378
rect 4529 4326 4541 4378
rect 4593 4326 12059 4378
rect 12111 4326 12123 4378
rect 12175 4326 12187 4378
rect 12239 4326 12251 4378
rect 12303 4326 12315 4378
rect 12367 4326 19833 4378
rect 19885 4326 19897 4378
rect 19949 4326 19961 4378
rect 20013 4326 20025 4378
rect 20077 4326 20089 4378
rect 20141 4326 27607 4378
rect 27659 4326 27671 4378
rect 27723 4326 27735 4378
rect 27787 4326 27799 4378
rect 27851 4326 27863 4378
rect 27915 4326 31648 4378
rect 552 4304 31648 4326
rect 1029 4267 1087 4273
rect 1029 4233 1041 4267
rect 1075 4264 1087 4267
rect 1118 4264 1124 4276
rect 1075 4236 1124 4264
rect 1075 4233 1087 4236
rect 1029 4227 1087 4233
rect 1118 4224 1124 4236
rect 1176 4224 1182 4276
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 4782 4267 4840 4273
rect 4782 4264 4794 4267
rect 4672 4236 4794 4264
rect 4672 4224 4678 4236
rect 4782 4233 4794 4236
rect 4828 4233 4840 4267
rect 4782 4227 4840 4233
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6730 4264 6736 4276
rect 6319 4236 6736 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7190 4224 7196 4276
rect 7248 4224 7254 4276
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 8205 4267 8263 4273
rect 8205 4233 8217 4267
rect 8251 4264 8263 4267
rect 8846 4264 8852 4276
rect 8251 4236 8852 4264
rect 8251 4233 8263 4236
rect 8205 4227 8263 4233
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9640 4236 9781 4264
rect 9640 4224 9646 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 9769 4227 9827 4233
rect 10410 4224 10416 4276
rect 10468 4224 10474 4276
rect 10873 4267 10931 4273
rect 10873 4233 10885 4267
rect 10919 4264 10931 4267
rect 10962 4264 10968 4276
rect 10919 4236 10968 4264
rect 10919 4233 10931 4236
rect 10873 4227 10931 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14332 4236 14749 4264
rect 14332 4224 14338 4236
rect 14737 4233 14749 4236
rect 14783 4233 14795 4267
rect 14737 4227 14795 4233
rect 15105 4267 15163 4273
rect 15105 4233 15117 4267
rect 15151 4264 15163 4267
rect 15654 4264 15660 4276
rect 15151 4236 15660 4264
rect 15151 4233 15163 4236
rect 15105 4227 15163 4233
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 16022 4224 16028 4276
rect 16080 4264 16086 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 16080 4236 18981 4264
rect 16080 4224 16086 4236
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 18969 4227 19027 4233
rect 19702 4224 19708 4276
rect 19760 4264 19766 4276
rect 19760 4236 22140 4264
rect 19760 4224 19766 4236
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 3878 4196 3884 4208
rect 2832 4168 3884 4196
rect 2832 4156 2838 4168
rect 3878 4156 3884 4168
rect 3936 4156 3942 4208
rect 7208 4196 7236 4224
rect 6196 4168 7236 4196
rect 7484 4196 7512 4224
rect 9306 4196 9312 4208
rect 7484 4168 8800 4196
rect 1026 4088 1032 4140
rect 1084 4088 1090 4140
rect 1121 4131 1179 4137
rect 1121 4097 1133 4131
rect 1167 4128 1179 4131
rect 2038 4128 2044 4140
rect 1167 4100 2044 4128
rect 1167 4097 1179 4100
rect 1121 4091 1179 4097
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3234 4128 3240 4140
rect 2924 4100 3240 4128
rect 2924 4088 2930 4100
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 6086 4128 6092 4140
rect 3835 4100 6092 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 845 4063 903 4069
rect 845 4029 857 4063
rect 891 4060 903 4063
rect 1044 4060 1072 4088
rect 891 4032 1072 4060
rect 891 4029 903 4032
rect 845 4023 903 4029
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 2464 4032 2728 4060
rect 2464 4020 2470 4032
rect 1394 3952 1400 4004
rect 1452 3952 1458 4004
rect 2700 3992 2728 4032
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 3050 4060 3056 4072
rect 2832 4032 3056 4060
rect 2832 4020 2838 4032
rect 3050 4020 3056 4032
rect 3108 4060 3114 4072
rect 3804 4060 3832 4091
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 3108 4032 3832 4060
rect 3108 4020 3114 4032
rect 4062 4020 4068 4072
rect 4120 4020 4126 4072
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 4080 3992 4108 4020
rect 2700 3964 4108 3992
rect 4448 3992 4476 4023
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6196 4060 6224 4168
rect 7558 4128 7564 4140
rect 7024 4100 7564 4128
rect 5960 4032 6224 4060
rect 6457 4063 6515 4069
rect 5960 4020 5966 4032
rect 6457 4029 6469 4063
rect 6503 4060 6515 4063
rect 7024 4060 7052 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7668 4137 7696 4168
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 8570 4128 8576 4140
rect 7653 4091 7711 4097
rect 8036 4100 8576 4128
rect 6503 4032 7052 4060
rect 6503 4029 6515 4032
rect 6457 4023 6515 4029
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 8036 4069 8064 4100
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8772 4137 8800 4168
rect 8956 4168 9312 4196
rect 8956 4137 8984 4168
rect 9306 4156 9312 4168
rect 9364 4156 9370 4208
rect 9401 4199 9459 4205
rect 9401 4165 9413 4199
rect 9447 4196 9459 4199
rect 10428 4196 10456 4224
rect 9447 4168 10456 4196
rect 9447 4165 9459 4168
rect 9401 4159 9459 4165
rect 13998 4156 14004 4208
rect 14056 4196 14062 4208
rect 15010 4196 15016 4208
rect 14056 4168 15016 4196
rect 14056 4156 14062 4168
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 10505 4131 10563 4137
rect 9272 4100 9996 4128
rect 9272 4088 9278 4100
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 7156 4032 7481 4060
rect 7156 4020 7162 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 9968 4060 9996 4100
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 11514 4128 11520 4140
rect 10735 4100 11520 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13596 4100 13645 4128
rect 13596 4088 13602 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 8435 4032 9904 4060
rect 9968 4032 11253 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 4890 3992 4896 4004
rect 4448 3964 4896 3992
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 6178 3952 6184 4004
rect 6236 3992 6242 4004
rect 7009 3995 7067 4001
rect 6236 3964 6408 3992
rect 6236 3952 6242 3964
rect 3234 3884 3240 3936
rect 3292 3884 3298 3936
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3384 3896 3617 3924
rect 3384 3884 3390 3896
rect 3605 3893 3617 3896
rect 3651 3893 3663 3927
rect 3605 3887 3663 3893
rect 3694 3884 3700 3936
rect 3752 3884 3758 3936
rect 4246 3884 4252 3936
rect 4304 3884 4310 3936
rect 6380 3924 6408 3964
rect 7009 3961 7021 3995
rect 7055 3992 7067 3995
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 7055 3964 7573 3992
rect 7055 3961 7067 3964
rect 7009 3955 7067 3961
rect 7561 3961 7573 3964
rect 7607 3961 7619 3995
rect 7561 3955 7619 3961
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 9030 3992 9036 4004
rect 8812 3964 9036 3992
rect 8812 3952 8818 3964
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9766 3952 9772 4004
rect 9824 3952 9830 4004
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 6380 3896 7113 3924
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9548 3896 9597 3924
rect 9548 3884 9554 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9876 3924 9904 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 13004 4060 13032 4088
rect 11379 4032 13032 4060
rect 14093 4063 14151 4069
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14200 4060 14228 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 15473 4199 15531 4205
rect 15473 4165 15485 4199
rect 15519 4196 15531 4199
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 15519 4168 17785 4196
rect 15519 4165 15531 4168
rect 15473 4159 15531 4165
rect 17773 4165 17785 4168
rect 17819 4165 17831 4199
rect 17773 4159 17831 4165
rect 17865 4199 17923 4205
rect 17865 4165 17877 4199
rect 17911 4196 17923 4199
rect 18230 4196 18236 4208
rect 17911 4168 18236 4196
rect 17911 4165 17923 4168
rect 17865 4159 17923 4165
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 20530 4196 20536 4208
rect 19352 4168 20536 4196
rect 16209 4131 16267 4137
rect 14292 4100 15516 4128
rect 14292 4069 14320 4100
rect 14139 4032 14228 4060
rect 14277 4063 14335 4069
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14277 4029 14289 4063
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4060 14427 4063
rect 14415 4032 14504 4060
rect 14415 4029 14427 4032
rect 14369 4023 14427 4029
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10502 3992 10508 4004
rect 9999 3964 10508 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 11256 3992 11284 4023
rect 11256 3964 11468 3992
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 9876 3896 10057 3924
rect 9585 3887 9643 3893
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 10410 3884 10416 3936
rect 10468 3884 10474 3936
rect 11440 3924 11468 3964
rect 11606 3952 11612 4004
rect 11664 3992 11670 4004
rect 13814 3992 13820 4004
rect 11664 3964 13820 3992
rect 11664 3952 11670 3964
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14476 3936 14504 4032
rect 15010 4020 15016 4072
rect 15068 4020 15074 4072
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 15378 4020 15384 4072
rect 15436 4020 15442 4072
rect 15194 3952 15200 4004
rect 15252 3952 15258 4004
rect 13538 3924 13544 3936
rect 11440 3896 13544 3924
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 14458 3884 14464 3936
rect 14516 3884 14522 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15396 3924 15424 4020
rect 15488 3992 15516 4100
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16298 4128 16304 4140
rect 16255 4100 16304 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16666 4128 16672 4140
rect 16531 4100 16672 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16666 4088 16672 4100
rect 16724 4128 16730 4140
rect 16724 4100 19288 4128
rect 16724 4088 16730 4100
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16022 4060 16028 4072
rect 15611 4032 16028 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16960 4069 16988 4100
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 16945 4063 17003 4069
rect 16945 4029 16957 4063
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 16206 3992 16212 4004
rect 15488 3964 16212 3992
rect 16206 3952 16212 3964
rect 16264 3952 16270 4004
rect 16408 3992 16436 4023
rect 16853 3995 16911 4001
rect 16408 3964 16712 3992
rect 16684 3936 16712 3964
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 17144 3992 17172 4023
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 17770 4060 17776 4072
rect 17368 4032 17776 4060
rect 17368 4020 17374 4032
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 18782 4060 18788 4072
rect 17972 4032 18788 4060
rect 17972 3992 18000 4032
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 19150 4020 19156 4072
rect 19208 4020 19214 4072
rect 19260 4069 19288 4100
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 16899 3964 18000 3992
rect 18049 3995 18107 4001
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 18049 3961 18061 3995
rect 18095 3992 18107 3995
rect 19352 3992 19380 4168
rect 20530 4156 20536 4168
rect 20588 4156 20594 4208
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 19668 4100 20208 4128
rect 19668 4088 19674 4100
rect 19426 4020 19432 4072
rect 19484 4020 19490 4072
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 19702 4060 19708 4072
rect 19567 4032 19708 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 19536 3992 19564 4023
rect 19702 4020 19708 4032
rect 19760 4020 19766 4072
rect 20070 4020 20076 4072
rect 20128 4020 20134 4072
rect 20180 4069 20208 4100
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20254 4060 20260 4072
rect 20211 4032 20260 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20346 4020 20352 4072
rect 20404 4020 20410 4072
rect 20438 4020 20444 4072
rect 20496 4020 20502 4072
rect 20640 4060 20668 4236
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4097 21971 4131
rect 21913 4091 21971 4097
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 20640 4032 20821 4060
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 20902 4063 20960 4069
rect 20902 4029 20914 4063
rect 20948 4029 20960 4063
rect 20902 4023 20960 4029
rect 18095 3964 19380 3992
rect 19444 3964 19564 3992
rect 20272 3992 20300 4020
rect 20917 3992 20945 4023
rect 21174 4020 21180 4072
rect 21232 4020 21238 4072
rect 21266 4020 21272 4072
rect 21324 4069 21330 4072
rect 21324 4060 21332 4069
rect 21729 4063 21787 4069
rect 21324 4032 21369 4060
rect 21324 4023 21332 4032
rect 21729 4029 21741 4063
rect 21775 4060 21787 4063
rect 21818 4060 21824 4072
rect 21775 4032 21824 4060
rect 21775 4029 21787 4032
rect 21729 4023 21787 4029
rect 21324 4020 21330 4023
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 21928 4060 21956 4091
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22112 4128 22140 4236
rect 22922 4224 22928 4276
rect 22980 4264 22986 4276
rect 22980 4236 24072 4264
rect 22980 4224 22986 4236
rect 22462 4196 22468 4208
rect 22388 4168 22468 4196
rect 22388 4137 22416 4168
rect 22462 4156 22468 4168
rect 22520 4196 22526 4208
rect 23198 4196 23204 4208
rect 22520 4168 23204 4196
rect 22520 4156 22526 4168
rect 23198 4156 23204 4168
rect 23256 4156 23262 4208
rect 23474 4156 23480 4208
rect 23532 4156 23538 4208
rect 24044 4196 24072 4236
rect 24118 4224 24124 4276
rect 24176 4224 24182 4276
rect 25866 4224 25872 4276
rect 25924 4224 25930 4276
rect 26237 4267 26295 4273
rect 26237 4233 26249 4267
rect 26283 4264 26295 4267
rect 26283 4236 28120 4264
rect 26283 4233 26295 4236
rect 26237 4227 26295 4233
rect 24670 4196 24676 4208
rect 24044 4168 24676 4196
rect 22373 4131 22431 4137
rect 22112 4100 22324 4128
rect 21928 4032 22048 4060
rect 20272 3964 20945 3992
rect 21085 3995 21143 4001
rect 18095 3961 18107 3964
rect 18049 3955 18107 3961
rect 19444 3936 19472 3964
rect 21085 3961 21097 3995
rect 21131 3992 21143 3995
rect 21131 3964 21864 3992
rect 21131 3961 21143 3964
rect 21085 3955 21143 3961
rect 15160 3896 15424 3924
rect 15160 3884 15166 3896
rect 16666 3884 16672 3936
rect 16724 3884 16730 3936
rect 17037 3927 17095 3933
rect 17037 3893 17049 3927
rect 17083 3924 17095 3927
rect 17126 3924 17132 3936
rect 17083 3896 17132 3924
rect 17083 3893 17095 3896
rect 17037 3887 17095 3893
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 19426 3884 19432 3936
rect 19484 3884 19490 3936
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 19889 3927 19947 3933
rect 19889 3924 19901 3927
rect 19760 3896 19901 3924
rect 19760 3884 19766 3896
rect 19889 3893 19901 3896
rect 19935 3893 19947 3927
rect 19889 3887 19947 3893
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 21100 3924 21128 3955
rect 21836 3936 21864 3964
rect 20312 3896 21128 3924
rect 20312 3884 20318 3896
rect 21450 3884 21456 3936
rect 21508 3884 21514 3936
rect 21542 3884 21548 3936
rect 21600 3884 21606 3936
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 22020 3924 22048 4032
rect 22296 3936 22324 4100
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 22741 4131 22799 4137
rect 22741 4097 22753 4131
rect 22787 4128 22799 4131
rect 24121 4131 24179 4137
rect 24121 4128 24133 4131
rect 22787 4100 24133 4128
rect 22787 4097 22799 4100
rect 22741 4091 22799 4097
rect 24121 4097 24133 4100
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 22557 4063 22615 4069
rect 22557 4029 22569 4063
rect 22603 4060 22615 4063
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22603 4032 23029 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 23017 4029 23029 4032
rect 23063 4060 23075 4063
rect 23201 4063 23259 4069
rect 23063 4032 23152 4060
rect 23063 4029 23075 4032
rect 23017 4023 23075 4029
rect 21876 3896 22048 3924
rect 21876 3884 21882 3896
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 23014 3924 23020 3936
rect 22336 3896 23020 3924
rect 22336 3884 22342 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23124 3924 23152 4032
rect 23201 4029 23213 4063
rect 23247 4060 23259 4063
rect 23290 4060 23296 4072
rect 23247 4032 23296 4060
rect 23247 4029 23259 4032
rect 23201 4023 23259 4029
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24412 4069 24440 4168
rect 24670 4156 24676 4168
rect 24728 4156 24734 4208
rect 26329 4199 26387 4205
rect 26329 4196 26341 4199
rect 26160 4168 26341 4196
rect 24949 4131 25007 4137
rect 24949 4097 24961 4131
rect 24995 4128 25007 4131
rect 25314 4128 25320 4140
rect 24995 4100 25320 4128
rect 24995 4097 25007 4100
rect 24949 4091 25007 4097
rect 25314 4088 25320 4100
rect 25372 4088 25378 4140
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4029 23535 4063
rect 23477 4023 23535 4029
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4060 23719 4063
rect 24397 4063 24455 4069
rect 23707 4032 24348 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 23492 3992 23520 4023
rect 24320 3992 24348 4032
rect 24397 4029 24409 4063
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24854 4020 24860 4072
rect 24912 4020 24918 4072
rect 25041 4063 25099 4069
rect 25041 4029 25053 4063
rect 25087 4060 25099 4063
rect 25130 4060 25136 4072
rect 25087 4032 25136 4060
rect 25087 4029 25099 4032
rect 25041 4023 25099 4029
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25498 4020 25504 4072
rect 25556 4020 25562 4072
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 25777 4063 25835 4069
rect 25777 4029 25789 4063
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 26053 4063 26111 4069
rect 26053 4029 26065 4063
rect 26099 4060 26111 4063
rect 26160 4060 26188 4168
rect 26329 4165 26341 4168
rect 26375 4165 26387 4199
rect 26329 4159 26387 4165
rect 27617 4199 27675 4205
rect 27617 4165 27629 4199
rect 27663 4196 27675 4199
rect 27985 4199 28043 4205
rect 27985 4196 27997 4199
rect 27663 4168 27997 4196
rect 27663 4165 27675 4168
rect 27617 4159 27675 4165
rect 27985 4165 27997 4168
rect 28031 4165 28043 4199
rect 27985 4159 28043 4165
rect 26418 4088 26424 4140
rect 26476 4128 26482 4140
rect 28092 4137 28120 4236
rect 28077 4131 28135 4137
rect 26476 4100 27844 4128
rect 26476 4088 26482 4100
rect 26510 4069 26516 4072
rect 26508 4060 26516 4069
rect 26099 4032 26188 4060
rect 26436 4032 26516 4060
rect 26099 4029 26111 4032
rect 26053 4023 26111 4029
rect 24872 3992 24900 4020
rect 23492 3964 23888 3992
rect 24320 3964 24900 3992
rect 23566 3924 23572 3936
rect 23124 3896 23572 3924
rect 23566 3884 23572 3896
rect 23624 3924 23630 3936
rect 23750 3924 23756 3936
rect 23624 3896 23756 3924
rect 23624 3884 23630 3896
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 23860 3933 23888 3964
rect 25590 3952 25596 4004
rect 25648 3952 25654 4004
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 24762 3884 24768 3936
rect 24820 3884 24826 3936
rect 25409 3927 25467 3933
rect 25409 3893 25421 3927
rect 25455 3924 25467 3927
rect 25700 3924 25728 4023
rect 25792 3992 25820 4023
rect 26436 3992 26464 4032
rect 26508 4023 26516 4032
rect 26510 4020 26516 4023
rect 26568 4020 26574 4072
rect 26620 4069 26648 4100
rect 26605 4063 26663 4069
rect 26605 4029 26617 4063
rect 26651 4029 26663 4063
rect 26878 4060 26884 4072
rect 26839 4032 26884 4060
rect 26605 4023 26663 4029
rect 26878 4020 26884 4032
rect 26936 4020 26942 4072
rect 26970 4020 26976 4072
rect 27028 4020 27034 4072
rect 27062 4020 27068 4072
rect 27120 4020 27126 4072
rect 27154 4020 27160 4072
rect 27212 4020 27218 4072
rect 27246 4020 27252 4072
rect 27304 4060 27310 4072
rect 27341 4063 27399 4069
rect 27341 4060 27353 4063
rect 27304 4032 27353 4060
rect 27304 4020 27310 4032
rect 27341 4029 27353 4032
rect 27387 4029 27399 4063
rect 27341 4023 27399 4029
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 25792 3964 26464 3992
rect 26694 3952 26700 4004
rect 26752 3952 26758 4004
rect 27448 3992 27476 4023
rect 26896 3964 27476 3992
rect 26712 3924 26740 3952
rect 26896 3936 26924 3964
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 27709 3995 27767 4001
rect 27709 3992 27721 3995
rect 27580 3964 27721 3992
rect 27580 3952 27586 3964
rect 27709 3961 27721 3964
rect 27755 3961 27767 3995
rect 27816 3992 27844 4100
rect 28077 4097 28089 4131
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 27893 4063 27951 4069
rect 27893 4029 27905 4063
rect 27939 4060 27951 4063
rect 27982 4060 27988 4072
rect 27939 4032 27988 4060
rect 27939 4029 27951 4032
rect 27893 4023 27951 4029
rect 27982 4020 27988 4032
rect 28040 4020 28046 4072
rect 28074 3992 28080 4004
rect 27816 3964 28080 3992
rect 27709 3955 27767 3961
rect 28074 3952 28080 3964
rect 28132 3952 28138 4004
rect 28166 3952 28172 4004
rect 28224 3952 28230 4004
rect 25455 3896 26740 3924
rect 25455 3893 25467 3896
rect 25409 3887 25467 3893
rect 26878 3884 26884 3936
rect 26936 3884 26942 3936
rect 552 3834 31808 3856
rect 552 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 15946 3834
rect 15998 3782 16010 3834
rect 16062 3782 16074 3834
rect 16126 3782 16138 3834
rect 16190 3782 16202 3834
rect 16254 3782 23720 3834
rect 23772 3782 23784 3834
rect 23836 3782 23848 3834
rect 23900 3782 23912 3834
rect 23964 3782 23976 3834
rect 24028 3782 31494 3834
rect 31546 3782 31558 3834
rect 31610 3782 31622 3834
rect 31674 3782 31686 3834
rect 31738 3782 31750 3834
rect 31802 3782 31808 3834
rect 552 3760 31808 3782
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 4522 3720 4528 3732
rect 2096 3692 4528 3720
rect 2096 3680 2102 3692
rect 4522 3680 4528 3692
rect 4580 3720 4586 3732
rect 4798 3720 4804 3732
rect 4580 3692 4804 3720
rect 4580 3680 4586 3692
rect 4798 3680 4804 3692
rect 4856 3720 4862 3732
rect 6822 3720 6828 3732
rect 4856 3692 6316 3720
rect 4856 3680 4862 3692
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 2056 3593 2084 3680
rect 4062 3652 4068 3664
rect 3542 3624 4068 3652
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 4157 3655 4215 3661
rect 4157 3621 4169 3655
rect 4203 3652 4215 3655
rect 4246 3652 4252 3664
rect 4203 3624 4252 3652
rect 4203 3621 4215 3624
rect 4157 3615 4215 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 5902 3652 5908 3664
rect 5382 3624 5908 3652
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 6178 3612 6184 3664
rect 6236 3612 6242 3664
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 3878 3544 3884 3596
rect 3936 3544 3942 3596
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 6196 3584 6224 3612
rect 6043 3556 6224 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 6288 3525 6316 3692
rect 6564 3692 6828 3720
rect 6564 3661 6592 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 9214 3720 9220 3732
rect 8496 3692 9220 3720
rect 8496 3664 8524 3692
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9364 3692 9965 3720
rect 9364 3680 9370 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 7006 3612 7012 3664
rect 7064 3612 7070 3664
rect 8386 3612 8392 3664
rect 8444 3612 8450 3664
rect 8478 3612 8484 3664
rect 8536 3612 8542 3664
rect 9122 3612 9128 3664
rect 9180 3612 9186 3664
rect 11256 3652 11284 3683
rect 11422 3680 11428 3732
rect 11480 3720 11486 3732
rect 11974 3720 11980 3732
rect 11480 3692 11980 3720
rect 11480 3680 11486 3692
rect 11974 3680 11980 3692
rect 12032 3720 12038 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12032 3692 13093 3720
rect 12032 3680 12038 3692
rect 13081 3689 13093 3692
rect 13127 3720 13139 3723
rect 14826 3720 14832 3732
rect 13127 3692 14832 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 14826 3680 14832 3692
rect 14884 3680 14890 3732
rect 14921 3723 14979 3729
rect 14921 3689 14933 3723
rect 14967 3720 14979 3723
rect 15194 3720 15200 3732
rect 14967 3692 15200 3720
rect 14967 3689 14979 3692
rect 14921 3683 14979 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 15344 3692 16221 3720
rect 15344 3680 15350 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 18138 3680 18144 3732
rect 18196 3680 18202 3732
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 20254 3720 20260 3732
rect 19116 3692 20260 3720
rect 19116 3680 19122 3692
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20404 3692 20913 3720
rect 20404 3680 20410 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 20990 3680 20996 3732
rect 21048 3680 21054 3732
rect 21450 3680 21456 3732
rect 21508 3680 21514 3732
rect 21726 3720 21732 3732
rect 21652 3692 21732 3720
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11256 3624 11621 3652
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 12618 3612 12624 3664
rect 12676 3612 12682 3664
rect 13814 3612 13820 3664
rect 13872 3612 13878 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 15304 3652 15332 3680
rect 21008 3652 21036 3680
rect 21468 3652 21496 3680
rect 21652 3661 21680 3692
rect 21726 3680 21732 3692
rect 21784 3680 21790 3732
rect 21818 3680 21824 3732
rect 21876 3680 21882 3732
rect 22002 3680 22008 3732
rect 22060 3720 22066 3732
rect 22060 3692 22324 3720
rect 22060 3680 22066 3692
rect 14056 3624 14320 3652
rect 14056 3612 14062 3624
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 9646 3556 10517 3584
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3516 6331 3519
rect 8018 3516 8024 3528
rect 6319 3488 8024 3516
rect 6319 3485 6331 3488
rect 6273 3479 6331 3485
rect 8018 3476 8024 3488
rect 8076 3516 8082 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 8076 3488 8125 3516
rect 8076 3476 8082 3488
rect 8113 3485 8125 3488
rect 8159 3516 8171 3519
rect 8846 3516 8852 3528
rect 8159 3488 8852 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9646 3516 9674 3556
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11146 3584 11152 3596
rect 11103 3556 11152 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 14292 3593 14320 3624
rect 15212 3624 15332 3652
rect 17420 3624 18276 3652
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11296 3556 11345 3584
rect 11296 3544 11302 3556
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11333 3547 11391 3553
rect 14277 3587 14335 3593
rect 14277 3553 14289 3587
rect 14323 3553 14335 3587
rect 14277 3547 14335 3553
rect 14458 3544 14464 3596
rect 14516 3544 14522 3596
rect 9456 3488 9674 3516
rect 9861 3519 9919 3525
rect 9456 3476 9462 3488
rect 9861 3485 9873 3519
rect 9907 3516 9919 3519
rect 9950 3516 9956 3528
rect 9907 3488 9956 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10410 3476 10416 3528
rect 10468 3476 10474 3528
rect 11606 3516 11612 3528
rect 11440 3488 11612 3516
rect 1394 3408 1400 3460
rect 1452 3448 1458 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 1452 3420 1501 3448
rect 1452 3408 1458 3420
rect 1489 3417 1501 3420
rect 1535 3417 1547 3451
rect 10428 3448 10456 3476
rect 11440 3448 11468 3488
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 10428 3420 11468 3448
rect 14476 3448 14504 3544
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 15212 3525 15240 3624
rect 17420 3596 17448 3624
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15378 3584 15384 3596
rect 15335 3556 15384 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3584 16635 3587
rect 17313 3587 17371 3593
rect 16623 3556 17172 3584
rect 16623 3553 16635 3556
rect 16577 3547 16635 3553
rect 17144 3528 17172 3556
rect 17313 3553 17325 3587
rect 17359 3584 17371 3587
rect 17402 3584 17408 3596
rect 17359 3556 17408 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17497 3587 17555 3593
rect 17497 3553 17509 3587
rect 17543 3584 17555 3587
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17543 3556 17601 3584
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 17589 3547 17647 3553
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3584 17831 3587
rect 17862 3584 17868 3596
rect 17819 3556 17868 3584
rect 17819 3553 17831 3556
rect 17773 3547 17831 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18248 3593 18276 3624
rect 18708 3624 19840 3652
rect 18708 3593 18736 3624
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3553 18567 3587
rect 18509 3547 18567 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 19058 3584 19064 3596
rect 18693 3547 18751 3553
rect 18800 3556 19064 3584
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 14476 3420 15516 3448
rect 1489 3411 1547 3417
rect 15488 3392 15516 3420
rect 16684 3392 16712 3479
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 18064 3516 18092 3547
rect 17184 3488 18092 3516
rect 18524 3516 18552 3547
rect 18800 3516 18828 3556
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 19812 3593 19840 3624
rect 20824 3624 21036 3652
rect 21284 3624 21496 3652
rect 21637 3655 21695 3661
rect 19797 3587 19855 3593
rect 19797 3553 19809 3587
rect 19843 3584 19855 3587
rect 20162 3584 20168 3596
rect 19843 3556 20168 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 20824 3593 20852 3624
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20312 3556 20821 3584
rect 20312 3544 20318 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 20990 3544 20996 3596
rect 21048 3544 21054 3596
rect 21284 3593 21312 3624
rect 21637 3621 21649 3655
rect 21683 3621 21695 3655
rect 21836 3652 21864 3680
rect 21836 3624 22232 3652
rect 21637 3615 21695 3621
rect 21450 3593 21456 3596
rect 21269 3587 21327 3593
rect 21269 3553 21281 3587
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 21417 3587 21456 3593
rect 21417 3553 21429 3587
rect 21417 3547 21456 3553
rect 21450 3544 21456 3547
rect 21508 3544 21514 3596
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3553 21603 3587
rect 21734 3587 21792 3593
rect 21734 3584 21746 3587
rect 21545 3547 21603 3553
rect 21652 3556 21746 3584
rect 18524 3488 18828 3516
rect 20717 3519 20775 3525
rect 17184 3476 17190 3488
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 20898 3516 20904 3528
rect 20763 3488 20904 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 20898 3476 20904 3488
rect 20956 3516 20962 3528
rect 21560 3516 21588 3547
rect 20956 3488 21588 3516
rect 20956 3476 20962 3488
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 18325 3451 18383 3457
rect 18325 3448 18337 3451
rect 17552 3420 18337 3448
rect 17552 3408 17558 3420
rect 18325 3417 18337 3420
rect 18371 3417 18383 3451
rect 18325 3411 18383 3417
rect 19610 3408 19616 3460
rect 19668 3448 19674 3460
rect 20070 3448 20076 3460
rect 19668 3420 20076 3448
rect 19668 3408 19674 3420
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 21652 3448 21680 3556
rect 21734 3553 21746 3556
rect 21780 3584 21792 3587
rect 21910 3584 21916 3596
rect 21780 3556 21916 3584
rect 21780 3553 21792 3556
rect 21734 3547 21792 3553
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22204 3593 22232 3624
rect 22296 3593 22324 3692
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 23842 3720 23848 3732
rect 23256 3692 23848 3720
rect 23256 3680 23262 3692
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24029 3723 24087 3729
rect 24029 3689 24041 3723
rect 24075 3720 24087 3723
rect 26050 3720 26056 3732
rect 24075 3692 26056 3720
rect 24075 3689 24087 3692
rect 24029 3683 24087 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 26694 3720 26700 3732
rect 26283 3692 26700 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 26694 3680 26700 3692
rect 26752 3680 26758 3732
rect 28166 3680 28172 3732
rect 28224 3680 28230 3732
rect 24394 3612 24400 3664
rect 24452 3612 24458 3664
rect 24854 3612 24860 3664
rect 24912 3652 24918 3664
rect 28184 3652 28212 3680
rect 24912 3624 28212 3652
rect 24912 3612 24918 3624
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22281 3587 22339 3593
rect 22281 3553 22293 3587
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 22922 3544 22928 3596
rect 22980 3584 22986 3596
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 22980 3556 23489 3584
rect 22980 3544 22986 3556
rect 23477 3553 23489 3556
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 23937 3587 23995 3593
rect 23937 3553 23949 3587
rect 23983 3584 23995 3587
rect 24026 3584 24032 3596
rect 23983 3556 24032 3584
rect 23983 3553 23995 3556
rect 23937 3547 23995 3553
rect 24026 3544 24032 3556
rect 24084 3544 24090 3596
rect 24213 3587 24271 3593
rect 24213 3553 24225 3587
rect 24259 3584 24271 3587
rect 24259 3556 24624 3584
rect 24259 3553 24271 3556
rect 24213 3547 24271 3553
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 21876 3488 21956 3516
rect 21876 3476 21882 3488
rect 21928 3457 21956 3488
rect 23290 3476 23296 3528
rect 23348 3476 23354 3528
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 20824 3420 21680 3448
rect 21913 3451 21971 3457
rect 20824 3392 20852 3420
rect 21913 3417 21925 3451
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6638 3380 6644 3392
rect 6227 3352 6644 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3380 8079 3383
rect 8754 3380 8760 3392
rect 8067 3352 8760 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 11422 3380 11428 3392
rect 9088 3352 11428 3380
rect 9088 3340 9094 3352
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 16666 3340 16672 3392
rect 16724 3340 16730 3392
rect 16850 3340 16856 3392
rect 16908 3380 16914 3392
rect 20530 3380 20536 3392
rect 16908 3352 20536 3380
rect 16908 3340 16914 3352
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 20806 3340 20812 3392
rect 20864 3340 20870 3392
rect 23106 3340 23112 3392
rect 23164 3340 23170 3392
rect 23400 3380 23428 3479
rect 23584 3448 23612 3479
rect 23658 3476 23664 3528
rect 23716 3516 23722 3528
rect 24305 3519 24363 3525
rect 24305 3516 24317 3519
rect 23716 3488 24317 3516
rect 23716 3476 23722 3488
rect 24305 3485 24317 3488
rect 24351 3485 24363 3519
rect 24596 3516 24624 3556
rect 24670 3544 24676 3596
rect 24728 3544 24734 3596
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3584 24823 3587
rect 25130 3584 25136 3596
rect 24811 3556 25136 3584
rect 24811 3553 24823 3556
rect 24765 3547 24823 3553
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 25682 3544 25688 3596
rect 25740 3544 25746 3596
rect 25866 3544 25872 3596
rect 25924 3584 25930 3596
rect 26053 3587 26111 3593
rect 26053 3584 26065 3587
rect 25924 3556 26065 3584
rect 25924 3544 25930 3556
rect 26053 3553 26065 3556
rect 26099 3553 26111 3587
rect 26053 3547 26111 3553
rect 26237 3587 26295 3593
rect 26237 3553 26249 3587
rect 26283 3584 26295 3587
rect 26510 3584 26516 3596
rect 26283 3556 26516 3584
rect 26283 3553 26295 3556
rect 26237 3547 26295 3553
rect 25700 3516 25728 3544
rect 24596 3488 25728 3516
rect 24305 3479 24363 3485
rect 25682 3448 25688 3460
rect 23584 3420 25688 3448
rect 25682 3408 25688 3420
rect 25740 3408 25746 3460
rect 26068 3448 26096 3547
rect 26510 3544 26516 3556
rect 26568 3584 26574 3596
rect 27430 3584 27436 3596
rect 26568 3556 27436 3584
rect 26568 3544 26574 3556
rect 27430 3544 27436 3556
rect 27488 3544 27494 3596
rect 27801 3587 27859 3593
rect 27801 3553 27813 3587
rect 27847 3584 27859 3587
rect 27847 3556 28028 3584
rect 27847 3553 27859 3556
rect 27801 3547 27859 3553
rect 26697 3519 26755 3525
rect 26697 3485 26709 3519
rect 26743 3516 26755 3519
rect 26786 3516 26792 3528
rect 26743 3488 26792 3516
rect 26743 3485 26755 3488
rect 26697 3479 26755 3485
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 27154 3476 27160 3528
rect 27212 3516 27218 3528
rect 27525 3519 27583 3525
rect 27525 3516 27537 3519
rect 27212 3488 27537 3516
rect 27212 3476 27218 3488
rect 27525 3485 27537 3488
rect 27571 3516 27583 3519
rect 27893 3519 27951 3525
rect 27893 3516 27905 3519
rect 27571 3488 27905 3516
rect 27571 3485 27583 3488
rect 27525 3479 27583 3485
rect 27893 3485 27905 3488
rect 27939 3485 27951 3519
rect 27893 3479 27951 3485
rect 26878 3448 26884 3460
rect 26068 3420 26884 3448
rect 26878 3408 26884 3420
rect 26936 3448 26942 3460
rect 28000 3448 28028 3556
rect 26936 3420 28028 3448
rect 26936 3408 26942 3420
rect 23566 3380 23572 3392
rect 23400 3352 23572 3380
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 24213 3383 24271 3389
rect 24213 3349 24225 3383
rect 24259 3380 24271 3383
rect 24486 3380 24492 3392
rect 24259 3352 24492 3380
rect 24259 3349 24271 3352
rect 24213 3343 24271 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 24946 3340 24952 3392
rect 25004 3340 25010 3392
rect 552 3290 31648 3312
rect 552 3238 4285 3290
rect 4337 3238 4349 3290
rect 4401 3238 4413 3290
rect 4465 3238 4477 3290
rect 4529 3238 4541 3290
rect 4593 3238 12059 3290
rect 12111 3238 12123 3290
rect 12175 3238 12187 3290
rect 12239 3238 12251 3290
rect 12303 3238 12315 3290
rect 12367 3238 19833 3290
rect 19885 3238 19897 3290
rect 19949 3238 19961 3290
rect 20013 3238 20025 3290
rect 20077 3238 20089 3290
rect 20141 3238 27607 3290
rect 27659 3238 27671 3290
rect 27723 3238 27735 3290
rect 27787 3238 27799 3290
rect 27851 3238 27863 3290
rect 27915 3238 31648 3290
rect 552 3216 31648 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1728 3148 1869 3176
rect 1728 3136 1734 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 1857 3139 1915 3145
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2777 3179 2835 3185
rect 2777 3176 2789 3179
rect 2372 3148 2789 3176
rect 2372 3136 2378 3148
rect 2777 3145 2789 3148
rect 2823 3145 2835 3179
rect 2777 3139 2835 3145
rect 3234 3136 3240 3188
rect 3292 3136 3298 3188
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3752 3148 3801 3176
rect 3752 3136 3758 3148
rect 3789 3145 3801 3148
rect 3835 3145 3847 3179
rect 3789 3139 3847 3145
rect 5810 3136 5816 3188
rect 5868 3136 5874 3188
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7892 3148 8033 3176
rect 7892 3136 7898 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8444 3148 8493 3176
rect 8444 3136 8450 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 8481 3139 8539 3145
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8628 3148 9996 3176
rect 8628 3136 8634 3148
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 2884 2972 2912 3000
rect 2363 2944 2912 2972
rect 2961 2975 3019 2981
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3252 2972 3280 3136
rect 8757 3111 8815 3117
rect 6840 3080 8064 3108
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 3844 3012 4353 3040
rect 3844 3000 3850 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3040 6515 3043
rect 6730 3040 6736 3052
rect 6503 3012 6736 3040
rect 6503 3009 6515 3012
rect 6457 3003 6515 3009
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 3007 2944 3280 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2498 2904 2504 2916
rect 2271 2876 2504 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2498 2864 2504 2876
rect 2556 2904 2562 2916
rect 6840 2904 6868 3080
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7742 3040 7748 3052
rect 7699 3012 7748 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 6963 2944 7052 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 2556 2876 6868 2904
rect 2556 2864 2562 2876
rect 7024 2845 7052 2944
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 7156 2944 7389 2972
rect 7156 2932 7162 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 7392 2904 7420 2935
rect 7669 2904 7697 3003
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8036 3040 8064 3080
rect 8757 3077 8769 3111
rect 8803 3077 8815 3111
rect 8757 3071 8815 3077
rect 8478 3040 8484 3052
rect 8036 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7984 2944 8217 2972
rect 7984 2932 7990 2944
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 8772 2972 8800 3071
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 8904 3080 9904 3108
rect 8904 3068 8910 3080
rect 9876 3049 9904 3080
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 8711 2944 8800 2972
rect 8864 3012 9321 3040
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 8864 2904 8892 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9968 3040 9996 3148
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11701 3179 11759 3185
rect 11701 3176 11713 3179
rect 11204 3148 11713 3176
rect 11204 3136 11210 3148
rect 11701 3145 11713 3148
rect 11747 3145 11759 3179
rect 11701 3139 11759 3145
rect 14918 3136 14924 3188
rect 14976 3136 14982 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15378 3176 15384 3188
rect 15335 3148 15384 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15470 3136 15476 3188
rect 15528 3136 15534 3188
rect 16666 3136 16672 3188
rect 16724 3136 16730 3188
rect 16850 3176 16856 3188
rect 16776 3148 16856 3176
rect 11422 3068 11428 3120
rect 11480 3068 11486 3120
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 11848 3080 13584 3108
rect 11848 3068 11854 3080
rect 10137 3043 10195 3049
rect 10137 3040 10149 3043
rect 9968 3012 10149 3040
rect 9861 3003 9919 3009
rect 10137 3009 10149 3012
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 9088 2944 9137 2972
rect 9088 2932 9094 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10410 2904 10416 2916
rect 7392 2876 7604 2904
rect 7669 2876 8892 2904
rect 9140 2876 10416 2904
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 7466 2796 7472 2848
rect 7524 2796 7530 2848
rect 7576 2836 7604 2876
rect 9140 2836 9168 2876
rect 10410 2864 10416 2876
rect 10468 2864 10474 2916
rect 11440 2904 11468 3068
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 13556 3049 13584 3080
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11572 3012 12265 3040
rect 11572 3000 11578 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14277 3043 14335 3049
rect 14277 3040 14289 3043
rect 13964 3012 14289 3040
rect 13964 3000 13970 3012
rect 14277 3009 14289 3012
rect 14323 3009 14335 3043
rect 14277 3003 14335 3009
rect 15286 3000 15292 3052
rect 15344 3000 15350 3052
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15620 3012 15945 3040
rect 15620 3000 15626 3012
rect 15933 3009 15945 3012
rect 15979 3040 15991 3043
rect 16776 3040 16804 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17494 3136 17500 3188
rect 17552 3136 17558 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 18656 3148 18889 3176
rect 18656 3136 18662 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 19797 3179 19855 3185
rect 19797 3145 19809 3179
rect 19843 3176 19855 3179
rect 19843 3148 20392 3176
rect 19843 3145 19855 3148
rect 19797 3139 19855 3145
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 15979 3012 16804 3040
rect 16868 3080 19993 3108
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 12032 2944 12173 2972
rect 12032 2932 12038 2944
rect 12161 2941 12173 2944
rect 12207 2941 12219 2975
rect 12161 2935 12219 2941
rect 13998 2932 14004 2984
rect 14056 2932 14062 2984
rect 14182 2932 14188 2984
rect 14240 2932 14246 2984
rect 15304 2972 15332 3000
rect 15381 2975 15439 2981
rect 15381 2972 15393 2975
rect 15304 2944 15393 2972
rect 15381 2941 15393 2944
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 15654 2932 15660 2984
rect 15712 2932 15718 2984
rect 15838 2932 15844 2984
rect 15896 2932 15902 2984
rect 16758 2932 16764 2984
rect 16816 2932 16822 2984
rect 16868 2981 16896 3080
rect 19981 3077 19993 3080
rect 20027 3077 20039 3111
rect 20364 3108 20392 3148
rect 20438 3136 20444 3188
rect 20496 3136 20502 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 22094 3176 22100 3188
rect 20588 3148 22100 3176
rect 20588 3136 20594 3148
rect 22094 3136 22100 3148
rect 22152 3176 22158 3188
rect 23014 3176 23020 3188
rect 22152 3148 23020 3176
rect 22152 3136 22158 3148
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 23106 3136 23112 3188
rect 23164 3136 23170 3188
rect 23290 3136 23296 3188
rect 23348 3136 23354 3188
rect 24029 3179 24087 3185
rect 24029 3176 24041 3179
rect 23492 3148 24041 3176
rect 20714 3108 20720 3120
rect 20364 3080 20720 3108
rect 19981 3071 20039 3077
rect 19610 3040 19616 3052
rect 16960 3012 19616 3040
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 10520 2876 10626 2904
rect 11440 2876 12081 2904
rect 7576 2808 9168 2836
rect 9214 2796 9220 2848
rect 9272 2796 9278 2848
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10520 2836 10548 2876
rect 12069 2873 12081 2876
rect 12115 2904 12127 2907
rect 13538 2904 13544 2916
rect 12115 2876 13544 2904
rect 12115 2873 12127 2876
rect 12069 2867 12127 2873
rect 13538 2864 13544 2876
rect 13596 2904 13602 2916
rect 16390 2904 16396 2916
rect 13596 2876 16396 2904
rect 13596 2864 13602 2876
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 16776 2904 16804 2932
rect 16960 2904 16988 3012
rect 17126 2932 17132 2984
rect 17184 2932 17190 2984
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17236 2904 17264 2935
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17972 2981 18000 3012
rect 19610 3000 19616 3012
rect 19668 3000 19674 3052
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19760 3012 19901 3040
rect 19760 3000 19766 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19996 3040 20024 3071
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 21818 3068 21824 3120
rect 21876 3068 21882 3120
rect 23124 3108 23152 3136
rect 22940 3080 23152 3108
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 19996 3012 21005 3040
rect 19889 3003 19947 3009
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 21726 3040 21732 3052
rect 20993 3003 21051 3009
rect 21468 3012 21732 3040
rect 17773 2975 17831 2981
rect 17773 2972 17785 2975
rect 17460 2944 17785 2972
rect 17460 2932 17466 2944
rect 17773 2941 17785 2944
rect 17819 2941 17831 2975
rect 17773 2935 17831 2941
rect 17957 2975 18015 2981
rect 17957 2941 17969 2975
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 19426 2975 19484 2981
rect 19426 2972 19438 2975
rect 18187 2944 19438 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 19426 2941 19438 2944
rect 19472 2972 19484 2975
rect 19794 2972 19800 2984
rect 19472 2944 19800 2972
rect 19472 2941 19484 2944
rect 19426 2935 19484 2941
rect 16776 2876 16988 2904
rect 17052 2876 17264 2904
rect 10376 2808 10548 2836
rect 10376 2796 10382 2808
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 10836 2808 11621 2836
rect 10836 2796 10842 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 17052 2845 17080 2876
rect 17586 2864 17592 2916
rect 17644 2904 17650 2916
rect 18156 2904 18184 2935
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 19978 2932 19984 2984
rect 20036 2932 20042 2984
rect 20165 2975 20223 2981
rect 20165 2941 20177 2975
rect 20211 2972 20223 2975
rect 20254 2972 20260 2984
rect 20211 2944 20260 2972
rect 20211 2941 20223 2944
rect 20165 2935 20223 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20901 2975 20959 2981
rect 20901 2941 20913 2975
rect 20947 2972 20959 2975
rect 21468 2972 21496 3012
rect 21726 3000 21732 3012
rect 21784 3000 21790 3052
rect 20947 2944 21496 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 21542 2932 21548 2984
rect 21600 2972 21606 2984
rect 21836 2981 21864 3068
rect 22940 2981 22968 3080
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 21600 2944 21649 2972
rect 21600 2932 21606 2944
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 21637 2935 21695 2941
rect 21821 2975 21879 2981
rect 21821 2941 21833 2975
rect 21867 2941 21879 2975
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 21821 2935 21879 2941
rect 21928 2944 22661 2972
rect 17644 2876 18184 2904
rect 17644 2864 17650 2876
rect 18414 2864 18420 2916
rect 18472 2904 18478 2916
rect 18690 2904 18696 2916
rect 18472 2876 18696 2904
rect 18472 2864 18478 2876
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 21266 2904 21272 2916
rect 20855 2876 21272 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 21928 2904 21956 2944
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 22833 2975 22891 2981
rect 22833 2941 22845 2975
rect 22879 2941 22891 2975
rect 22833 2935 22891 2941
rect 22925 2975 22983 2981
rect 22925 2941 22937 2975
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 21376 2876 21956 2904
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16632 2808 17049 2836
rect 16632 2796 16638 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17678 2796 17684 2848
rect 17736 2796 17742 2848
rect 18874 2796 18880 2848
rect 18932 2845 18938 2848
rect 18932 2839 18951 2845
rect 18939 2805 18951 2839
rect 18932 2799 18951 2805
rect 18932 2796 18938 2799
rect 19058 2796 19064 2848
rect 19116 2796 19122 2848
rect 19245 2839 19303 2845
rect 19245 2805 19257 2839
rect 19291 2836 19303 2839
rect 19334 2836 19340 2848
rect 19291 2808 19340 2836
rect 19291 2805 19303 2808
rect 19245 2799 19303 2805
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19429 2839 19487 2845
rect 19429 2805 19441 2839
rect 19475 2836 19487 2839
rect 19978 2836 19984 2848
rect 19475 2808 19984 2836
rect 19475 2805 19487 2808
rect 19429 2799 19487 2805
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 21376 2836 21404 2876
rect 22094 2864 22100 2916
rect 22152 2904 22158 2916
rect 22189 2907 22247 2913
rect 22189 2904 22201 2907
rect 22152 2876 22201 2904
rect 22152 2864 22158 2876
rect 22189 2873 22201 2876
rect 22235 2873 22247 2907
rect 22189 2867 22247 2873
rect 22370 2864 22376 2916
rect 22428 2864 22434 2916
rect 20128 2808 21404 2836
rect 20128 2796 20134 2808
rect 21450 2796 21456 2848
rect 21508 2796 21514 2848
rect 22002 2796 22008 2848
rect 22060 2796 22066 2848
rect 22848 2836 22876 2935
rect 23124 2904 23152 3003
rect 23198 2932 23204 2984
rect 23256 2972 23262 2984
rect 23382 2972 23388 2984
rect 23256 2944 23388 2972
rect 23256 2932 23262 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23492 2981 23520 3148
rect 24029 3145 24041 3148
rect 24075 3176 24087 3179
rect 24118 3176 24124 3188
rect 24075 3148 24124 3176
rect 24075 3145 24087 3148
rect 24029 3139 24087 3145
rect 24118 3136 24124 3148
rect 24176 3136 24182 3188
rect 24854 3136 24860 3188
rect 24912 3136 24918 3188
rect 24946 3136 24952 3188
rect 25004 3176 25010 3188
rect 25004 3148 25268 3176
rect 25004 3136 25010 3148
rect 23750 3068 23756 3120
rect 23808 3068 23814 3120
rect 23768 3040 23796 3068
rect 23768 3012 24072 3040
rect 23477 2975 23535 2981
rect 23477 2941 23489 2975
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 23842 2932 23848 2984
rect 23900 2932 23906 2984
rect 24044 2981 24072 3012
rect 24136 2981 24164 3136
rect 24872 3108 24900 3136
rect 24596 3080 24900 3108
rect 25041 3111 25099 3117
rect 24210 3000 24216 3052
rect 24268 3040 24274 3052
rect 24268 3012 24348 3040
rect 24268 3000 24274 3012
rect 24320 2981 24348 3012
rect 24596 2981 24624 3080
rect 25041 3077 25053 3111
rect 25087 3077 25099 3111
rect 25041 3071 25099 3077
rect 24670 3000 24676 3052
rect 24728 3000 24734 3052
rect 24029 2975 24087 2981
rect 24029 2941 24041 2975
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 24121 2975 24179 2981
rect 24121 2941 24133 2975
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24305 2975 24363 2981
rect 24305 2941 24317 2975
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 24545 2975 24624 2981
rect 24545 2941 24557 2975
rect 24591 2944 24624 2975
rect 24688 2972 24716 3000
rect 24946 2981 24952 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24688 2944 24777 2972
rect 24591 2941 24603 2944
rect 24545 2935 24603 2941
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 24765 2935 24823 2941
rect 24903 2975 24952 2981
rect 24903 2941 24915 2975
rect 24949 2941 24952 2975
rect 24903 2935 24952 2941
rect 23661 2907 23719 2913
rect 23661 2904 23673 2907
rect 23124 2876 23673 2904
rect 23661 2873 23673 2876
rect 23707 2904 23719 2907
rect 23934 2904 23940 2916
rect 23707 2876 23940 2904
rect 23707 2873 23719 2876
rect 23661 2867 23719 2873
rect 23934 2864 23940 2876
rect 23992 2864 23998 2916
rect 24210 2904 24216 2916
rect 24044 2876 24216 2904
rect 24044 2836 24072 2876
rect 24210 2864 24216 2876
rect 24268 2864 24274 2916
rect 22848 2808 24072 2836
rect 24118 2796 24124 2848
rect 24176 2796 24182 2848
rect 24412 2836 24440 2935
rect 24946 2932 24952 2935
rect 25004 2932 25010 2984
rect 25056 2972 25084 3071
rect 25240 2981 25268 3148
rect 25682 3136 25688 3188
rect 25740 3136 25746 3188
rect 26789 3179 26847 3185
rect 26789 3145 26801 3179
rect 26835 3176 26847 3179
rect 27154 3176 27160 3188
rect 26835 3148 27160 3176
rect 26835 3145 26847 3148
rect 26789 3139 26847 3145
rect 27154 3136 27160 3148
rect 27212 3136 27218 3188
rect 26970 3108 26976 3120
rect 25424 3080 26976 3108
rect 25424 2981 25452 3080
rect 26970 3068 26976 3080
rect 27028 3068 27034 3120
rect 27065 3043 27123 3049
rect 26620 3012 27016 3040
rect 25133 2975 25191 2981
rect 25133 2972 25145 2975
rect 25056 2944 25145 2972
rect 25133 2941 25145 2944
rect 25179 2941 25191 2975
rect 25133 2935 25191 2941
rect 25225 2975 25283 2981
rect 25225 2941 25237 2975
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 25409 2975 25467 2981
rect 25409 2941 25421 2975
rect 25455 2941 25467 2975
rect 25409 2935 25467 2941
rect 25501 2975 25559 2981
rect 25501 2941 25513 2975
rect 25547 2941 25559 2975
rect 25501 2935 25559 2941
rect 24670 2864 24676 2916
rect 24728 2864 24734 2916
rect 25038 2864 25044 2916
rect 25096 2864 25102 2916
rect 25314 2864 25320 2916
rect 25372 2904 25378 2916
rect 25516 2904 25544 2935
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 26620 2981 26648 3012
rect 26988 2981 27016 3012
rect 27065 3009 27077 3043
rect 27111 3040 27123 3043
rect 27430 3040 27436 3052
rect 27111 3012 27436 3040
rect 27111 3009 27123 3012
rect 27065 3003 27123 3009
rect 26605 2975 26663 2981
rect 26605 2972 26617 2975
rect 25648 2944 26617 2972
rect 25648 2932 25654 2944
rect 26605 2941 26617 2944
rect 26651 2941 26663 2975
rect 26605 2935 26663 2941
rect 26881 2975 26939 2981
rect 26881 2941 26893 2975
rect 26927 2941 26939 2975
rect 26881 2935 26939 2941
rect 26973 2975 27031 2981
rect 26973 2941 26985 2975
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 25372 2876 25544 2904
rect 26896 2904 26924 2935
rect 27080 2904 27108 3003
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 26896 2876 27108 2904
rect 25372 2864 25378 2876
rect 25056 2836 25084 2864
rect 24412 2808 25084 2836
rect 26418 2796 26424 2848
rect 26476 2796 26482 2848
rect 27338 2796 27344 2848
rect 27396 2796 27402 2848
rect 552 2746 31808 2768
rect 552 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 15946 2746
rect 15998 2694 16010 2746
rect 16062 2694 16074 2746
rect 16126 2694 16138 2746
rect 16190 2694 16202 2746
rect 16254 2694 23720 2746
rect 23772 2694 23784 2746
rect 23836 2694 23848 2746
rect 23900 2694 23912 2746
rect 23964 2694 23976 2746
rect 24028 2694 31494 2746
rect 31546 2694 31558 2746
rect 31610 2694 31622 2746
rect 31674 2694 31686 2746
rect 31738 2694 31750 2746
rect 31802 2694 31808 2746
rect 552 2672 31808 2694
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 7524 2604 7757 2632
rect 7524 2592 7530 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 7745 2595 7803 2601
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9272 2604 9597 2632
rect 9272 2592 9278 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 15654 2632 15660 2644
rect 15611 2604 15660 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 17310 2592 17316 2644
rect 17368 2592 17374 2644
rect 17586 2592 17592 2644
rect 17644 2592 17650 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17736 2604 17816 2632
rect 17736 2592 17742 2604
rect 13538 2524 13544 2576
rect 13596 2524 13602 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 15396 2536 15761 2564
rect 15396 2508 15424 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15749 2527 15807 2533
rect 15838 2524 15844 2576
rect 15896 2524 15902 2576
rect 17604 2564 17632 2592
rect 16960 2536 17632 2564
rect 17788 2564 17816 2604
rect 18230 2592 18236 2644
rect 18288 2592 18294 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 18874 2632 18880 2644
rect 18564 2604 18880 2632
rect 18564 2592 18570 2604
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 21358 2632 21364 2644
rect 18984 2604 21364 2632
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 17788 2536 18797 2564
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8662 2496 8668 2508
rect 8435 2468 8668 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9732 2468 10149 2496
rect 9732 2456 9738 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 13998 2456 14004 2508
rect 14056 2456 14062 2508
rect 14182 2456 14188 2508
rect 14240 2456 14246 2508
rect 14274 2456 14280 2508
rect 14332 2456 14338 2508
rect 15194 2456 15200 2508
rect 15252 2456 15258 2508
rect 15378 2456 15384 2508
rect 15436 2456 15442 2508
rect 15657 2499 15715 2505
rect 15657 2465 15669 2499
rect 15703 2465 15715 2499
rect 15856 2495 15884 2524
rect 15657 2459 15715 2465
rect 15841 2489 15899 2495
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15120 2360 15148 2391
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 15672 2428 15700 2459
rect 15841 2455 15853 2489
rect 15887 2455 15899 2489
rect 16666 2456 16672 2508
rect 16724 2456 16730 2508
rect 16960 2505 16988 2536
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 18984 2564 19012 2604
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 21910 2632 21916 2644
rect 21468 2604 21916 2632
rect 20898 2564 20904 2576
rect 18785 2527 18843 2533
rect 18908 2536 19012 2564
rect 19536 2536 20904 2564
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 17589 2499 17647 2505
rect 17589 2465 17601 2499
rect 17635 2496 17647 2499
rect 17678 2496 17684 2508
rect 17635 2468 17684 2496
rect 17635 2465 17647 2468
rect 17589 2459 17647 2465
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 17954 2496 17960 2508
rect 17788 2468 17960 2496
rect 15841 2449 15899 2455
rect 15746 2428 15752 2440
rect 15672 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16209 2431 16267 2437
rect 16209 2397 16221 2431
rect 16255 2428 16267 2431
rect 16574 2428 16580 2440
rect 16255 2400 16580 2428
rect 16255 2397 16267 2400
rect 16209 2391 16267 2397
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2428 17371 2431
rect 17788 2428 17816 2468
rect 17954 2456 17960 2468
rect 18012 2496 18018 2508
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 18012 2468 18429 2496
rect 18012 2456 18018 2468
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 18506 2456 18512 2508
rect 18564 2456 18570 2508
rect 18598 2456 18604 2508
rect 18656 2456 18662 2508
rect 18908 2496 18936 2536
rect 18800 2468 18936 2496
rect 17359 2400 17816 2428
rect 17865 2431 17923 2437
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 17865 2397 17877 2431
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 18524 2428 18552 2456
rect 18095 2400 18552 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 17880 2360 17908 2391
rect 18138 2360 18144 2372
rect 15120 2332 17080 2360
rect 17880 2332 18144 2360
rect 17052 2292 17080 2332
rect 18138 2320 18144 2332
rect 18196 2360 18202 2372
rect 18616 2360 18644 2456
rect 18800 2440 18828 2468
rect 19058 2456 19064 2508
rect 19116 2456 19122 2508
rect 19153 2499 19211 2505
rect 19153 2465 19165 2499
rect 19199 2496 19211 2499
rect 19242 2496 19248 2508
rect 19199 2468 19248 2496
rect 19199 2465 19211 2468
rect 19153 2459 19211 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19334 2456 19340 2508
rect 19392 2456 19398 2508
rect 19426 2456 19432 2508
rect 19484 2456 19490 2508
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 19536 2428 19564 2536
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 21468 2564 21496 2604
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 22370 2592 22376 2644
rect 22428 2632 22434 2644
rect 22649 2635 22707 2641
rect 22649 2632 22661 2635
rect 22428 2604 22661 2632
rect 22428 2592 22434 2604
rect 22649 2601 22661 2604
rect 22695 2601 22707 2635
rect 22649 2595 22707 2601
rect 23293 2635 23351 2641
rect 23293 2601 23305 2635
rect 23339 2632 23351 2635
rect 23382 2632 23388 2644
rect 23339 2604 23388 2632
rect 23339 2601 23351 2604
rect 23293 2595 23351 2601
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 23952 2604 24992 2632
rect 21100 2536 21496 2564
rect 19610 2456 19616 2508
rect 19668 2494 19674 2508
rect 19797 2499 19855 2505
rect 19797 2494 19809 2499
rect 19668 2466 19809 2494
rect 19668 2456 19674 2466
rect 19797 2465 19809 2466
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 19978 2456 19984 2508
rect 20036 2456 20042 2508
rect 20806 2456 20812 2508
rect 20864 2456 20870 2508
rect 20990 2456 20996 2508
rect 21048 2456 21054 2508
rect 21100 2505 21128 2536
rect 21542 2524 21548 2576
rect 21600 2524 21606 2576
rect 23477 2567 23535 2573
rect 23477 2564 23489 2567
rect 22112 2536 23489 2564
rect 21085 2499 21143 2505
rect 21085 2465 21097 2499
rect 21131 2465 21143 2499
rect 21085 2459 21143 2465
rect 21266 2456 21272 2508
rect 21324 2456 21330 2508
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21560 2468 21741 2496
rect 19024 2400 19564 2428
rect 19705 2431 19763 2437
rect 19024 2388 19030 2400
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 19996 2428 20024 2456
rect 19751 2400 20024 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 21008 2428 21036 2456
rect 21450 2428 21456 2440
rect 20404 2400 21456 2428
rect 20404 2388 20410 2400
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 18196 2332 18644 2360
rect 18196 2320 18202 2332
rect 19794 2320 19800 2372
rect 19852 2360 19858 2372
rect 21560 2369 21588 2468
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 22002 2456 22008 2508
rect 22060 2456 22066 2508
rect 22112 2372 22140 2536
rect 23477 2533 23489 2536
rect 23523 2533 23535 2567
rect 23477 2527 23535 2533
rect 22186 2456 22192 2508
rect 22244 2456 22250 2508
rect 22373 2499 22431 2505
rect 22373 2465 22385 2499
rect 22419 2465 22431 2499
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22373 2459 22431 2465
rect 22848 2468 23397 2496
rect 22388 2428 22416 2459
rect 22848 2437 22876 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 23385 2459 23443 2465
rect 23566 2456 23572 2508
rect 23624 2456 23630 2508
rect 23952 2505 23980 2604
rect 24964 2576 24992 2604
rect 25406 2592 25412 2644
rect 25464 2632 25470 2644
rect 26145 2635 26203 2641
rect 26145 2632 26157 2635
rect 25464 2604 26157 2632
rect 25464 2592 25470 2604
rect 26145 2601 26157 2604
rect 26191 2601 26203 2635
rect 26602 2632 26608 2644
rect 26145 2595 26203 2601
rect 26252 2604 26608 2632
rect 24762 2564 24768 2576
rect 24228 2536 24768 2564
rect 24228 2505 24256 2536
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 24946 2524 24952 2576
rect 25004 2564 25010 2576
rect 25593 2567 25651 2573
rect 25593 2564 25605 2567
rect 25004 2536 25605 2564
rect 25004 2524 25010 2536
rect 25593 2533 25605 2536
rect 25639 2533 25651 2567
rect 25593 2527 25651 2533
rect 23937 2499 23995 2505
rect 23937 2465 23949 2499
rect 23983 2465 23995 2499
rect 23937 2459 23995 2465
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2465 24179 2499
rect 24121 2459 24179 2465
rect 24213 2499 24271 2505
rect 24213 2465 24225 2499
rect 24259 2465 24271 2499
rect 24213 2459 24271 2465
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22388 2400 22845 2428
rect 20625 2363 20683 2369
rect 20625 2360 20637 2363
rect 19852 2332 20637 2360
rect 19852 2320 19858 2332
rect 20625 2329 20637 2332
rect 20671 2329 20683 2363
rect 20625 2323 20683 2329
rect 21545 2363 21603 2369
rect 21545 2329 21557 2363
rect 21591 2329 21603 2363
rect 22094 2360 22100 2372
rect 21545 2323 21603 2329
rect 21652 2332 22100 2360
rect 18877 2295 18935 2301
rect 18877 2292 18889 2295
rect 17052 2264 18889 2292
rect 18877 2261 18889 2264
rect 18923 2261 18935 2295
rect 18877 2255 18935 2261
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 21652 2292 21680 2332
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 19024 2264 21680 2292
rect 21729 2295 21787 2301
rect 19024 2252 19030 2264
rect 21729 2261 21741 2295
rect 21775 2292 21787 2295
rect 21818 2292 21824 2304
rect 21775 2264 21824 2292
rect 21775 2261 21787 2264
rect 21729 2255 21787 2261
rect 21818 2252 21824 2264
rect 21876 2252 21882 2304
rect 22278 2252 22284 2304
rect 22336 2292 22342 2304
rect 22388 2292 22416 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23584 2428 23612 2456
rect 24026 2428 24032 2440
rect 22971 2400 24032 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24136 2428 24164 2459
rect 24302 2456 24308 2508
rect 24360 2496 24366 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 24360 2468 24409 2496
rect 24360 2456 24366 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 24578 2456 24584 2508
rect 24636 2456 24642 2508
rect 25222 2496 25228 2508
rect 24688 2468 25228 2496
rect 24688 2428 24716 2468
rect 25222 2456 25228 2468
rect 25280 2456 25286 2508
rect 25498 2456 25504 2508
rect 25556 2456 25562 2508
rect 25682 2456 25688 2508
rect 25740 2456 25746 2508
rect 25958 2456 25964 2508
rect 26016 2456 26022 2508
rect 26160 2440 26188 2595
rect 26252 2505 26280 2604
rect 26602 2592 26608 2604
rect 26660 2632 26666 2644
rect 27065 2635 27123 2641
rect 27065 2632 27077 2635
rect 26660 2604 27077 2632
rect 26660 2592 26666 2604
rect 27065 2601 27077 2604
rect 27111 2601 27123 2635
rect 27065 2595 27123 2601
rect 27525 2567 27583 2573
rect 27525 2564 27537 2567
rect 26436 2536 27537 2564
rect 26436 2508 26464 2536
rect 27525 2533 27537 2536
rect 27571 2533 27583 2567
rect 27525 2527 27583 2533
rect 26237 2499 26295 2505
rect 26237 2465 26249 2499
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 26418 2456 26424 2508
rect 26476 2456 26482 2508
rect 26789 2499 26847 2505
rect 26789 2465 26801 2499
rect 26835 2465 26847 2499
rect 26789 2459 26847 2465
rect 24136 2400 24716 2428
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25317 2431 25375 2437
rect 25317 2428 25329 2431
rect 24820 2400 25329 2428
rect 24820 2388 24826 2400
rect 25317 2397 25329 2400
rect 25363 2428 25375 2431
rect 25590 2428 25596 2440
rect 25363 2400 25596 2428
rect 25363 2397 25375 2400
rect 25317 2391 25375 2397
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 26142 2388 26148 2440
rect 26200 2428 26206 2440
rect 26804 2428 26832 2459
rect 26200 2400 26832 2428
rect 26973 2431 27031 2437
rect 26200 2388 26206 2400
rect 26973 2397 26985 2431
rect 27019 2428 27031 2431
rect 27019 2400 27292 2428
rect 27019 2397 27031 2400
rect 26973 2391 27031 2397
rect 23474 2320 23480 2372
rect 23532 2360 23538 2372
rect 23532 2332 24164 2360
rect 23532 2320 23538 2332
rect 22336 2264 22416 2292
rect 22336 2252 22342 2264
rect 23750 2252 23756 2304
rect 23808 2252 23814 2304
rect 24136 2292 24164 2332
rect 24210 2320 24216 2372
rect 24268 2360 24274 2372
rect 25961 2363 26019 2369
rect 25961 2360 25973 2363
rect 24268 2332 25973 2360
rect 24268 2320 24274 2332
rect 25961 2329 25973 2332
rect 26007 2329 26019 2363
rect 25961 2323 26019 2329
rect 26510 2320 26516 2372
rect 26568 2320 26574 2372
rect 27264 2369 27292 2400
rect 27249 2363 27307 2369
rect 27249 2329 27261 2363
rect 27295 2360 27307 2363
rect 27338 2360 27344 2372
rect 27295 2332 27344 2360
rect 27295 2329 27307 2332
rect 27249 2323 27307 2329
rect 27338 2320 27344 2332
rect 27396 2320 27402 2372
rect 24302 2292 24308 2304
rect 24136 2264 24308 2292
rect 24302 2252 24308 2264
rect 24360 2292 24366 2304
rect 24670 2292 24676 2304
rect 24360 2264 24676 2292
rect 24360 2252 24366 2264
rect 24670 2252 24676 2264
rect 24728 2252 24734 2304
rect 552 2202 31648 2224
rect 552 2150 4285 2202
rect 4337 2150 4349 2202
rect 4401 2150 4413 2202
rect 4465 2150 4477 2202
rect 4529 2150 4541 2202
rect 4593 2150 12059 2202
rect 12111 2150 12123 2202
rect 12175 2150 12187 2202
rect 12239 2150 12251 2202
rect 12303 2150 12315 2202
rect 12367 2150 19833 2202
rect 19885 2150 19897 2202
rect 19949 2150 19961 2202
rect 20013 2150 20025 2202
rect 20077 2150 20089 2202
rect 20141 2150 27607 2202
rect 27659 2150 27671 2202
rect 27723 2150 27735 2202
rect 27787 2150 27799 2202
rect 27851 2150 27863 2202
rect 27915 2150 31648 2202
rect 552 2128 31648 2150
rect 14553 2091 14611 2097
rect 14553 2057 14565 2091
rect 14599 2088 14611 2091
rect 15286 2088 15292 2100
rect 14599 2060 15292 2088
rect 14599 2057 14611 2060
rect 14553 2051 14611 2057
rect 15286 2048 15292 2060
rect 15344 2048 15350 2100
rect 15838 2048 15844 2100
rect 15896 2048 15902 2100
rect 17126 2088 17132 2100
rect 17052 2060 17132 2088
rect 15105 2023 15163 2029
rect 15105 1989 15117 2023
rect 15151 2020 15163 2023
rect 15856 2020 15884 2048
rect 15151 1992 15884 2020
rect 15151 1989 15163 1992
rect 15105 1983 15163 1989
rect 14921 1887 14979 1893
rect 14921 1853 14933 1887
rect 14967 1884 14979 1887
rect 15120 1884 15148 1983
rect 15565 1955 15623 1961
rect 15565 1921 15577 1955
rect 15611 1952 15623 1955
rect 17052 1952 17080 2060
rect 17126 2048 17132 2060
rect 17184 2088 17190 2100
rect 17184 2060 17632 2088
rect 17184 2048 17190 2060
rect 17494 2020 17500 2032
rect 17144 1992 17500 2020
rect 17144 1961 17172 1992
rect 17494 1980 17500 1992
rect 17552 1980 17558 2032
rect 17604 2020 17632 2060
rect 18138 2048 18144 2100
rect 18196 2048 18202 2100
rect 18874 2048 18880 2100
rect 18932 2048 18938 2100
rect 19334 2048 19340 2100
rect 19392 2088 19398 2100
rect 19392 2060 20852 2088
rect 19392 2048 19398 2060
rect 19610 2020 19616 2032
rect 17604 1992 19616 2020
rect 19610 1980 19616 1992
rect 19668 1980 19674 2032
rect 19981 2023 20039 2029
rect 19981 1989 19993 2023
rect 20027 2020 20039 2023
rect 20027 1992 20760 2020
rect 20027 1989 20039 1992
rect 19981 1983 20039 1989
rect 15611 1924 17080 1952
rect 17129 1955 17187 1961
rect 15611 1921 15623 1924
rect 15565 1915 15623 1921
rect 17129 1921 17141 1955
rect 17175 1921 17187 1955
rect 17129 1915 17187 1921
rect 17405 1955 17463 1961
rect 17405 1921 17417 1955
rect 17451 1921 17463 1955
rect 19058 1952 19064 1964
rect 17405 1915 17463 1921
rect 18248 1924 19064 1952
rect 14967 1856 15148 1884
rect 15473 1887 15531 1893
rect 14967 1853 14979 1856
rect 14921 1847 14979 1853
rect 15473 1853 15485 1887
rect 15519 1884 15531 1887
rect 16574 1884 16580 1896
rect 15519 1856 16580 1884
rect 15519 1853 15531 1856
rect 15473 1847 15531 1853
rect 16574 1844 16580 1856
rect 16632 1884 16638 1896
rect 17037 1887 17095 1893
rect 17037 1884 17049 1887
rect 16632 1856 17049 1884
rect 16632 1844 16638 1856
rect 17037 1853 17049 1856
rect 17083 1853 17095 1887
rect 17037 1847 17095 1853
rect 14737 1819 14795 1825
rect 14737 1785 14749 1819
rect 14783 1816 14795 1819
rect 17420 1816 17448 1915
rect 18248 1816 18276 1924
rect 19058 1912 19064 1924
rect 19116 1952 19122 1964
rect 19153 1955 19211 1961
rect 19153 1952 19165 1955
rect 19116 1924 19165 1952
rect 19116 1912 19122 1924
rect 19153 1921 19165 1924
rect 19199 1921 19211 1955
rect 19996 1952 20024 1983
rect 20732 1961 20760 1992
rect 19153 1915 19211 1921
rect 19444 1924 20024 1952
rect 20441 1955 20499 1961
rect 19444 1893 19472 1924
rect 20441 1921 20453 1955
rect 20487 1921 20499 1955
rect 20441 1915 20499 1921
rect 20717 1955 20775 1961
rect 20717 1921 20729 1955
rect 20763 1921 20775 1955
rect 20717 1915 20775 1921
rect 18325 1887 18383 1893
rect 18325 1853 18337 1887
rect 18371 1884 18383 1887
rect 19429 1887 19487 1893
rect 18371 1856 19012 1884
rect 18371 1853 18383 1856
rect 18325 1847 18383 1853
rect 18509 1819 18567 1825
rect 18509 1816 18521 1819
rect 14783 1788 15792 1816
rect 17420 1788 18521 1816
rect 14783 1785 14795 1788
rect 14737 1779 14795 1785
rect 15764 1760 15792 1788
rect 18509 1785 18521 1788
rect 18555 1785 18567 1819
rect 18984 1816 19012 1856
rect 19429 1853 19441 1887
rect 19475 1853 19487 1887
rect 19429 1847 19487 1853
rect 19527 1887 19585 1893
rect 19527 1853 19539 1887
rect 19573 1884 19585 1887
rect 19573 1856 19656 1884
rect 19573 1853 19585 1856
rect 19527 1847 19585 1853
rect 19628 1816 19656 1856
rect 19702 1844 19708 1896
rect 19760 1884 19766 1896
rect 20346 1884 20352 1896
rect 19760 1856 20352 1884
rect 19760 1844 19766 1856
rect 20346 1844 20352 1856
rect 20404 1844 20410 1896
rect 20456 1828 20484 1915
rect 20824 1896 20852 2060
rect 20898 2048 20904 2100
rect 20956 2048 20962 2100
rect 21085 2091 21143 2097
rect 21085 2057 21097 2091
rect 21131 2088 21143 2091
rect 21266 2088 21272 2100
rect 21131 2060 21272 2088
rect 21131 2057 21143 2060
rect 21085 2051 21143 2057
rect 21266 2048 21272 2060
rect 21324 2048 21330 2100
rect 22278 2048 22284 2100
rect 22336 2048 22342 2100
rect 23750 2048 23756 2100
rect 23808 2048 23814 2100
rect 24394 2048 24400 2100
rect 24452 2048 24458 2100
rect 24578 2088 24584 2100
rect 24504 2060 24584 2088
rect 20916 2020 20944 2048
rect 23474 2020 23480 2032
rect 20916 1992 23480 2020
rect 20806 1844 20812 1896
rect 20864 1844 20870 1896
rect 20916 1884 20944 1992
rect 23474 1980 23480 1992
rect 23532 1980 23538 2032
rect 21910 1952 21916 1964
rect 21871 1924 21916 1952
rect 21910 1912 21916 1924
rect 21968 1952 21974 1964
rect 23768 1952 23796 2048
rect 24504 2020 24532 2060
rect 24578 2048 24584 2060
rect 24636 2088 24642 2100
rect 25133 2091 25191 2097
rect 24636 2060 24992 2088
rect 24636 2048 24642 2060
rect 21968 1924 23796 1952
rect 24412 1992 24532 2020
rect 24964 2020 24992 2060
rect 25133 2057 25145 2091
rect 25179 2088 25191 2091
rect 25314 2088 25320 2100
rect 25179 2060 25320 2088
rect 25179 2057 25191 2060
rect 25133 2051 25191 2057
rect 25314 2048 25320 2060
rect 25372 2048 25378 2100
rect 25409 2091 25467 2097
rect 25409 2057 25421 2091
rect 25455 2088 25467 2091
rect 25498 2088 25504 2100
rect 25455 2060 25504 2088
rect 25455 2057 25467 2060
rect 25409 2051 25467 2057
rect 25498 2048 25504 2060
rect 25556 2088 25562 2100
rect 25556 2060 25820 2088
rect 25556 2048 25562 2060
rect 25682 2020 25688 2032
rect 24964 1992 25688 2020
rect 21968 1912 21974 1924
rect 21269 1887 21327 1893
rect 21269 1884 21281 1887
rect 20916 1856 21281 1884
rect 21269 1853 21281 1856
rect 21315 1853 21327 1887
rect 21269 1847 21327 1853
rect 21453 1887 21511 1893
rect 21453 1853 21465 1887
rect 21499 1853 21511 1887
rect 21453 1847 21511 1853
rect 20438 1816 20444 1828
rect 18984 1788 19196 1816
rect 19628 1788 20444 1816
rect 18509 1779 18567 1785
rect 19168 1760 19196 1788
rect 20438 1776 20444 1788
rect 20496 1816 20502 1828
rect 21361 1819 21419 1825
rect 21361 1816 21373 1819
rect 20496 1788 21373 1816
rect 20496 1776 20502 1788
rect 21361 1785 21373 1788
rect 21407 1785 21419 1819
rect 21468 1816 21496 1847
rect 21542 1844 21548 1896
rect 21600 1884 21606 1896
rect 22005 1887 22063 1893
rect 22005 1884 22017 1887
rect 21600 1856 22017 1884
rect 21600 1844 21606 1856
rect 22005 1853 22017 1856
rect 22051 1853 22063 1887
rect 22005 1847 22063 1853
rect 21726 1816 21732 1828
rect 21468 1788 21732 1816
rect 21361 1779 21419 1785
rect 21726 1776 21732 1788
rect 21784 1816 21790 1828
rect 24412 1816 24440 1992
rect 24854 1912 24860 1964
rect 24912 1912 24918 1964
rect 24765 1887 24823 1893
rect 24765 1886 24777 1887
rect 24811 1886 24823 1887
rect 24762 1834 24768 1886
rect 24820 1834 24826 1886
rect 24964 1884 24992 1992
rect 25682 1980 25688 1992
rect 25740 1980 25746 2032
rect 25792 1952 25820 2060
rect 25958 2048 25964 2100
rect 26016 2088 26022 2100
rect 26513 2091 26571 2097
rect 26513 2088 26525 2091
rect 26016 2060 26525 2088
rect 26016 2048 26022 2060
rect 26513 2057 26525 2060
rect 26559 2057 26571 2091
rect 26513 2051 26571 2057
rect 26602 2048 26608 2100
rect 26660 2048 26666 2100
rect 26142 1980 26148 2032
rect 26200 1980 26206 2032
rect 25240 1924 25820 1952
rect 25240 1893 25268 1924
rect 25041 1887 25099 1893
rect 25041 1884 25053 1887
rect 24964 1856 25053 1884
rect 25041 1853 25053 1856
rect 25087 1853 25099 1887
rect 25041 1847 25099 1853
rect 25225 1887 25283 1893
rect 25225 1853 25237 1887
rect 25271 1853 25283 1887
rect 25225 1847 25283 1853
rect 25317 1887 25375 1893
rect 25317 1853 25329 1887
rect 25363 1853 25375 1887
rect 26160 1884 26188 1980
rect 26234 1912 26240 1964
rect 26292 1952 26298 1964
rect 26421 1955 26479 1961
rect 26421 1952 26433 1955
rect 26292 1924 26433 1952
rect 26292 1912 26298 1924
rect 26421 1921 26433 1924
rect 26467 1952 26479 1955
rect 27982 1952 27988 1964
rect 26467 1924 27988 1952
rect 26467 1921 26479 1924
rect 26421 1915 26479 1921
rect 27982 1912 27988 1924
rect 28040 1912 28046 1964
rect 26697 1887 26755 1893
rect 26697 1884 26709 1887
rect 26160 1856 26709 1884
rect 25317 1847 25375 1853
rect 26697 1853 26709 1856
rect 26743 1853 26755 1887
rect 26697 1847 26755 1853
rect 21784 1788 24440 1816
rect 21784 1776 21790 1788
rect 24854 1776 24860 1828
rect 24912 1816 24918 1828
rect 25332 1816 25360 1847
rect 24912 1788 25360 1816
rect 24912 1776 24918 1788
rect 26510 1776 26516 1828
rect 26568 1776 26574 1828
rect 15746 1708 15752 1760
rect 15804 1748 15810 1760
rect 18966 1748 18972 1760
rect 15804 1720 18972 1748
rect 15804 1708 15810 1720
rect 18966 1708 18972 1720
rect 19024 1708 19030 1760
rect 19150 1708 19156 1760
rect 19208 1748 19214 1760
rect 19613 1751 19671 1757
rect 19613 1748 19625 1751
rect 19208 1720 19625 1748
rect 19208 1708 19214 1720
rect 19613 1717 19625 1720
rect 19659 1717 19671 1751
rect 19613 1711 19671 1717
rect 20806 1708 20812 1760
rect 20864 1748 20870 1760
rect 26528 1748 26556 1776
rect 20864 1720 26556 1748
rect 20864 1708 20870 1720
rect 552 1658 31808 1680
rect 552 1606 8172 1658
rect 8224 1606 8236 1658
rect 8288 1606 8300 1658
rect 8352 1606 8364 1658
rect 8416 1606 8428 1658
rect 8480 1606 15946 1658
rect 15998 1606 16010 1658
rect 16062 1606 16074 1658
rect 16126 1606 16138 1658
rect 16190 1606 16202 1658
rect 16254 1606 23720 1658
rect 23772 1606 23784 1658
rect 23836 1606 23848 1658
rect 23900 1606 23912 1658
rect 23964 1606 23976 1658
rect 24028 1606 31494 1658
rect 31546 1606 31558 1658
rect 31610 1606 31622 1658
rect 31674 1606 31686 1658
rect 31738 1606 31750 1658
rect 31802 1606 31808 1658
rect 552 1584 31808 1606
rect 18969 1547 19027 1553
rect 18969 1513 18981 1547
rect 19015 1544 19027 1547
rect 19242 1544 19248 1556
rect 19015 1516 19248 1544
rect 19015 1513 19027 1516
rect 18969 1507 19027 1513
rect 19242 1504 19248 1516
rect 19300 1504 19306 1556
rect 19334 1504 19340 1556
rect 19392 1504 19398 1556
rect 20438 1544 20444 1556
rect 19536 1516 20444 1544
rect 14182 1436 14188 1488
rect 14240 1476 14246 1488
rect 14240 1448 19288 1476
rect 14240 1436 14246 1448
rect 18969 1411 19027 1417
rect 18969 1377 18981 1411
rect 19015 1408 19027 1411
rect 19150 1408 19156 1420
rect 19015 1380 19156 1408
rect 19015 1377 19027 1380
rect 18969 1371 19027 1377
rect 19150 1368 19156 1380
rect 19208 1368 19214 1420
rect 19058 1300 19064 1352
rect 19116 1300 19122 1352
rect 19260 1340 19288 1448
rect 19352 1417 19380 1504
rect 19536 1417 19564 1516
rect 20438 1504 20444 1516
rect 20496 1504 20502 1556
rect 21358 1504 21364 1556
rect 21416 1544 21422 1556
rect 26234 1544 26240 1556
rect 21416 1516 26240 1544
rect 21416 1504 21422 1516
rect 26234 1504 26240 1516
rect 26292 1504 26298 1556
rect 21818 1476 21824 1488
rect 19628 1448 21824 1476
rect 19337 1411 19395 1417
rect 19337 1377 19349 1411
rect 19383 1377 19395 1411
rect 19337 1371 19395 1377
rect 19521 1411 19579 1417
rect 19521 1377 19533 1411
rect 19567 1377 19579 1411
rect 19521 1371 19579 1377
rect 19628 1340 19656 1448
rect 21818 1436 21824 1448
rect 21876 1436 21882 1488
rect 19702 1368 19708 1420
rect 19760 1368 19766 1420
rect 19260 1312 19656 1340
rect 19245 1207 19303 1213
rect 19245 1173 19257 1207
rect 19291 1204 19303 1207
rect 19521 1207 19579 1213
rect 19521 1204 19533 1207
rect 19291 1176 19533 1204
rect 19291 1173 19303 1176
rect 19245 1167 19303 1173
rect 19521 1173 19533 1176
rect 19567 1173 19579 1207
rect 19521 1167 19579 1173
rect 552 1114 31648 1136
rect 552 1062 4285 1114
rect 4337 1062 4349 1114
rect 4401 1062 4413 1114
rect 4465 1062 4477 1114
rect 4529 1062 4541 1114
rect 4593 1062 12059 1114
rect 12111 1062 12123 1114
rect 12175 1062 12187 1114
rect 12239 1062 12251 1114
rect 12303 1062 12315 1114
rect 12367 1062 19833 1114
rect 19885 1062 19897 1114
rect 19949 1062 19961 1114
rect 20013 1062 20025 1114
rect 20077 1062 20089 1114
rect 20141 1062 27607 1114
rect 27659 1062 27671 1114
rect 27723 1062 27735 1114
rect 27787 1062 27799 1114
rect 27851 1062 27863 1114
rect 27915 1062 31648 1114
rect 552 1040 31648 1062
rect 552 570 31808 592
rect 552 518 8172 570
rect 8224 518 8236 570
rect 8288 518 8300 570
rect 8352 518 8364 570
rect 8416 518 8428 570
rect 8480 518 15946 570
rect 15998 518 16010 570
rect 16062 518 16074 570
rect 16126 518 16138 570
rect 16190 518 16202 570
rect 16254 518 23720 570
rect 23772 518 23784 570
rect 23836 518 23848 570
rect 23900 518 23912 570
rect 23964 518 23976 570
rect 24028 518 31494 570
rect 31546 518 31558 570
rect 31610 518 31622 570
rect 31674 518 31686 570
rect 31738 518 31750 570
rect 31802 518 31808 570
rect 552 496 31808 518
<< via1 >>
rect 5080 21972 5132 22024
rect 15200 21972 15252 22024
rect 24584 21972 24636 22024
rect 26884 21972 26936 22024
rect 30380 21972 30432 22024
rect 4068 21904 4120 21956
rect 10140 21904 10192 21956
rect 10324 21904 10376 21956
rect 3516 21836 3568 21888
rect 15844 21836 15896 21888
rect 25320 21836 25372 21888
rect 30840 21836 30892 21888
rect 4285 21734 4337 21786
rect 4349 21734 4401 21786
rect 4413 21734 4465 21786
rect 4477 21734 4529 21786
rect 4541 21734 4593 21786
rect 12059 21734 12111 21786
rect 12123 21734 12175 21786
rect 12187 21734 12239 21786
rect 12251 21734 12303 21786
rect 12315 21734 12367 21786
rect 19833 21734 19885 21786
rect 19897 21734 19949 21786
rect 19961 21734 20013 21786
rect 20025 21734 20077 21786
rect 20089 21734 20141 21786
rect 27607 21734 27659 21786
rect 27671 21734 27723 21786
rect 27735 21734 27787 21786
rect 27799 21734 27851 21786
rect 27863 21734 27915 21786
rect 6368 21632 6420 21684
rect 7012 21675 7064 21684
rect 7012 21641 7021 21675
rect 7021 21641 7055 21675
rect 7055 21641 7064 21675
rect 7012 21632 7064 21641
rect 4988 21564 5040 21616
rect 1308 21539 1360 21548
rect 1308 21505 1317 21539
rect 1317 21505 1351 21539
rect 1351 21505 1360 21539
rect 1308 21496 1360 21505
rect 5540 21496 5592 21548
rect 6276 21496 6328 21548
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 2228 21360 2280 21412
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 8852 21632 8904 21684
rect 12532 21675 12584 21684
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 13820 21632 13872 21684
rect 16580 21675 16632 21684
rect 16580 21641 16589 21675
rect 16589 21641 16623 21675
rect 16623 21641 16632 21675
rect 16580 21632 16632 21641
rect 9036 21496 9088 21548
rect 9772 21496 9824 21548
rect 12348 21564 12400 21616
rect 13636 21564 13688 21616
rect 20444 21632 20496 21684
rect 13176 21496 13228 21548
rect 9680 21428 9732 21480
rect 3608 21360 3660 21412
rect 3884 21403 3936 21412
rect 3884 21369 3893 21403
rect 3893 21369 3927 21403
rect 3927 21369 3936 21403
rect 3884 21360 3936 21369
rect 6920 21360 6972 21412
rect 7012 21360 7064 21412
rect 7288 21403 7340 21412
rect 7288 21369 7297 21403
rect 7297 21369 7331 21403
rect 7331 21369 7340 21403
rect 7288 21360 7340 21369
rect 7380 21360 7432 21412
rect 2964 21292 3016 21344
rect 3792 21292 3844 21344
rect 4620 21292 4672 21344
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 6368 21292 6420 21344
rect 7196 21292 7248 21344
rect 10508 21428 10560 21480
rect 13544 21428 13596 21480
rect 13912 21496 13964 21548
rect 20260 21564 20312 21616
rect 20720 21632 20772 21684
rect 22008 21632 22060 21684
rect 28448 21632 28500 21684
rect 21456 21564 21508 21616
rect 15292 21428 15344 21480
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 9128 21292 9180 21344
rect 11244 21360 11296 21412
rect 11336 21360 11388 21412
rect 11704 21360 11756 21412
rect 12348 21360 12400 21412
rect 12992 21360 13044 21412
rect 13268 21403 13320 21412
rect 13268 21369 13277 21403
rect 13277 21369 13311 21403
rect 13311 21369 13320 21403
rect 13268 21360 13320 21369
rect 12256 21292 12308 21344
rect 13360 21292 13412 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 14188 21292 14240 21301
rect 14372 21335 14424 21344
rect 14372 21301 14399 21335
rect 14399 21301 14424 21335
rect 14372 21292 14424 21301
rect 14556 21403 14608 21412
rect 14556 21369 14565 21403
rect 14565 21369 14599 21403
rect 14599 21369 14608 21403
rect 14556 21360 14608 21369
rect 15108 21360 15160 21412
rect 16672 21292 16724 21344
rect 19064 21471 19116 21480
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 19156 21471 19208 21480
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 19524 21428 19576 21480
rect 20536 21428 20588 21480
rect 21456 21428 21508 21480
rect 23940 21428 23992 21480
rect 20996 21360 21048 21412
rect 25872 21496 25924 21548
rect 24676 21471 24728 21480
rect 24676 21437 24685 21471
rect 24685 21437 24719 21471
rect 24719 21437 24728 21471
rect 24676 21428 24728 21437
rect 24860 21428 24912 21480
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 26608 21471 26660 21480
rect 26608 21437 26617 21471
rect 26617 21437 26651 21471
rect 26651 21437 26660 21471
rect 26608 21428 26660 21437
rect 27436 21471 27488 21480
rect 27436 21437 27445 21471
rect 27445 21437 27479 21471
rect 27479 21437 27488 21471
rect 27436 21428 27488 21437
rect 27528 21428 27580 21480
rect 28816 21496 28868 21548
rect 27712 21471 27764 21480
rect 27712 21437 27721 21471
rect 27721 21437 27755 21471
rect 27755 21437 27764 21471
rect 27712 21428 27764 21437
rect 28080 21471 28132 21480
rect 28080 21437 28089 21471
rect 28089 21437 28123 21471
rect 28123 21437 28132 21471
rect 28080 21428 28132 21437
rect 29000 21471 29052 21480
rect 29000 21437 29009 21471
rect 29009 21437 29043 21471
rect 29043 21437 29052 21471
rect 29000 21428 29052 21437
rect 29184 21428 29236 21480
rect 19616 21292 19668 21344
rect 20628 21292 20680 21344
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 24860 21292 24912 21344
rect 26332 21360 26384 21412
rect 29736 21471 29788 21480
rect 29736 21437 29745 21471
rect 29745 21437 29779 21471
rect 29779 21437 29788 21471
rect 29736 21428 29788 21437
rect 30012 21471 30064 21480
rect 30012 21437 30021 21471
rect 30021 21437 30055 21471
rect 30055 21437 30064 21471
rect 30012 21428 30064 21437
rect 30288 21428 30340 21480
rect 29644 21360 29696 21412
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 27252 21335 27304 21344
rect 27252 21301 27261 21335
rect 27261 21301 27295 21335
rect 27295 21301 27304 21335
rect 27252 21292 27304 21301
rect 29000 21292 29052 21344
rect 29368 21335 29420 21344
rect 29368 21301 29377 21335
rect 29377 21301 29411 21335
rect 29411 21301 29420 21335
rect 29368 21292 29420 21301
rect 30288 21335 30340 21344
rect 30288 21301 30297 21335
rect 30297 21301 30331 21335
rect 30331 21301 30340 21335
rect 30288 21292 30340 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 15946 21190 15998 21242
rect 16010 21190 16062 21242
rect 16074 21190 16126 21242
rect 16138 21190 16190 21242
rect 16202 21190 16254 21242
rect 23720 21190 23772 21242
rect 23784 21190 23836 21242
rect 23848 21190 23900 21242
rect 23912 21190 23964 21242
rect 23976 21190 24028 21242
rect 31494 21190 31546 21242
rect 31558 21190 31610 21242
rect 31622 21190 31674 21242
rect 31686 21190 31738 21242
rect 31750 21190 31802 21242
rect 2136 21088 2188 21140
rect 3884 21088 3936 21140
rect 3976 21131 4028 21140
rect 3976 21097 3985 21131
rect 3985 21097 4019 21131
rect 4019 21097 4028 21131
rect 3976 21088 4028 21097
rect 4068 21131 4120 21140
rect 4068 21097 4077 21131
rect 4077 21097 4111 21131
rect 4111 21097 4120 21131
rect 4068 21088 4120 21097
rect 4988 21131 5040 21140
rect 4988 21097 4997 21131
rect 4997 21097 5031 21131
rect 5031 21097 5040 21131
rect 4988 21088 5040 21097
rect 5080 21131 5132 21140
rect 5080 21097 5089 21131
rect 5089 21097 5123 21131
rect 5123 21097 5132 21131
rect 5080 21088 5132 21097
rect 6460 21131 6512 21140
rect 6460 21097 6469 21131
rect 6469 21097 6503 21131
rect 6503 21097 6512 21131
rect 6460 21088 6512 21097
rect 6644 21088 6696 21140
rect 2228 20952 2280 21004
rect 4712 21020 4764 21072
rect 7012 21063 7064 21072
rect 7012 21029 7021 21063
rect 7021 21029 7055 21063
rect 7055 21029 7064 21063
rect 7012 21020 7064 21029
rect 8944 21088 8996 21140
rect 9036 21088 9088 21140
rect 9404 21088 9456 21140
rect 13084 21088 13136 21140
rect 13176 21088 13228 21140
rect 13728 21131 13780 21140
rect 13728 21097 13753 21131
rect 13753 21097 13780 21131
rect 13728 21088 13780 21097
rect 14372 21088 14424 21140
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 1216 20884 1268 20936
rect 3792 20884 3844 20936
rect 5448 20995 5500 21004
rect 5448 20961 5457 20995
rect 5457 20961 5491 20995
rect 5491 20961 5500 20995
rect 5448 20952 5500 20961
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 6276 20884 6328 20936
rect 940 20748 992 20800
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 5632 20791 5684 20800
rect 5632 20757 5641 20791
rect 5641 20757 5675 20791
rect 5675 20757 5684 20791
rect 5632 20748 5684 20757
rect 6092 20748 6144 20800
rect 6920 20952 6972 21004
rect 10324 20952 10376 21004
rect 10600 20952 10652 21004
rect 10784 20952 10836 21004
rect 11244 20952 11296 21004
rect 12256 21020 12308 21072
rect 14740 21020 14792 21072
rect 18512 21131 18564 21140
rect 18512 21097 18521 21131
rect 18521 21097 18555 21131
rect 18555 21097 18564 21131
rect 18512 21088 18564 21097
rect 19064 21131 19116 21140
rect 19064 21097 19073 21131
rect 19073 21097 19107 21131
rect 19107 21097 19116 21131
rect 19064 21088 19116 21097
rect 19248 21131 19300 21140
rect 19248 21097 19275 21131
rect 19275 21097 19300 21131
rect 19248 21088 19300 21097
rect 16028 21020 16080 21072
rect 12348 20952 12400 21004
rect 12808 20952 12860 21004
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 13268 20952 13320 20961
rect 13912 20952 13964 21004
rect 14096 20952 14148 21004
rect 14648 20952 14700 21004
rect 15200 20995 15252 21004
rect 15200 20961 15210 20995
rect 15210 20961 15244 20995
rect 15244 20961 15252 20995
rect 15200 20952 15252 20961
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 7288 20884 7340 20936
rect 9036 20927 9088 20936
rect 9036 20893 9045 20927
rect 9045 20893 9079 20927
rect 9079 20893 9088 20927
rect 9036 20884 9088 20893
rect 9680 20884 9732 20936
rect 9956 20884 10008 20936
rect 9772 20816 9824 20868
rect 10876 20816 10928 20868
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 13084 20884 13136 20936
rect 13820 20884 13872 20936
rect 15660 20952 15712 21004
rect 15844 20952 15896 21004
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 16488 20995 16540 21004
rect 16488 20961 16497 20995
rect 16497 20961 16531 20995
rect 16531 20961 16540 20995
rect 16488 20952 16540 20961
rect 16672 21063 16724 21072
rect 16672 21029 16681 21063
rect 16681 21029 16715 21063
rect 16715 21029 16724 21063
rect 16672 21020 16724 21029
rect 17960 21020 18012 21072
rect 20536 21088 20588 21140
rect 19432 21063 19484 21072
rect 19432 21029 19441 21063
rect 19441 21029 19475 21063
rect 19475 21029 19484 21063
rect 19432 21020 19484 21029
rect 18236 20952 18288 21004
rect 18328 20952 18380 21004
rect 11980 20816 12032 20868
rect 16396 20884 16448 20936
rect 10784 20748 10836 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 11612 20748 11664 20800
rect 12394 20748 12446 20800
rect 13728 20791 13780 20800
rect 13728 20757 13737 20791
rect 13737 20757 13771 20791
rect 13771 20757 13780 20791
rect 13728 20748 13780 20757
rect 17316 20748 17368 20800
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 19064 20884 19116 20936
rect 19340 20816 19392 20868
rect 20260 20995 20312 21004
rect 20260 20961 20269 20995
rect 20269 20961 20303 20995
rect 20303 20961 20312 20995
rect 20260 20952 20312 20961
rect 20720 20952 20772 21004
rect 21456 21063 21508 21072
rect 21456 21029 21465 21063
rect 21465 21029 21499 21063
rect 21499 21029 21508 21063
rect 22376 21088 22428 21140
rect 21456 21020 21508 21029
rect 21824 20952 21876 21004
rect 22468 21020 22520 21072
rect 23848 21020 23900 21072
rect 24124 21088 24176 21140
rect 22376 20884 22428 20936
rect 22836 20995 22888 21004
rect 22836 20961 22845 20995
rect 22845 20961 22879 20995
rect 22879 20961 22888 20995
rect 22836 20952 22888 20961
rect 22928 20995 22980 21004
rect 22928 20961 22937 20995
rect 22937 20961 22971 20995
rect 22971 20961 22980 20995
rect 22928 20952 22980 20961
rect 23296 20995 23348 21004
rect 23296 20961 23305 20995
rect 23305 20961 23339 20995
rect 23339 20961 23348 20995
rect 23296 20952 23348 20961
rect 23388 20952 23440 21004
rect 23572 20995 23624 21004
rect 23572 20961 23581 20995
rect 23581 20961 23615 20995
rect 23615 20961 23624 20995
rect 23572 20952 23624 20961
rect 24492 20995 24544 21004
rect 24492 20961 24501 20995
rect 24501 20961 24535 20995
rect 24535 20961 24544 20995
rect 24492 20952 24544 20961
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 23664 20884 23716 20936
rect 21916 20816 21968 20868
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 25412 20995 25464 21004
rect 25412 20961 25421 20995
rect 25421 20961 25455 20995
rect 25455 20961 25464 20995
rect 25412 20952 25464 20961
rect 25504 20995 25556 21004
rect 25504 20961 25513 20995
rect 25513 20961 25547 20995
rect 25547 20961 25556 20995
rect 25504 20952 25556 20961
rect 25688 20995 25740 21004
rect 25688 20961 25697 20995
rect 25697 20961 25731 20995
rect 25731 20961 25740 20995
rect 25688 20952 25740 20961
rect 25780 20995 25832 21004
rect 25780 20961 25789 20995
rect 25789 20961 25823 20995
rect 25823 20961 25832 20995
rect 25780 20952 25832 20961
rect 18788 20748 18840 20800
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 23848 20816 23900 20868
rect 26700 20995 26752 21004
rect 26700 20961 26709 20995
rect 26709 20961 26743 20995
rect 26743 20961 26752 20995
rect 26700 20952 26752 20961
rect 26884 21088 26936 21140
rect 27068 21020 27120 21072
rect 27344 21020 27396 21072
rect 29184 21088 29236 21140
rect 30840 21131 30892 21140
rect 30840 21097 30849 21131
rect 30849 21097 30883 21131
rect 30883 21097 30892 21131
rect 30840 21088 30892 21097
rect 27804 20952 27856 21004
rect 27896 20995 27948 21004
rect 27896 20961 27904 20995
rect 27904 20961 27938 20995
rect 27938 20961 27948 20995
rect 27896 20952 27948 20961
rect 29092 21020 29144 21072
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 28540 20952 28592 21004
rect 30932 20952 30984 21004
rect 30564 20927 30616 20936
rect 25596 20816 25648 20868
rect 30564 20893 30573 20927
rect 30573 20893 30607 20927
rect 30607 20893 30616 20927
rect 30564 20884 30616 20893
rect 27344 20791 27396 20800
rect 27344 20757 27353 20791
rect 27353 20757 27387 20791
rect 27387 20757 27396 20791
rect 27344 20748 27396 20757
rect 27804 20748 27856 20800
rect 28080 20748 28132 20800
rect 30472 20791 30524 20800
rect 30472 20757 30481 20791
rect 30481 20757 30515 20791
rect 30515 20757 30524 20791
rect 30472 20748 30524 20757
rect 4285 20646 4337 20698
rect 4349 20646 4401 20698
rect 4413 20646 4465 20698
rect 4477 20646 4529 20698
rect 4541 20646 4593 20698
rect 12059 20646 12111 20698
rect 12123 20646 12175 20698
rect 12187 20646 12239 20698
rect 12251 20646 12303 20698
rect 12315 20646 12367 20698
rect 19833 20646 19885 20698
rect 19897 20646 19949 20698
rect 19961 20646 20013 20698
rect 20025 20646 20077 20698
rect 20089 20646 20141 20698
rect 27607 20646 27659 20698
rect 27671 20646 27723 20698
rect 27735 20646 27787 20698
rect 27799 20646 27851 20698
rect 27863 20646 27915 20698
rect 2688 20544 2740 20596
rect 1124 20247 1176 20256
rect 1124 20213 1133 20247
rect 1133 20213 1167 20247
rect 1167 20213 1176 20247
rect 1124 20204 1176 20213
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 2504 20408 2556 20460
rect 2872 20340 2924 20392
rect 2780 20272 2832 20324
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 2596 20204 2648 20256
rect 4620 20544 4672 20596
rect 4528 20476 4580 20528
rect 3608 20408 3660 20460
rect 4160 20408 4212 20460
rect 7196 20408 7248 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8668 20587 8720 20596
rect 8668 20553 8677 20587
rect 8677 20553 8711 20587
rect 8711 20553 8720 20587
rect 8668 20544 8720 20553
rect 10508 20587 10560 20596
rect 10508 20553 10517 20587
rect 10517 20553 10551 20587
rect 10551 20553 10560 20587
rect 10508 20544 10560 20553
rect 11796 20544 11848 20596
rect 8024 20476 8076 20528
rect 14004 20544 14056 20596
rect 15292 20544 15344 20596
rect 16028 20544 16080 20596
rect 16304 20587 16356 20596
rect 16304 20553 16313 20587
rect 16313 20553 16347 20587
rect 16347 20553 16356 20587
rect 16304 20544 16356 20553
rect 17960 20544 18012 20596
rect 18236 20544 18288 20596
rect 3240 20272 3292 20324
rect 4988 20272 5040 20324
rect 4160 20204 4212 20256
rect 4528 20204 4580 20256
rect 6460 20204 6512 20256
rect 6920 20204 6972 20256
rect 7840 20204 7892 20256
rect 9404 20340 9456 20392
rect 8852 20272 8904 20324
rect 9036 20272 9088 20324
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 10784 20408 10836 20460
rect 13820 20476 13872 20528
rect 16580 20476 16632 20528
rect 12992 20408 13044 20460
rect 15752 20451 15804 20460
rect 8576 20204 8628 20256
rect 11612 20340 11664 20392
rect 12900 20340 12952 20392
rect 13176 20383 13228 20392
rect 13176 20349 13185 20383
rect 13185 20349 13219 20383
rect 13219 20349 13228 20383
rect 13176 20340 13228 20349
rect 14188 20340 14240 20392
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 12256 20272 12308 20324
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 14740 20383 14792 20392
rect 14740 20349 14749 20383
rect 14749 20349 14783 20383
rect 14783 20349 14792 20383
rect 14740 20340 14792 20349
rect 14832 20383 14884 20392
rect 14832 20349 14841 20383
rect 14841 20349 14875 20383
rect 14875 20349 14884 20383
rect 14832 20340 14884 20349
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 15108 20340 15160 20392
rect 15568 20340 15620 20392
rect 15660 20383 15712 20392
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 15936 20383 15988 20392
rect 15936 20349 15945 20383
rect 15945 20349 15979 20383
rect 15979 20349 15988 20383
rect 15936 20340 15988 20349
rect 16488 20340 16540 20392
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 17040 20340 17092 20392
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 17592 20340 17644 20392
rect 18420 20476 18472 20528
rect 18604 20476 18656 20528
rect 19800 20476 19852 20528
rect 20260 20476 20312 20528
rect 20720 20544 20772 20596
rect 21916 20544 21968 20596
rect 22560 20544 22612 20596
rect 23296 20544 23348 20596
rect 23572 20544 23624 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 25136 20544 25188 20596
rect 18512 20408 18564 20460
rect 19156 20408 19208 20460
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 10600 20204 10652 20256
rect 11612 20204 11664 20256
rect 15384 20272 15436 20324
rect 17868 20315 17920 20324
rect 14924 20204 14976 20256
rect 17868 20281 17895 20315
rect 17895 20281 17920 20315
rect 17868 20272 17920 20281
rect 19708 20340 19760 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 20720 20340 20772 20392
rect 21272 20383 21324 20392
rect 21272 20349 21281 20383
rect 21281 20349 21315 20383
rect 21315 20349 21324 20383
rect 21272 20340 21324 20349
rect 16580 20204 16632 20256
rect 16948 20204 17000 20256
rect 17500 20204 17552 20256
rect 20904 20315 20956 20324
rect 20904 20281 20913 20315
rect 20913 20281 20947 20315
rect 20947 20281 20956 20315
rect 20904 20272 20956 20281
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 25504 20476 25556 20528
rect 22192 20408 22244 20460
rect 23572 20408 23624 20460
rect 23664 20408 23716 20460
rect 24308 20340 24360 20392
rect 23388 20272 23440 20324
rect 23756 20272 23808 20324
rect 18328 20204 18380 20256
rect 19340 20204 19392 20256
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20260 20204 20312 20256
rect 20536 20204 20588 20256
rect 21456 20204 21508 20256
rect 22468 20204 22520 20256
rect 22652 20204 22704 20256
rect 24584 20408 24636 20460
rect 25596 20408 25648 20460
rect 28448 20408 28500 20460
rect 29092 20544 29144 20596
rect 29460 20587 29512 20596
rect 29460 20553 29469 20587
rect 29469 20553 29503 20587
rect 29503 20553 29512 20587
rect 29460 20544 29512 20553
rect 30472 20544 30524 20596
rect 30564 20519 30616 20528
rect 30564 20485 30573 20519
rect 30573 20485 30607 20519
rect 30607 20485 30616 20519
rect 30564 20476 30616 20485
rect 24952 20340 25004 20392
rect 27068 20340 27120 20392
rect 24860 20272 24912 20324
rect 28632 20340 28684 20392
rect 30196 20408 30248 20460
rect 30840 20408 30892 20460
rect 29184 20315 29236 20324
rect 29184 20281 29219 20315
rect 29219 20281 29236 20315
rect 29920 20340 29972 20392
rect 30748 20383 30800 20392
rect 30748 20349 30757 20383
rect 30757 20349 30791 20383
rect 30791 20349 30800 20383
rect 30748 20340 30800 20349
rect 31024 20383 31076 20392
rect 31024 20349 31033 20383
rect 31033 20349 31067 20383
rect 31067 20349 31076 20383
rect 31024 20340 31076 20349
rect 29184 20272 29236 20281
rect 29552 20272 29604 20324
rect 30288 20272 30340 20324
rect 25320 20204 25372 20256
rect 25688 20204 25740 20256
rect 26792 20204 26844 20256
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 28356 20204 28408 20256
rect 30104 20204 30156 20256
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 15946 20102 15998 20154
rect 16010 20102 16062 20154
rect 16074 20102 16126 20154
rect 16138 20102 16190 20154
rect 16202 20102 16254 20154
rect 23720 20102 23772 20154
rect 23784 20102 23836 20154
rect 23848 20102 23900 20154
rect 23912 20102 23964 20154
rect 23976 20102 24028 20154
rect 31494 20102 31546 20154
rect 31558 20102 31610 20154
rect 31622 20102 31674 20154
rect 31686 20102 31738 20154
rect 31750 20102 31802 20154
rect 1124 20000 1176 20052
rect 3976 20000 4028 20052
rect 3332 19932 3384 19984
rect 4988 19932 5040 19984
rect 9036 20000 9088 20052
rect 5632 19932 5684 19984
rect 6920 19932 6972 19984
rect 7472 19932 7524 19984
rect 2228 19864 2280 19916
rect 2688 19864 2740 19916
rect 3608 19907 3660 19916
rect 3608 19873 3617 19907
rect 3617 19873 3651 19907
rect 3651 19873 3660 19907
rect 3608 19864 3660 19873
rect 3056 19796 3108 19848
rect 5540 19864 5592 19916
rect 7840 19864 7892 19916
rect 6184 19796 6236 19848
rect 6644 19796 6696 19848
rect 8944 19796 8996 19848
rect 940 19660 992 19712
rect 3608 19728 3660 19780
rect 10416 20043 10468 20052
rect 10416 20009 10425 20043
rect 10425 20009 10459 20043
rect 10459 20009 10468 20043
rect 10416 20000 10468 20009
rect 10048 19864 10100 19916
rect 12256 20000 12308 20052
rect 13176 20000 13228 20052
rect 16488 20000 16540 20052
rect 17684 20000 17736 20052
rect 18512 20000 18564 20052
rect 18880 20000 18932 20052
rect 21640 20000 21692 20052
rect 23296 20000 23348 20052
rect 24952 20000 25004 20052
rect 26792 20000 26844 20052
rect 10968 19864 11020 19916
rect 11152 19864 11204 19916
rect 11612 19864 11664 19916
rect 11980 19864 12032 19916
rect 12256 19907 12308 19916
rect 12256 19873 12265 19907
rect 12265 19873 12299 19907
rect 12299 19873 12308 19907
rect 12256 19864 12308 19873
rect 12808 19932 12860 19984
rect 12992 19932 13044 19984
rect 13084 19932 13136 19984
rect 14832 19932 14884 19984
rect 17316 19932 17368 19984
rect 15568 19864 15620 19916
rect 17040 19864 17092 19916
rect 17500 19864 17552 19916
rect 17960 19864 18012 19916
rect 18420 19932 18472 19984
rect 19156 19932 19208 19984
rect 21548 19932 21600 19984
rect 22284 19932 22336 19984
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 11796 19796 11848 19848
rect 12532 19796 12584 19848
rect 12624 19796 12676 19848
rect 16488 19796 16540 19848
rect 17868 19796 17920 19848
rect 18144 19796 18196 19848
rect 9496 19728 9548 19780
rect 2688 19660 2740 19712
rect 3976 19660 4028 19712
rect 5356 19660 5408 19712
rect 6920 19660 6972 19712
rect 10232 19728 10284 19780
rect 14556 19728 14608 19780
rect 17500 19728 17552 19780
rect 18880 19907 18932 19916
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 19340 19864 19392 19916
rect 19432 19864 19484 19916
rect 19524 19864 19576 19916
rect 20076 19907 20128 19916
rect 20076 19873 20085 19907
rect 20085 19873 20119 19907
rect 20119 19873 20128 19907
rect 20076 19864 20128 19873
rect 20720 19864 20772 19916
rect 21180 19864 21232 19916
rect 21456 19864 21508 19916
rect 21916 19864 21968 19916
rect 19800 19771 19852 19780
rect 19800 19737 19809 19771
rect 19809 19737 19843 19771
rect 19843 19737 19852 19771
rect 19800 19728 19852 19737
rect 20904 19796 20956 19848
rect 22100 19839 22152 19848
rect 22100 19805 22108 19839
rect 22108 19805 22142 19839
rect 22142 19805 22152 19839
rect 22100 19796 22152 19805
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 24400 19932 24452 19984
rect 24676 19932 24728 19984
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 23480 19864 23532 19916
rect 23940 19864 23992 19916
rect 24308 19907 24360 19916
rect 24308 19873 24317 19907
rect 24317 19873 24351 19907
rect 24351 19873 24360 19907
rect 24308 19864 24360 19873
rect 21456 19728 21508 19780
rect 23020 19796 23072 19848
rect 24768 19907 24820 19916
rect 24768 19873 24777 19907
rect 24777 19873 24811 19907
rect 24811 19873 24820 19907
rect 24768 19864 24820 19873
rect 26700 19932 26752 19984
rect 10600 19660 10652 19712
rect 10968 19703 11020 19712
rect 10968 19669 10977 19703
rect 10977 19669 11011 19703
rect 11011 19669 11020 19703
rect 10968 19660 11020 19669
rect 11060 19660 11112 19712
rect 14188 19660 14240 19712
rect 16396 19660 16448 19712
rect 17408 19660 17460 19712
rect 17868 19660 17920 19712
rect 18512 19660 18564 19712
rect 20812 19660 20864 19712
rect 20904 19660 20956 19712
rect 25136 19796 25188 19848
rect 25320 19907 25372 19916
rect 25320 19873 25329 19907
rect 25329 19873 25363 19907
rect 25363 19873 25372 19907
rect 25320 19864 25372 19873
rect 25596 19864 25648 19916
rect 26332 19864 26384 19916
rect 26516 19864 26568 19916
rect 26608 19907 26660 19916
rect 26608 19873 26617 19907
rect 26617 19873 26651 19907
rect 26651 19873 26660 19907
rect 26608 19864 26660 19873
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 27160 20000 27212 20052
rect 29184 20000 29236 20052
rect 29460 20000 29512 20052
rect 27436 19864 27488 19916
rect 28080 19907 28132 19916
rect 28080 19873 28089 19907
rect 28089 19873 28123 19907
rect 28123 19873 28132 19907
rect 28080 19864 28132 19873
rect 30748 20000 30800 20052
rect 29736 19932 29788 19984
rect 31024 19932 31076 19984
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 30748 19864 30800 19916
rect 28080 19728 28132 19780
rect 28540 19728 28592 19780
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 23756 19660 23808 19712
rect 26056 19660 26108 19712
rect 4285 19558 4337 19610
rect 4349 19558 4401 19610
rect 4413 19558 4465 19610
rect 4477 19558 4529 19610
rect 4541 19558 4593 19610
rect 12059 19558 12111 19610
rect 12123 19558 12175 19610
rect 12187 19558 12239 19610
rect 12251 19558 12303 19610
rect 12315 19558 12367 19610
rect 19833 19558 19885 19610
rect 19897 19558 19949 19610
rect 19961 19558 20013 19610
rect 20025 19558 20077 19610
rect 20089 19558 20141 19610
rect 27607 19558 27659 19610
rect 27671 19558 27723 19610
rect 27735 19558 27787 19610
rect 27799 19558 27851 19610
rect 27863 19558 27915 19610
rect 940 19456 992 19508
rect 3056 19499 3108 19508
rect 3056 19465 3065 19499
rect 3065 19465 3099 19499
rect 3099 19465 3108 19499
rect 3056 19456 3108 19465
rect 2688 19252 2740 19304
rect 4344 19363 4396 19372
rect 4344 19329 4353 19363
rect 4353 19329 4387 19363
rect 4387 19329 4396 19363
rect 4344 19320 4396 19329
rect 4620 19320 4672 19372
rect 1124 19227 1176 19236
rect 1124 19193 1133 19227
rect 1133 19193 1167 19227
rect 1167 19193 1176 19227
rect 1124 19184 1176 19193
rect 3240 19227 3292 19236
rect 3240 19193 3249 19227
rect 3249 19193 3283 19227
rect 3283 19193 3292 19227
rect 3240 19184 3292 19193
rect 5356 19252 5408 19304
rect 6000 19252 6052 19304
rect 7932 19431 7984 19440
rect 7932 19397 7941 19431
rect 7941 19397 7975 19431
rect 7975 19397 7984 19431
rect 7932 19388 7984 19397
rect 9036 19456 9088 19508
rect 10048 19456 10100 19508
rect 10232 19456 10284 19508
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 11428 19456 11480 19508
rect 12808 19456 12860 19508
rect 6276 19320 6328 19372
rect 13636 19456 13688 19508
rect 14372 19456 14424 19508
rect 14740 19456 14792 19508
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 15384 19456 15436 19508
rect 16488 19456 16540 19508
rect 9956 19320 10008 19372
rect 7380 19252 7432 19304
rect 8024 19252 8076 19304
rect 10600 19252 10652 19304
rect 10968 19252 11020 19304
rect 11428 19295 11480 19304
rect 11428 19261 11437 19295
rect 11437 19261 11471 19295
rect 11471 19261 11480 19295
rect 11428 19252 11480 19261
rect 12624 19320 12676 19372
rect 14464 19388 14516 19440
rect 17500 19388 17552 19440
rect 18880 19456 18932 19508
rect 19064 19456 19116 19508
rect 20904 19456 20956 19508
rect 18604 19388 18656 19440
rect 19432 19388 19484 19440
rect 11888 19295 11940 19304
rect 11888 19261 11897 19295
rect 11897 19261 11931 19295
rect 11931 19261 11940 19295
rect 11888 19252 11940 19261
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 3332 19116 3384 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 5448 19184 5500 19236
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 4896 19159 4948 19168
rect 4896 19125 4905 19159
rect 4905 19125 4939 19159
rect 4939 19125 4948 19159
rect 4896 19116 4948 19125
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 5356 19116 5408 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 6000 19116 6052 19168
rect 6644 19227 6696 19236
rect 6644 19193 6653 19227
rect 6653 19193 6687 19227
rect 6687 19193 6696 19227
rect 6644 19184 6696 19193
rect 7932 19184 7984 19236
rect 9036 19184 9088 19236
rect 6552 19116 6604 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 9864 19227 9916 19236
rect 9864 19193 9873 19227
rect 9873 19193 9907 19227
rect 9907 19193 9916 19227
rect 9864 19184 9916 19193
rect 11612 19227 11664 19236
rect 11612 19193 11621 19227
rect 11621 19193 11655 19227
rect 11655 19193 11664 19227
rect 11612 19184 11664 19193
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 13636 19252 13688 19304
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 13912 19252 13964 19261
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 16396 19320 16448 19329
rect 17132 19320 17184 19372
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 14648 19252 14700 19304
rect 13728 19184 13780 19236
rect 13820 19116 13872 19168
rect 14740 19184 14792 19236
rect 15292 19252 15344 19304
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 15200 19184 15252 19236
rect 16396 19184 16448 19236
rect 16580 19295 16632 19304
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 16856 19252 16908 19304
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 16580 19116 16632 19168
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 18420 19320 18472 19372
rect 19616 19388 19668 19440
rect 22284 19456 22336 19508
rect 23388 19456 23440 19508
rect 24860 19499 24912 19508
rect 24860 19465 24869 19499
rect 24869 19465 24903 19499
rect 24903 19465 24912 19499
rect 24860 19456 24912 19465
rect 17500 19252 17552 19304
rect 17684 19252 17736 19304
rect 18972 19252 19024 19304
rect 19064 19252 19116 19304
rect 17776 19184 17828 19236
rect 18604 19184 18656 19236
rect 17684 19116 17736 19168
rect 17868 19116 17920 19168
rect 19432 19116 19484 19168
rect 19708 19184 19760 19236
rect 20720 19320 20772 19372
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20628 19252 20680 19304
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 21640 19363 21692 19372
rect 21640 19329 21649 19363
rect 21649 19329 21683 19363
rect 21683 19329 21692 19363
rect 21640 19320 21692 19329
rect 22100 19388 22152 19440
rect 24768 19388 24820 19440
rect 25136 19388 25188 19440
rect 26608 19456 26660 19508
rect 29460 19456 29512 19508
rect 29920 19499 29972 19508
rect 29920 19465 29929 19499
rect 29929 19465 29963 19499
rect 29963 19465 29972 19499
rect 29920 19456 29972 19465
rect 22192 19320 22244 19372
rect 22652 19320 22704 19372
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 23940 19320 23992 19372
rect 24216 19320 24268 19372
rect 27436 19388 27488 19440
rect 29092 19388 29144 19440
rect 30288 19388 30340 19440
rect 27344 19320 27396 19372
rect 20720 19184 20772 19236
rect 21732 19295 21784 19304
rect 21732 19261 21741 19295
rect 21741 19261 21775 19295
rect 21775 19261 21784 19295
rect 21732 19252 21784 19261
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 19800 19116 19852 19168
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 20168 19116 20220 19168
rect 20352 19116 20404 19168
rect 22192 19184 22244 19236
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 23204 19252 23256 19304
rect 23664 19252 23716 19304
rect 23848 19295 23900 19304
rect 23848 19261 23857 19295
rect 23857 19261 23891 19295
rect 23891 19261 23900 19295
rect 23848 19252 23900 19261
rect 22652 19184 22704 19236
rect 22376 19116 22428 19168
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 23112 19184 23164 19236
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 25872 19252 25924 19304
rect 26056 19252 26108 19304
rect 26148 19227 26200 19236
rect 26148 19193 26157 19227
rect 26157 19193 26191 19227
rect 26191 19193 26200 19227
rect 26148 19184 26200 19193
rect 23296 19116 23348 19168
rect 24124 19116 24176 19168
rect 26424 19295 26476 19304
rect 26424 19261 26433 19295
rect 26433 19261 26467 19295
rect 26467 19261 26476 19295
rect 26424 19252 26476 19261
rect 26884 19295 26936 19304
rect 26884 19261 26893 19295
rect 26893 19261 26927 19295
rect 26927 19261 26936 19295
rect 26884 19252 26936 19261
rect 27160 19295 27212 19304
rect 27160 19261 27169 19295
rect 27169 19261 27203 19295
rect 27203 19261 27212 19295
rect 27160 19252 27212 19261
rect 29000 19252 29052 19304
rect 29184 19295 29236 19304
rect 29184 19261 29193 19295
rect 29193 19261 29227 19295
rect 29227 19261 29236 19295
rect 29184 19252 29236 19261
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 29368 19295 29420 19304
rect 29368 19261 29377 19295
rect 29377 19261 29411 19295
rect 29411 19261 29420 19295
rect 29368 19252 29420 19261
rect 29644 19295 29696 19304
rect 29644 19261 29653 19295
rect 29653 19261 29687 19295
rect 29687 19261 29696 19295
rect 29644 19252 29696 19261
rect 29828 19252 29880 19304
rect 30196 19252 30248 19304
rect 26700 19116 26752 19168
rect 30840 19320 30892 19372
rect 31024 19320 31076 19372
rect 30656 19252 30708 19304
rect 30656 19159 30708 19168
rect 30656 19125 30665 19159
rect 30665 19125 30699 19159
rect 30699 19125 30708 19159
rect 30656 19116 30708 19125
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 15946 19014 15998 19066
rect 16010 19014 16062 19066
rect 16074 19014 16126 19066
rect 16138 19014 16190 19066
rect 16202 19014 16254 19066
rect 23720 19014 23772 19066
rect 23784 19014 23836 19066
rect 23848 19014 23900 19066
rect 23912 19014 23964 19066
rect 23976 19014 24028 19066
rect 31494 19014 31546 19066
rect 31558 19014 31610 19066
rect 31622 19014 31674 19066
rect 31686 19014 31738 19066
rect 31750 19014 31802 19066
rect 1124 18912 1176 18964
rect 2044 18912 2096 18964
rect 2136 18912 2188 18964
rect 2780 18912 2832 18964
rect 3240 18912 3292 18964
rect 4068 18912 4120 18964
rect 4712 18912 4764 18964
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 5264 18912 5316 18964
rect 6276 18912 6328 18964
rect 8392 18912 8444 18964
rect 8668 18912 8720 18964
rect 2596 18844 2648 18896
rect 3700 18844 3752 18896
rect 7840 18844 7892 18896
rect 3424 18776 3476 18828
rect 3516 18819 3568 18828
rect 3516 18785 3525 18819
rect 3525 18785 3559 18819
rect 3559 18785 3568 18819
rect 3516 18776 3568 18785
rect 1216 18572 1268 18624
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 2872 18640 2924 18692
rect 4068 18708 4120 18760
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 5080 18776 5132 18828
rect 4252 18640 4304 18692
rect 4712 18708 4764 18760
rect 5448 18751 5500 18760
rect 5448 18717 5457 18751
rect 5457 18717 5491 18751
rect 5491 18717 5500 18751
rect 5448 18708 5500 18717
rect 5724 18708 5776 18760
rect 4804 18640 4856 18692
rect 4988 18572 5040 18624
rect 6920 18708 6972 18760
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 8668 18776 8720 18828
rect 9772 18912 9824 18964
rect 9864 18912 9916 18964
rect 11244 18912 11296 18964
rect 10140 18844 10192 18896
rect 12532 18912 12584 18964
rect 17132 18912 17184 18964
rect 17224 18912 17276 18964
rect 17684 18912 17736 18964
rect 17776 18955 17828 18964
rect 17776 18921 17785 18955
rect 17785 18921 17819 18955
rect 17819 18921 17828 18955
rect 17776 18912 17828 18921
rect 12992 18844 13044 18896
rect 16672 18844 16724 18896
rect 10324 18776 10376 18828
rect 11060 18776 11112 18828
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 9956 18708 10008 18760
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 10968 18640 11020 18692
rect 11060 18683 11112 18692
rect 11060 18649 11069 18683
rect 11069 18649 11103 18683
rect 11103 18649 11112 18683
rect 11060 18640 11112 18649
rect 11612 18819 11664 18828
rect 11612 18785 11621 18819
rect 11621 18785 11655 18819
rect 11655 18785 11664 18819
rect 11612 18776 11664 18785
rect 11888 18776 11940 18828
rect 13360 18776 13412 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 13728 18776 13780 18785
rect 13912 18819 13964 18828
rect 13912 18785 13921 18819
rect 13921 18785 13955 18819
rect 13955 18785 13964 18819
rect 13912 18776 13964 18785
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 18328 18912 18380 18964
rect 18420 18912 18472 18964
rect 19524 18912 19576 18964
rect 18144 18844 18196 18896
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 19064 18819 19116 18828
rect 19064 18785 19073 18819
rect 19073 18785 19107 18819
rect 19107 18785 19116 18819
rect 19064 18776 19116 18785
rect 19156 18776 19208 18828
rect 15568 18708 15620 18760
rect 16580 18708 16632 18760
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 7380 18572 7432 18624
rect 8668 18572 8720 18624
rect 9128 18572 9180 18624
rect 11796 18572 11848 18624
rect 12624 18572 12676 18624
rect 13084 18572 13136 18624
rect 14556 18640 14608 18692
rect 15200 18640 15252 18692
rect 16856 18640 16908 18692
rect 17684 18640 17736 18692
rect 18420 18708 18472 18760
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 19800 18776 19852 18828
rect 19984 18819 20036 18828
rect 19984 18785 19993 18819
rect 19993 18785 20027 18819
rect 20027 18785 20036 18819
rect 19984 18776 20036 18785
rect 20904 18912 20956 18964
rect 20996 18912 21048 18964
rect 21640 18912 21692 18964
rect 22376 18912 22428 18964
rect 22560 18912 22612 18964
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 23020 18912 23072 18964
rect 20536 18819 20588 18828
rect 20536 18785 20545 18819
rect 20545 18785 20579 18819
rect 20579 18785 20588 18819
rect 20536 18776 20588 18785
rect 21180 18776 21232 18828
rect 21456 18776 21508 18828
rect 23756 18844 23808 18896
rect 24676 18912 24728 18964
rect 26884 18955 26936 18964
rect 26884 18921 26893 18955
rect 26893 18921 26927 18955
rect 26927 18921 26936 18955
rect 26884 18912 26936 18921
rect 29276 18912 29328 18964
rect 30656 18912 30708 18964
rect 14188 18572 14240 18624
rect 14372 18572 14424 18624
rect 14832 18572 14884 18624
rect 15016 18572 15068 18624
rect 17776 18572 17828 18624
rect 19340 18572 19392 18624
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 21548 18708 21600 18760
rect 19984 18572 20036 18624
rect 20260 18572 20312 18624
rect 21180 18640 21232 18692
rect 23204 18776 23256 18828
rect 26608 18776 26660 18828
rect 20996 18572 21048 18624
rect 21272 18572 21324 18624
rect 22100 18572 22152 18624
rect 22928 18708 22980 18760
rect 24124 18708 24176 18760
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 25044 18751 25096 18760
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 22652 18640 22704 18692
rect 26148 18708 26200 18760
rect 28908 18819 28960 18828
rect 28908 18785 28917 18819
rect 28917 18785 28951 18819
rect 28951 18785 28960 18819
rect 28908 18776 28960 18785
rect 29092 18776 29144 18828
rect 23480 18572 23532 18624
rect 24032 18572 24084 18624
rect 24860 18572 24912 18624
rect 26976 18572 27028 18624
rect 29920 18708 29972 18760
rect 28172 18572 28224 18624
rect 28908 18572 28960 18624
rect 4285 18470 4337 18522
rect 4349 18470 4401 18522
rect 4413 18470 4465 18522
rect 4477 18470 4529 18522
rect 4541 18470 4593 18522
rect 12059 18470 12111 18522
rect 12123 18470 12175 18522
rect 12187 18470 12239 18522
rect 12251 18470 12303 18522
rect 12315 18470 12367 18522
rect 19833 18470 19885 18522
rect 19897 18470 19949 18522
rect 19961 18470 20013 18522
rect 20025 18470 20077 18522
rect 20089 18470 20141 18522
rect 27607 18470 27659 18522
rect 27671 18470 27723 18522
rect 27735 18470 27787 18522
rect 27799 18470 27851 18522
rect 27863 18470 27915 18522
rect 2596 18368 2648 18420
rect 2780 18411 2832 18420
rect 2780 18377 2789 18411
rect 2789 18377 2823 18411
rect 2823 18377 2832 18411
rect 2780 18368 2832 18377
rect 3056 18368 3108 18420
rect 3516 18368 3568 18420
rect 1032 18275 1084 18284
rect 1032 18241 1041 18275
rect 1041 18241 1075 18275
rect 1075 18241 1084 18275
rect 1032 18232 1084 18241
rect 3240 18300 3292 18352
rect 4896 18368 4948 18420
rect 4988 18368 5040 18420
rect 4160 18343 4212 18352
rect 4160 18309 4169 18343
rect 4169 18309 4203 18343
rect 4203 18309 4212 18343
rect 4160 18300 4212 18309
rect 3608 18232 3660 18284
rect 2688 18096 2740 18148
rect 3332 18096 3384 18148
rect 3792 18096 3844 18148
rect 4068 18096 4120 18148
rect 4988 18232 5040 18284
rect 5448 18368 5500 18420
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 10508 18368 10560 18420
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 11060 18368 11112 18420
rect 11612 18368 11664 18420
rect 8300 18300 8352 18352
rect 4436 18139 4488 18148
rect 4436 18105 4445 18139
rect 4445 18105 4479 18139
rect 4479 18105 4488 18139
rect 4436 18096 4488 18105
rect 5356 18164 5408 18216
rect 6092 18164 6144 18216
rect 6184 18207 6236 18216
rect 6184 18173 6193 18207
rect 6193 18173 6227 18207
rect 6227 18173 6236 18207
rect 6184 18164 6236 18173
rect 8392 18232 8444 18284
rect 10324 18343 10376 18352
rect 10324 18309 10333 18343
rect 10333 18309 10367 18343
rect 10367 18309 10376 18343
rect 10324 18300 10376 18309
rect 11428 18300 11480 18352
rect 11796 18343 11848 18352
rect 11796 18309 11805 18343
rect 11805 18309 11839 18343
rect 11839 18309 11848 18343
rect 11796 18300 11848 18309
rect 15844 18368 15896 18420
rect 17040 18411 17092 18420
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 17224 18368 17276 18420
rect 17500 18368 17552 18420
rect 12624 18300 12676 18352
rect 7472 18096 7524 18148
rect 7748 18096 7800 18148
rect 9956 18164 10008 18216
rect 10324 18164 10376 18216
rect 10692 18164 10744 18216
rect 8576 18096 8628 18148
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 4804 18028 4856 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 6000 18028 6052 18080
rect 7196 18028 7248 18080
rect 7840 18028 7892 18080
rect 11428 18207 11480 18216
rect 11428 18173 11437 18207
rect 11437 18173 11471 18207
rect 11471 18173 11480 18207
rect 11428 18164 11480 18173
rect 11612 18207 11664 18216
rect 11612 18173 11621 18207
rect 11621 18173 11655 18207
rect 11655 18173 11664 18207
rect 11612 18164 11664 18173
rect 11796 18164 11848 18216
rect 12992 18300 13044 18352
rect 15108 18300 15160 18352
rect 15200 18300 15252 18352
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 20444 18411 20496 18420
rect 20444 18377 20453 18411
rect 20453 18377 20487 18411
rect 20487 18377 20496 18411
rect 20444 18368 20496 18377
rect 20720 18368 20772 18420
rect 22376 18368 22428 18420
rect 24124 18368 24176 18420
rect 24492 18368 24544 18420
rect 24860 18368 24912 18420
rect 26148 18368 26200 18420
rect 26700 18368 26752 18420
rect 29276 18368 29328 18420
rect 29552 18368 29604 18420
rect 30196 18368 30248 18420
rect 30472 18368 30524 18420
rect 12348 18096 12400 18148
rect 13268 18164 13320 18216
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 13912 18164 13964 18173
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 15016 18164 15068 18216
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 15476 18207 15528 18216
rect 15476 18173 15485 18207
rect 15485 18173 15519 18207
rect 15519 18173 15528 18207
rect 15476 18164 15528 18173
rect 15660 18164 15712 18216
rect 16120 18232 16172 18284
rect 16028 18207 16080 18216
rect 16028 18173 16037 18207
rect 16037 18173 16071 18207
rect 16071 18173 16080 18207
rect 16028 18164 16080 18173
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 16948 18164 17000 18216
rect 17224 18164 17276 18216
rect 17868 18164 17920 18216
rect 18696 18164 18748 18216
rect 18972 18232 19024 18284
rect 19064 18207 19116 18216
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 20260 18300 20312 18352
rect 20628 18300 20680 18352
rect 20812 18343 20864 18352
rect 20812 18309 20821 18343
rect 20821 18309 20855 18343
rect 20855 18309 20864 18343
rect 20812 18300 20864 18309
rect 21272 18300 21324 18352
rect 22468 18300 22520 18352
rect 19708 18207 19760 18216
rect 9680 18028 9732 18080
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 10600 18028 10652 18080
rect 10968 18028 11020 18080
rect 11980 18028 12032 18080
rect 13452 18028 13504 18080
rect 16764 18096 16816 18148
rect 17684 18096 17736 18148
rect 16028 18028 16080 18080
rect 16488 18028 16540 18080
rect 16580 18028 16632 18080
rect 17224 18028 17276 18080
rect 17592 18028 17644 18080
rect 18512 18028 18564 18080
rect 19156 18028 19208 18080
rect 19340 18096 19392 18148
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 19708 18164 19760 18173
rect 20076 18096 20128 18148
rect 23020 18300 23072 18352
rect 25872 18300 25924 18352
rect 26240 18300 26292 18352
rect 22744 18275 22796 18284
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 23112 18232 23164 18284
rect 24308 18232 24360 18284
rect 24492 18232 24544 18284
rect 27252 18232 27304 18284
rect 27344 18232 27396 18284
rect 22836 18164 22888 18216
rect 23020 18207 23072 18216
rect 23020 18173 23029 18207
rect 23029 18173 23063 18207
rect 23063 18173 23072 18207
rect 23020 18164 23072 18173
rect 23480 18164 23532 18216
rect 23756 18164 23808 18216
rect 24032 18164 24084 18216
rect 24860 18164 24912 18216
rect 24676 18096 24728 18148
rect 20996 18028 21048 18080
rect 21916 18028 21968 18080
rect 25412 18096 25464 18148
rect 25688 18096 25740 18148
rect 25872 18096 25924 18148
rect 26976 18096 27028 18148
rect 25228 18028 25280 18080
rect 28080 18300 28132 18352
rect 28632 18164 28684 18216
rect 30104 18164 30156 18216
rect 30656 18207 30708 18216
rect 30656 18173 30665 18207
rect 30665 18173 30699 18207
rect 30699 18173 30708 18207
rect 30656 18164 30708 18173
rect 27804 18096 27856 18148
rect 30012 18096 30064 18148
rect 30472 18028 30524 18080
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 15946 17926 15998 17978
rect 16010 17926 16062 17978
rect 16074 17926 16126 17978
rect 16138 17926 16190 17978
rect 16202 17926 16254 17978
rect 23720 17926 23772 17978
rect 23784 17926 23836 17978
rect 23848 17926 23900 17978
rect 23912 17926 23964 17978
rect 23976 17926 24028 17978
rect 31494 17926 31546 17978
rect 31558 17926 31610 17978
rect 31622 17926 31674 17978
rect 31686 17926 31738 17978
rect 31750 17926 31802 17978
rect 2596 17756 2648 17808
rect 2780 17824 2832 17876
rect 3792 17824 3844 17876
rect 3976 17824 4028 17876
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 5816 17824 5868 17876
rect 4528 17756 4580 17808
rect 4436 17688 4488 17740
rect 5632 17756 5684 17808
rect 6828 17824 6880 17876
rect 7748 17824 7800 17876
rect 8024 17824 8076 17876
rect 7196 17756 7248 17808
rect 8300 17756 8352 17808
rect 8668 17824 8720 17876
rect 9036 17824 9088 17876
rect 1124 17663 1176 17672
rect 1124 17629 1133 17663
rect 1133 17629 1167 17663
rect 1167 17629 1176 17663
rect 1124 17620 1176 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3976 17620 4028 17672
rect 5448 17620 5500 17672
rect 6460 17620 6512 17672
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 7104 17620 7156 17672
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 3056 17484 3108 17536
rect 3700 17484 3752 17536
rect 4712 17484 4764 17536
rect 4896 17484 4948 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6736 17484 6788 17536
rect 7840 17484 7892 17536
rect 8208 17527 8260 17536
rect 8208 17493 8217 17527
rect 8217 17493 8251 17527
rect 8251 17493 8260 17527
rect 8208 17484 8260 17493
rect 8760 17731 8812 17740
rect 8760 17697 8769 17731
rect 8769 17697 8803 17731
rect 8803 17697 8812 17731
rect 8760 17688 8812 17697
rect 9404 17756 9456 17808
rect 9220 17731 9272 17740
rect 9220 17697 9229 17731
rect 9229 17697 9263 17731
rect 9263 17697 9272 17731
rect 9220 17688 9272 17697
rect 9588 17731 9640 17740
rect 9588 17697 9597 17731
rect 9597 17697 9631 17731
rect 9631 17697 9640 17731
rect 9588 17688 9640 17697
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 9864 17756 9916 17808
rect 10416 17824 10468 17876
rect 10600 17824 10652 17876
rect 10140 17731 10192 17740
rect 10140 17697 10144 17731
rect 10144 17697 10178 17731
rect 10178 17697 10192 17731
rect 10140 17688 10192 17697
rect 10968 17756 11020 17808
rect 12348 17867 12400 17876
rect 12348 17833 12350 17867
rect 12350 17833 12384 17867
rect 12384 17833 12400 17867
rect 12348 17824 12400 17833
rect 11428 17756 11480 17808
rect 10508 17731 10560 17740
rect 10508 17697 10516 17731
rect 10516 17697 10550 17731
rect 10550 17697 10560 17731
rect 10508 17688 10560 17697
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 10784 17688 10836 17740
rect 11796 17731 11848 17740
rect 11796 17697 11805 17731
rect 11805 17697 11839 17731
rect 11839 17697 11848 17731
rect 11796 17688 11848 17697
rect 11980 17688 12032 17740
rect 12624 17756 12676 17808
rect 16580 17824 16632 17876
rect 16948 17867 17000 17876
rect 16948 17833 16957 17867
rect 16957 17833 16991 17867
rect 16991 17833 17000 17867
rect 16948 17824 17000 17833
rect 17776 17824 17828 17876
rect 18512 17824 18564 17876
rect 18696 17824 18748 17876
rect 8484 17552 8536 17604
rect 9496 17552 9548 17604
rect 8668 17484 8720 17536
rect 10232 17552 10284 17604
rect 10692 17552 10744 17604
rect 10876 17484 10928 17536
rect 11244 17552 11296 17604
rect 11980 17484 12032 17536
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13544 17688 13596 17740
rect 13636 17688 13688 17740
rect 16672 17688 16724 17740
rect 18972 17756 19024 17808
rect 12808 17620 12860 17672
rect 13360 17620 13412 17672
rect 16212 17620 16264 17672
rect 17316 17688 17368 17740
rect 17500 17688 17552 17740
rect 17868 17688 17920 17740
rect 18880 17688 18932 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 19432 17799 19484 17808
rect 19432 17765 19441 17799
rect 19441 17765 19475 17799
rect 19475 17765 19484 17799
rect 19432 17756 19484 17765
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 21548 17824 21600 17876
rect 23296 17824 23348 17876
rect 23480 17824 23532 17876
rect 20168 17799 20220 17808
rect 20168 17765 20177 17799
rect 20177 17765 20211 17799
rect 20211 17765 20220 17799
rect 20168 17756 20220 17765
rect 20812 17756 20864 17808
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 19800 17688 19852 17740
rect 14004 17552 14056 17604
rect 14096 17484 14148 17536
rect 15200 17484 15252 17536
rect 17500 17552 17552 17604
rect 18236 17552 18288 17604
rect 19432 17620 19484 17672
rect 19340 17552 19392 17604
rect 20536 17620 20588 17672
rect 20720 17688 20772 17740
rect 21640 17799 21692 17808
rect 21640 17765 21649 17799
rect 21649 17765 21683 17799
rect 21683 17765 21692 17799
rect 21640 17756 21692 17765
rect 23204 17756 23256 17808
rect 23572 17756 23624 17808
rect 20812 17620 20864 17672
rect 20996 17620 21048 17672
rect 21824 17731 21876 17740
rect 21824 17697 21833 17731
rect 21833 17697 21867 17731
rect 21867 17697 21876 17731
rect 21824 17688 21876 17697
rect 25044 17824 25096 17876
rect 27068 17824 27120 17876
rect 28080 17824 28132 17876
rect 26056 17756 26108 17808
rect 28448 17756 28500 17808
rect 28908 17867 28960 17876
rect 28908 17833 28917 17867
rect 28917 17833 28951 17867
rect 28951 17833 28960 17867
rect 28908 17824 28960 17833
rect 29920 17867 29972 17876
rect 29920 17833 29929 17867
rect 29929 17833 29963 17867
rect 29963 17833 29972 17867
rect 29920 17824 29972 17833
rect 29184 17756 29236 17808
rect 24492 17731 24544 17740
rect 24492 17697 24501 17731
rect 24501 17697 24535 17731
rect 24535 17697 24544 17731
rect 24492 17688 24544 17697
rect 24308 17620 24360 17672
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 25320 17688 25372 17740
rect 25780 17688 25832 17740
rect 26424 17688 26476 17740
rect 26516 17688 26568 17740
rect 26608 17731 26660 17740
rect 26608 17697 26617 17731
rect 26617 17697 26651 17731
rect 26651 17697 26660 17731
rect 26608 17688 26660 17697
rect 19156 17484 19208 17536
rect 22928 17552 22980 17604
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 22284 17484 22336 17536
rect 23940 17527 23992 17536
rect 23940 17493 23949 17527
rect 23949 17493 23983 17527
rect 23983 17493 23992 17527
rect 23940 17484 23992 17493
rect 24860 17484 24912 17536
rect 25780 17595 25832 17604
rect 25780 17561 25789 17595
rect 25789 17561 25823 17595
rect 25823 17561 25832 17595
rect 25780 17552 25832 17561
rect 28356 17731 28408 17740
rect 28356 17697 28365 17731
rect 28365 17697 28399 17731
rect 28399 17697 28408 17731
rect 28356 17688 28408 17697
rect 28724 17731 28776 17740
rect 28724 17697 28733 17731
rect 28733 17697 28767 17731
rect 28767 17697 28776 17731
rect 28724 17688 28776 17697
rect 28540 17620 28592 17672
rect 28632 17552 28684 17604
rect 26516 17484 26568 17536
rect 26976 17484 27028 17536
rect 30196 17731 30248 17740
rect 30196 17697 30205 17731
rect 30205 17697 30239 17731
rect 30239 17697 30248 17731
rect 30196 17688 30248 17697
rect 30288 17552 30340 17604
rect 30472 17688 30524 17740
rect 29460 17484 29512 17536
rect 4285 17382 4337 17434
rect 4349 17382 4401 17434
rect 4413 17382 4465 17434
rect 4477 17382 4529 17434
rect 4541 17382 4593 17434
rect 12059 17382 12111 17434
rect 12123 17382 12175 17434
rect 12187 17382 12239 17434
rect 12251 17382 12303 17434
rect 12315 17382 12367 17434
rect 19833 17382 19885 17434
rect 19897 17382 19949 17434
rect 19961 17382 20013 17434
rect 20025 17382 20077 17434
rect 20089 17382 20141 17434
rect 27607 17382 27659 17434
rect 27671 17382 27723 17434
rect 27735 17382 27787 17434
rect 27799 17382 27851 17434
rect 27863 17382 27915 17434
rect 1124 17280 1176 17332
rect 2964 17280 3016 17332
rect 3424 17280 3476 17332
rect 2872 17212 2924 17264
rect 4712 17212 4764 17264
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 5632 17280 5684 17332
rect 5908 17280 5960 17332
rect 8116 17323 8168 17332
rect 8116 17289 8125 17323
rect 8125 17289 8159 17323
rect 8159 17289 8168 17323
rect 8116 17280 8168 17289
rect 8208 17280 8260 17332
rect 8760 17323 8812 17332
rect 8760 17289 8769 17323
rect 8769 17289 8803 17323
rect 8803 17289 8812 17323
rect 8760 17280 8812 17289
rect 8944 17280 8996 17332
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 10140 17280 10192 17332
rect 10416 17280 10468 17332
rect 11060 17280 11112 17332
rect 11244 17280 11296 17332
rect 13912 17280 13964 17332
rect 14740 17280 14792 17332
rect 15476 17280 15528 17332
rect 15844 17280 15896 17332
rect 16948 17280 17000 17332
rect 17684 17280 17736 17332
rect 17868 17280 17920 17332
rect 18328 17280 18380 17332
rect 19248 17323 19300 17332
rect 19248 17289 19257 17323
rect 19257 17289 19291 17323
rect 19291 17289 19300 17323
rect 19248 17280 19300 17289
rect 19892 17280 19944 17332
rect 20996 17280 21048 17332
rect 2872 17076 2924 17128
rect 2964 17008 3016 17060
rect 2504 16940 2556 16992
rect 4160 17076 4212 17128
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 5172 17076 5224 17128
rect 6184 17144 6236 17196
rect 7656 17144 7708 17196
rect 6920 17076 6972 17128
rect 4528 17051 4580 17060
rect 4528 17017 4537 17051
rect 4537 17017 4571 17051
rect 4571 17017 4580 17051
rect 4528 17008 4580 17017
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 3608 16940 3660 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 4160 16940 4212 16992
rect 5632 16940 5684 16992
rect 7932 17076 7984 17128
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 7748 16940 7800 16949
rect 7840 16940 7892 16992
rect 9864 17212 9916 17264
rect 10232 17212 10284 17264
rect 8300 17076 8352 17128
rect 9128 17076 9180 17128
rect 8576 17051 8628 17060
rect 8576 17017 8585 17051
rect 8585 17017 8619 17051
rect 8619 17017 8628 17051
rect 8576 17008 8628 17017
rect 8760 17008 8812 17060
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 9772 17144 9824 17196
rect 9772 17008 9824 17060
rect 9956 17076 10008 17128
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10324 17076 10376 17128
rect 10692 17144 10744 17196
rect 10968 17144 11020 17196
rect 11796 17212 11848 17264
rect 11520 17076 11572 17128
rect 11796 17076 11848 17128
rect 12532 17212 12584 17264
rect 20628 17212 20680 17264
rect 24124 17280 24176 17332
rect 24676 17280 24728 17332
rect 12532 17076 12584 17128
rect 13636 17144 13688 17196
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13912 17144 13964 17196
rect 13176 17076 13228 17085
rect 14556 17076 14608 17128
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 15200 17076 15252 17128
rect 15292 17076 15344 17128
rect 16304 17144 16356 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 19708 17144 19760 17196
rect 20260 17144 20312 17196
rect 10784 17008 10836 17060
rect 10968 17051 11020 17060
rect 10968 17017 10977 17051
rect 10977 17017 11011 17051
rect 11011 17017 11020 17051
rect 10968 17008 11020 17017
rect 11980 17051 12032 17060
rect 11980 17017 11989 17051
rect 11989 17017 12023 17051
rect 12023 17017 12032 17051
rect 11980 17008 12032 17017
rect 12808 17051 12860 17060
rect 12808 17017 12817 17051
rect 12817 17017 12851 17051
rect 12851 17017 12860 17051
rect 12808 17008 12860 17017
rect 11060 16940 11112 16992
rect 11428 16940 11480 16992
rect 11612 16940 11664 16992
rect 12164 16940 12216 16992
rect 12716 16940 12768 16992
rect 13176 16940 13228 16992
rect 15016 17008 15068 17060
rect 15752 17119 15804 17128
rect 15752 17085 15764 17119
rect 15764 17085 15798 17119
rect 15798 17085 15804 17119
rect 15752 17076 15804 17085
rect 16396 17076 16448 17128
rect 17132 17076 17184 17128
rect 16488 17008 16540 17060
rect 13452 16940 13504 16992
rect 17224 16940 17276 16992
rect 17408 17008 17460 17060
rect 17960 17076 18012 17128
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 17960 16940 18012 16992
rect 19064 17076 19116 17128
rect 18696 17008 18748 17060
rect 18788 17008 18840 17060
rect 19248 17051 19300 17060
rect 19248 17017 19275 17051
rect 19275 17017 19300 17051
rect 19248 17008 19300 17017
rect 20536 17076 20588 17128
rect 20812 17119 20864 17128
rect 20812 17085 20821 17119
rect 20821 17085 20855 17119
rect 20855 17085 20864 17119
rect 20812 17076 20864 17085
rect 18512 16940 18564 16992
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 22376 17212 22428 17264
rect 23480 17212 23532 17264
rect 23756 17212 23808 17264
rect 24216 17212 24268 17264
rect 25320 17255 25372 17264
rect 25320 17221 25329 17255
rect 25329 17221 25363 17255
rect 25363 17221 25372 17255
rect 25320 17212 25372 17221
rect 25504 17212 25556 17264
rect 27160 17280 27212 17332
rect 27988 17280 28040 17332
rect 30656 17280 30708 17332
rect 28264 17212 28316 17264
rect 29184 17212 29236 17264
rect 21088 17051 21140 17060
rect 21088 17017 21097 17051
rect 21097 17017 21131 17051
rect 21131 17017 21140 17051
rect 21088 17008 21140 17017
rect 21272 17051 21324 17060
rect 21272 17017 21281 17051
rect 21281 17017 21315 17051
rect 21315 17017 21324 17051
rect 21272 17008 21324 17017
rect 22008 17076 22060 17128
rect 23572 17144 23624 17196
rect 23940 17144 23992 17196
rect 26240 17144 26292 17196
rect 26608 17144 26660 17196
rect 22284 17076 22336 17128
rect 22928 17076 22980 17128
rect 26976 17144 27028 17196
rect 21364 16983 21416 16992
rect 21364 16949 21373 16983
rect 21373 16949 21407 16983
rect 21407 16949 21416 16983
rect 21364 16940 21416 16949
rect 21640 16940 21692 16992
rect 23756 17008 23808 17060
rect 26884 17119 26936 17128
rect 26884 17085 26893 17119
rect 26893 17085 26927 17119
rect 26927 17085 26936 17119
rect 26884 17076 26936 17085
rect 27068 17076 27120 17128
rect 26976 17008 27028 17060
rect 27160 17008 27212 17060
rect 27252 17008 27304 17060
rect 27436 17076 27488 17128
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 28632 17144 28684 17196
rect 28908 17144 28960 17196
rect 29092 17144 29144 17196
rect 29368 17076 29420 17128
rect 30840 17212 30892 17264
rect 30472 17144 30524 17196
rect 28356 17008 28408 17060
rect 30380 17051 30432 17060
rect 30380 17017 30389 17051
rect 30389 17017 30423 17051
rect 30423 17017 30432 17051
rect 30380 17008 30432 17017
rect 23112 16940 23164 16992
rect 25320 16940 25372 16992
rect 26424 16940 26476 16992
rect 27068 16940 27120 16992
rect 30196 16940 30248 16992
rect 30564 16940 30616 16992
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 15946 16838 15998 16890
rect 16010 16838 16062 16890
rect 16074 16838 16126 16890
rect 16138 16838 16190 16890
rect 16202 16838 16254 16890
rect 23720 16838 23772 16890
rect 23784 16838 23836 16890
rect 23848 16838 23900 16890
rect 23912 16838 23964 16890
rect 23976 16838 24028 16890
rect 31494 16838 31546 16890
rect 31558 16838 31610 16890
rect 31622 16838 31674 16890
rect 31686 16838 31738 16890
rect 31750 16838 31802 16890
rect 2780 16600 2832 16652
rect 3700 16736 3752 16788
rect 5172 16736 5224 16788
rect 4712 16600 4764 16652
rect 5632 16668 5684 16720
rect 1124 16575 1176 16584
rect 1124 16541 1133 16575
rect 1133 16541 1167 16575
rect 1167 16541 1176 16575
rect 1124 16532 1176 16541
rect 3424 16532 3476 16584
rect 3792 16532 3844 16584
rect 7748 16736 7800 16788
rect 8576 16736 8628 16788
rect 9588 16736 9640 16788
rect 9772 16736 9824 16788
rect 10048 16736 10100 16788
rect 7380 16668 7432 16720
rect 10600 16736 10652 16788
rect 5264 16464 5316 16516
rect 7104 16532 7156 16584
rect 7840 16600 7892 16652
rect 8760 16532 8812 16584
rect 8944 16532 8996 16584
rect 9312 16532 9364 16584
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 3792 16396 3844 16448
rect 3884 16396 3936 16448
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 5172 16396 5224 16448
rect 5356 16396 5408 16448
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9404 16396 9456 16448
rect 9956 16600 10008 16652
rect 10324 16643 10376 16652
rect 10324 16609 10328 16643
rect 10328 16609 10362 16643
rect 10362 16609 10376 16643
rect 10324 16600 10376 16609
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 10600 16643 10652 16652
rect 11428 16668 11480 16720
rect 10600 16609 10645 16643
rect 10645 16609 10652 16643
rect 10600 16600 10652 16609
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 11060 16600 11112 16652
rect 11888 16668 11940 16720
rect 12164 16668 12216 16720
rect 13084 16736 13136 16788
rect 14464 16736 14516 16788
rect 15568 16736 15620 16788
rect 12072 16643 12124 16652
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 13912 16668 13964 16720
rect 13360 16600 13412 16652
rect 12624 16532 12676 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 10232 16464 10284 16516
rect 10968 16464 11020 16516
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 13176 16396 13228 16448
rect 13360 16464 13412 16516
rect 14372 16600 14424 16652
rect 14648 16600 14700 16652
rect 14740 16600 14792 16652
rect 14924 16600 14976 16652
rect 18420 16736 18472 16788
rect 20628 16736 20680 16788
rect 21272 16736 21324 16788
rect 21640 16736 21692 16788
rect 16580 16711 16632 16720
rect 16580 16677 16589 16711
rect 16589 16677 16623 16711
rect 16623 16677 16632 16711
rect 16580 16668 16632 16677
rect 16396 16600 16448 16652
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17500 16600 17552 16652
rect 17868 16668 17920 16720
rect 14464 16464 14516 16516
rect 14096 16396 14148 16448
rect 14372 16396 14424 16448
rect 14740 16507 14792 16516
rect 14740 16473 14749 16507
rect 14749 16473 14783 16507
rect 14783 16473 14792 16507
rect 14740 16464 14792 16473
rect 14924 16464 14976 16516
rect 16304 16464 16356 16516
rect 16856 16532 16908 16584
rect 18604 16532 18656 16584
rect 19708 16600 19760 16652
rect 18052 16464 18104 16516
rect 19156 16464 19208 16516
rect 19432 16464 19484 16516
rect 19708 16464 19760 16516
rect 19892 16643 19944 16652
rect 19892 16609 19901 16643
rect 19901 16609 19935 16643
rect 19935 16609 19944 16643
rect 19892 16600 19944 16609
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 20536 16600 20588 16652
rect 20904 16600 20956 16652
rect 21548 16600 21600 16652
rect 22284 16668 22336 16720
rect 22744 16668 22796 16720
rect 22560 16600 22612 16652
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 23296 16600 23348 16652
rect 24216 16668 24268 16720
rect 24308 16668 24360 16720
rect 24400 16711 24452 16720
rect 24400 16677 24409 16711
rect 24409 16677 24443 16711
rect 24443 16677 24452 16711
rect 24400 16668 24452 16677
rect 24676 16736 24728 16788
rect 25780 16736 25832 16788
rect 26608 16736 26660 16788
rect 26976 16736 27028 16788
rect 27160 16779 27212 16788
rect 27160 16745 27169 16779
rect 27169 16745 27203 16779
rect 27203 16745 27212 16779
rect 27160 16736 27212 16745
rect 27436 16736 27488 16788
rect 30564 16736 30616 16788
rect 25044 16668 25096 16720
rect 25228 16668 25280 16720
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 21364 16532 21416 16584
rect 26240 16600 26292 16652
rect 20168 16464 20220 16516
rect 20720 16464 20772 16516
rect 22928 16464 22980 16516
rect 23572 16464 23624 16516
rect 16764 16396 16816 16448
rect 16948 16396 17000 16448
rect 17132 16396 17184 16448
rect 17408 16439 17460 16448
rect 17408 16405 17417 16439
rect 17417 16405 17451 16439
rect 17451 16405 17460 16439
rect 17408 16396 17460 16405
rect 17960 16396 18012 16448
rect 18604 16396 18656 16448
rect 19616 16396 19668 16448
rect 21272 16396 21324 16448
rect 22192 16396 22244 16448
rect 22744 16396 22796 16448
rect 22836 16439 22888 16448
rect 22836 16405 22845 16439
rect 22845 16405 22879 16439
rect 22879 16405 22888 16439
rect 22836 16396 22888 16405
rect 24584 16396 24636 16448
rect 25228 16396 25280 16448
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 26976 16600 27028 16652
rect 27252 16600 27304 16652
rect 25504 16507 25556 16516
rect 25504 16473 25513 16507
rect 25513 16473 25547 16507
rect 25547 16473 25556 16507
rect 25504 16464 25556 16473
rect 25780 16464 25832 16516
rect 26976 16464 27028 16516
rect 27160 16464 27212 16516
rect 27620 16464 27672 16516
rect 28264 16600 28316 16652
rect 28540 16600 28592 16652
rect 28816 16507 28868 16516
rect 28816 16473 28825 16507
rect 28825 16473 28859 16507
rect 28859 16473 28868 16507
rect 28816 16464 28868 16473
rect 28908 16507 28960 16516
rect 28908 16473 28917 16507
rect 28917 16473 28951 16507
rect 28951 16473 28960 16507
rect 28908 16464 28960 16473
rect 28356 16396 28408 16448
rect 29184 16600 29236 16652
rect 29368 16643 29420 16652
rect 29368 16609 29377 16643
rect 29377 16609 29411 16643
rect 29411 16609 29420 16643
rect 29368 16600 29420 16609
rect 29552 16643 29604 16652
rect 29552 16609 29561 16643
rect 29561 16609 29595 16643
rect 29595 16609 29604 16643
rect 29552 16600 29604 16609
rect 30380 16600 30432 16652
rect 30656 16600 30708 16652
rect 29276 16396 29328 16448
rect 4285 16294 4337 16346
rect 4349 16294 4401 16346
rect 4413 16294 4465 16346
rect 4477 16294 4529 16346
rect 4541 16294 4593 16346
rect 12059 16294 12111 16346
rect 12123 16294 12175 16346
rect 12187 16294 12239 16346
rect 12251 16294 12303 16346
rect 12315 16294 12367 16346
rect 19833 16294 19885 16346
rect 19897 16294 19949 16346
rect 19961 16294 20013 16346
rect 20025 16294 20077 16346
rect 20089 16294 20141 16346
rect 27607 16294 27659 16346
rect 27671 16294 27723 16346
rect 27735 16294 27787 16346
rect 27799 16294 27851 16346
rect 27863 16294 27915 16346
rect 1124 16192 1176 16244
rect 1032 16124 1084 16176
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 4068 16124 4120 16176
rect 2136 16056 2188 16065
rect 3148 16056 3200 16108
rect 2596 15988 2648 16040
rect 2872 15988 2924 16040
rect 3608 15988 3660 16040
rect 4988 16056 5040 16108
rect 5172 16099 5224 16108
rect 5172 16065 5181 16099
rect 5181 16065 5215 16099
rect 5215 16065 5224 16099
rect 5172 16056 5224 16065
rect 5540 16056 5592 16108
rect 7288 16056 7340 16108
rect 7748 16056 7800 16108
rect 8760 16192 8812 16244
rect 8668 16124 8720 16176
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 9404 16192 9456 16244
rect 9680 16192 9732 16244
rect 9864 16192 9916 16244
rect 10876 16192 10928 16244
rect 11336 16192 11388 16244
rect 11980 16192 12032 16244
rect 13360 16192 13412 16244
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 7380 15988 7432 16040
rect 11060 16056 11112 16108
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 8484 15988 8536 16040
rect 9312 15988 9364 16040
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 11888 16056 11940 16108
rect 12808 16124 12860 16176
rect 14004 16124 14056 16176
rect 12992 16056 13044 16108
rect 13636 16056 13688 16108
rect 5632 15920 5684 15972
rect 6092 15963 6144 15972
rect 6092 15929 6101 15963
rect 6101 15929 6135 15963
rect 6135 15929 6144 15963
rect 6092 15920 6144 15929
rect 3240 15852 3292 15904
rect 3332 15895 3384 15904
rect 3332 15861 3341 15895
rect 3341 15861 3375 15895
rect 3375 15861 3384 15895
rect 3332 15852 3384 15861
rect 4620 15852 4672 15904
rect 5172 15852 5224 15904
rect 8576 15852 8628 15904
rect 8944 15852 8996 15904
rect 9404 15963 9456 15972
rect 9404 15929 9413 15963
rect 9413 15929 9447 15963
rect 9447 15929 9456 15963
rect 9404 15920 9456 15929
rect 9956 15920 10008 15972
rect 11244 15852 11296 15904
rect 14372 15920 14424 15972
rect 14556 16192 14608 16244
rect 14924 16192 14976 16244
rect 16304 16192 16356 16244
rect 17316 16192 17368 16244
rect 15384 16124 15436 16176
rect 16396 16124 16448 16176
rect 16764 16124 16816 16176
rect 17408 16124 17460 16176
rect 17960 16124 18012 16176
rect 18144 16124 18196 16176
rect 18696 16124 18748 16176
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 15752 16056 15804 16108
rect 15292 15988 15344 16040
rect 17316 15988 17368 16040
rect 17408 16031 17460 16040
rect 17408 15997 17417 16031
rect 17417 15997 17451 16031
rect 17451 15997 17460 16031
rect 17408 15988 17460 15997
rect 17500 16031 17552 16040
rect 17500 15997 17509 16031
rect 17509 15997 17543 16031
rect 17543 15997 17552 16031
rect 17500 15988 17552 15997
rect 17776 15988 17828 16040
rect 17960 15988 18012 16040
rect 18604 15988 18656 16040
rect 18972 16192 19024 16244
rect 19248 16192 19300 16244
rect 20904 16192 20956 16244
rect 21824 16192 21876 16244
rect 21916 16192 21968 16244
rect 23020 16192 23072 16244
rect 23112 16192 23164 16244
rect 23388 16192 23440 16244
rect 24216 16235 24268 16244
rect 24216 16201 24225 16235
rect 24225 16201 24259 16235
rect 24259 16201 24268 16235
rect 24216 16192 24268 16201
rect 24400 16192 24452 16244
rect 25780 16192 25832 16244
rect 26056 16192 26108 16244
rect 29368 16192 29420 16244
rect 29644 16192 29696 16244
rect 30196 16235 30248 16244
rect 30196 16201 30205 16235
rect 30205 16201 30239 16235
rect 30239 16201 30248 16235
rect 30196 16192 30248 16201
rect 19248 16056 19300 16108
rect 18328 15920 18380 15972
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 13084 15852 13136 15904
rect 13452 15852 13504 15904
rect 17592 15852 17644 15904
rect 19432 15920 19484 15972
rect 19616 15920 19668 15972
rect 18880 15852 18932 15904
rect 20168 15920 20220 15972
rect 20352 15920 20404 15972
rect 20628 16031 20680 16040
rect 20628 15997 20637 16031
rect 20637 15997 20671 16031
rect 20671 15997 20680 16031
rect 20628 15988 20680 15997
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 20996 16056 21048 16108
rect 21180 16056 21232 16108
rect 21272 16099 21324 16108
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 20996 15852 21048 15904
rect 21916 15988 21968 16040
rect 27068 16167 27120 16176
rect 27068 16133 27077 16167
rect 27077 16133 27111 16167
rect 27111 16133 27120 16167
rect 27068 16124 27120 16133
rect 22836 16056 22888 16108
rect 22928 16031 22980 16040
rect 22928 15997 22949 16031
rect 22949 15997 22980 16031
rect 25688 16056 25740 16108
rect 25780 16056 25832 16108
rect 28632 16124 28684 16176
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 28172 16056 28224 16108
rect 30196 16056 30248 16108
rect 22928 15988 22980 15997
rect 23572 15988 23624 16040
rect 21180 15963 21232 15972
rect 21180 15929 21189 15963
rect 21189 15929 21223 15963
rect 21223 15929 21232 15963
rect 21180 15920 21232 15929
rect 21548 15920 21600 15972
rect 21272 15852 21324 15904
rect 23296 15852 23348 15904
rect 23940 15920 23992 15972
rect 28724 15988 28776 16040
rect 30380 16031 30432 16040
rect 30380 15997 30389 16031
rect 30389 15997 30423 16031
rect 30423 15997 30432 16031
rect 30380 15988 30432 15997
rect 26700 15920 26752 15972
rect 27436 15920 27488 15972
rect 29736 15920 29788 15972
rect 30748 15988 30800 16040
rect 24400 15852 24452 15904
rect 27528 15895 27580 15904
rect 27528 15861 27537 15895
rect 27537 15861 27571 15895
rect 27571 15861 27580 15895
rect 27528 15852 27580 15861
rect 30472 15852 30524 15904
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 15946 15750 15998 15802
rect 16010 15750 16062 15802
rect 16074 15750 16126 15802
rect 16138 15750 16190 15802
rect 16202 15750 16254 15802
rect 23720 15750 23772 15802
rect 23784 15750 23836 15802
rect 23848 15750 23900 15802
rect 23912 15750 23964 15802
rect 23976 15750 24028 15802
rect 31494 15750 31546 15802
rect 31558 15750 31610 15802
rect 31622 15750 31674 15802
rect 31686 15750 31738 15802
rect 31750 15750 31802 15802
rect 1032 15648 1084 15700
rect 2780 15580 2832 15632
rect 5356 15648 5408 15700
rect 6092 15648 6144 15700
rect 6184 15648 6236 15700
rect 6644 15648 6696 15700
rect 3332 15512 3384 15564
rect 4804 15512 4856 15564
rect 2688 15444 2740 15496
rect 3792 15444 3844 15496
rect 4068 15444 4120 15496
rect 940 15308 992 15360
rect 2872 15308 2924 15360
rect 4988 15308 5040 15360
rect 9312 15648 9364 15700
rect 9404 15648 9456 15700
rect 9496 15648 9548 15700
rect 9588 15648 9640 15700
rect 11060 15648 11112 15700
rect 11704 15648 11756 15700
rect 12532 15691 12584 15700
rect 12532 15657 12541 15691
rect 12541 15657 12575 15691
rect 12575 15657 12584 15691
rect 12532 15648 12584 15657
rect 12716 15648 12768 15700
rect 14188 15648 14240 15700
rect 14372 15648 14424 15700
rect 16304 15648 16356 15700
rect 16488 15648 16540 15700
rect 17500 15648 17552 15700
rect 17592 15648 17644 15700
rect 18328 15691 18380 15700
rect 18328 15657 18337 15691
rect 18337 15657 18371 15691
rect 18371 15657 18380 15691
rect 18328 15648 18380 15657
rect 18512 15648 18564 15700
rect 18972 15648 19024 15700
rect 7932 15580 7984 15632
rect 6736 15512 6788 15564
rect 6828 15512 6880 15564
rect 7012 15512 7064 15564
rect 8024 15512 8076 15564
rect 8484 15512 8536 15564
rect 9128 15512 9180 15564
rect 9956 15580 10008 15632
rect 10876 15580 10928 15632
rect 11796 15580 11848 15632
rect 9312 15376 9364 15428
rect 9404 15376 9456 15428
rect 9772 15444 9824 15496
rect 9864 15376 9916 15428
rect 8668 15308 8720 15360
rect 11152 15555 11204 15564
rect 11152 15521 11161 15555
rect 11161 15521 11195 15555
rect 11195 15521 11204 15555
rect 11152 15512 11204 15521
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 12716 15555 12768 15564
rect 11612 15512 11664 15521
rect 12716 15521 12728 15555
rect 12728 15521 12762 15555
rect 12762 15521 12768 15555
rect 12716 15512 12768 15521
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 14648 15512 14700 15564
rect 14832 15512 14884 15564
rect 16212 15580 16264 15632
rect 16028 15512 16080 15564
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 10784 15444 10836 15496
rect 10508 15376 10560 15428
rect 11060 15376 11112 15428
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 11888 15376 11940 15428
rect 11980 15376 12032 15428
rect 10692 15308 10744 15360
rect 12992 15308 13044 15360
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 16580 15555 16632 15564
rect 16580 15521 16589 15555
rect 16589 15521 16623 15555
rect 16623 15521 16632 15555
rect 16580 15512 16632 15521
rect 16948 15580 17000 15632
rect 17408 15580 17460 15632
rect 18880 15623 18932 15632
rect 18880 15589 18889 15623
rect 18889 15589 18923 15623
rect 18923 15589 18932 15623
rect 18880 15580 18932 15589
rect 19432 15648 19484 15700
rect 22560 15691 22612 15700
rect 22560 15657 22569 15691
rect 22569 15657 22603 15691
rect 22603 15657 22612 15691
rect 22560 15648 22612 15657
rect 23204 15648 23256 15700
rect 23388 15648 23440 15700
rect 24032 15648 24084 15700
rect 19708 15580 19760 15632
rect 21548 15580 21600 15632
rect 18052 15444 18104 15496
rect 18604 15487 18656 15496
rect 18604 15453 18609 15487
rect 18609 15453 18643 15487
rect 18643 15453 18656 15487
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 15752 15308 15804 15360
rect 16764 15376 16816 15428
rect 17776 15376 17828 15428
rect 18604 15444 18656 15453
rect 18972 15487 19024 15496
rect 18972 15453 18981 15487
rect 18981 15453 19015 15487
rect 19015 15453 19024 15487
rect 18972 15444 19024 15453
rect 19524 15512 19576 15564
rect 20628 15512 20680 15564
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 21364 15512 21416 15564
rect 21456 15512 21508 15564
rect 23020 15580 23072 15632
rect 22192 15555 22244 15564
rect 22192 15521 22201 15555
rect 22201 15521 22235 15555
rect 22235 15521 22244 15555
rect 22192 15512 22244 15521
rect 22744 15555 22796 15564
rect 22744 15521 22753 15555
rect 22753 15521 22787 15555
rect 22787 15521 22796 15555
rect 22744 15512 22796 15521
rect 20444 15444 20496 15496
rect 20536 15444 20588 15496
rect 17592 15308 17644 15360
rect 17868 15308 17920 15360
rect 18328 15308 18380 15360
rect 19248 15308 19300 15360
rect 20812 15376 20864 15428
rect 23204 15512 23256 15564
rect 23756 15580 23808 15632
rect 24308 15648 24360 15700
rect 24676 15648 24728 15700
rect 24860 15648 24912 15700
rect 26148 15648 26200 15700
rect 24216 15623 24268 15632
rect 24216 15589 24225 15623
rect 24225 15589 24259 15623
rect 24259 15589 24268 15623
rect 24216 15580 24268 15589
rect 23940 15555 23992 15564
rect 23940 15521 23950 15555
rect 23950 15521 23984 15555
rect 23984 15521 23992 15555
rect 23940 15512 23992 15521
rect 24400 15512 24452 15564
rect 25044 15512 25096 15564
rect 23480 15444 23532 15496
rect 26424 15580 26476 15632
rect 25228 15444 25280 15496
rect 25412 15444 25464 15496
rect 25688 15487 25740 15496
rect 25688 15453 25697 15487
rect 25697 15453 25731 15487
rect 25731 15453 25740 15487
rect 25688 15444 25740 15453
rect 20076 15308 20128 15360
rect 24216 15376 24268 15428
rect 24584 15376 24636 15428
rect 24676 15376 24728 15428
rect 22560 15308 22612 15360
rect 23572 15308 23624 15360
rect 25320 15308 25372 15360
rect 26148 15512 26200 15564
rect 26792 15555 26844 15564
rect 26792 15521 26801 15555
rect 26801 15521 26835 15555
rect 26835 15521 26844 15555
rect 26792 15512 26844 15521
rect 27528 15648 27580 15700
rect 29552 15648 29604 15700
rect 27712 15623 27764 15632
rect 27712 15589 27721 15623
rect 27721 15589 27755 15623
rect 27755 15589 27764 15623
rect 27712 15580 27764 15589
rect 27436 15555 27488 15564
rect 27436 15521 27445 15555
rect 27445 15521 27479 15555
rect 27479 15521 27488 15555
rect 27436 15512 27488 15521
rect 27528 15512 27580 15564
rect 27988 15512 28040 15564
rect 28264 15512 28316 15564
rect 28632 15512 28684 15564
rect 30380 15580 30432 15632
rect 29368 15555 29420 15564
rect 29368 15521 29377 15555
rect 29377 15521 29411 15555
rect 29411 15521 29420 15555
rect 29368 15512 29420 15521
rect 29644 15555 29696 15564
rect 29644 15521 29653 15555
rect 29653 15521 29687 15555
rect 29687 15521 29696 15555
rect 29644 15512 29696 15521
rect 29736 15512 29788 15564
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 30564 15512 30616 15564
rect 29828 15444 29880 15496
rect 30380 15487 30432 15496
rect 30380 15453 30389 15487
rect 30389 15453 30423 15487
rect 30423 15453 30432 15487
rect 30380 15444 30432 15453
rect 26056 15376 26108 15428
rect 28540 15351 28592 15360
rect 28540 15317 28549 15351
rect 28549 15317 28583 15351
rect 28583 15317 28592 15351
rect 28540 15308 28592 15317
rect 4285 15206 4337 15258
rect 4349 15206 4401 15258
rect 4413 15206 4465 15258
rect 4477 15206 4529 15258
rect 4541 15206 4593 15258
rect 12059 15206 12111 15258
rect 12123 15206 12175 15258
rect 12187 15206 12239 15258
rect 12251 15206 12303 15258
rect 12315 15206 12367 15258
rect 19833 15206 19885 15258
rect 19897 15206 19949 15258
rect 19961 15206 20013 15258
rect 20025 15206 20077 15258
rect 20089 15206 20141 15258
rect 27607 15206 27659 15258
rect 27671 15206 27723 15258
rect 27735 15206 27787 15258
rect 27799 15206 27851 15258
rect 27863 15206 27915 15258
rect 3424 15104 3476 15156
rect 3700 15104 3752 15156
rect 5540 15104 5592 15156
rect 8852 15104 8904 15156
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 756 14968 808 15020
rect 3148 15036 3200 15088
rect 2688 14968 2740 15020
rect 3516 14968 3568 15020
rect 9128 15036 9180 15088
rect 11888 15104 11940 15156
rect 11796 15036 11848 15088
rect 12440 15079 12492 15088
rect 12440 15045 12449 15079
rect 12449 15045 12483 15079
rect 12483 15045 12492 15079
rect 12440 15036 12492 15045
rect 6828 14968 6880 15020
rect 8576 14968 8628 15020
rect 940 14900 992 14952
rect 1216 14943 1268 14952
rect 1216 14909 1225 14943
rect 1225 14909 1259 14943
rect 1259 14909 1268 14943
rect 1216 14900 1268 14909
rect 3608 14900 3660 14952
rect 6920 14900 6972 14952
rect 7380 14900 7432 14952
rect 7932 14900 7984 14952
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 8944 14900 8996 14952
rect 9588 14968 9640 15020
rect 9956 14968 10008 15020
rect 10692 14968 10744 15020
rect 11060 14968 11112 15020
rect 11612 14968 11664 15020
rect 16212 15104 16264 15156
rect 16764 15104 16816 15156
rect 17592 15104 17644 15156
rect 12808 15036 12860 15088
rect 13360 15036 13412 15088
rect 17040 15036 17092 15088
rect 17868 15036 17920 15088
rect 18420 15104 18472 15156
rect 19524 15104 19576 15156
rect 20168 15104 20220 15156
rect 19984 15036 20036 15088
rect 9312 14900 9364 14952
rect 9496 14943 9548 14952
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 2228 14832 2280 14884
rect 2780 14832 2832 14884
rect 4804 14875 4856 14884
rect 4804 14841 4813 14875
rect 4813 14841 4847 14875
rect 4847 14841 4856 14875
rect 4804 14832 4856 14841
rect 2596 14764 2648 14816
rect 3608 14764 3660 14816
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 4252 14764 4304 14816
rect 4620 14764 4672 14816
rect 8024 14832 8076 14884
rect 8484 14832 8536 14884
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 7104 14764 7156 14816
rect 9036 14764 9088 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 12992 14900 13044 14952
rect 15292 15011 15344 15020
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 22560 15104 22612 15156
rect 22744 15104 22796 15156
rect 22836 15147 22888 15156
rect 22836 15113 22845 15147
rect 22845 15113 22879 15147
rect 22879 15113 22888 15147
rect 22836 15104 22888 15113
rect 23020 15104 23072 15156
rect 23480 15104 23532 15156
rect 20444 15036 20496 15088
rect 25412 15036 25464 15088
rect 15292 14968 15344 14977
rect 10600 14832 10652 14884
rect 10876 14832 10928 14884
rect 14280 14900 14332 14952
rect 11888 14764 11940 14816
rect 13912 14764 13964 14816
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 15752 14900 15804 14952
rect 16028 14900 16080 14952
rect 16304 14900 16356 14952
rect 16764 14900 16816 14952
rect 17224 14900 17276 14952
rect 17408 14832 17460 14884
rect 14740 14764 14792 14816
rect 15476 14764 15528 14816
rect 17224 14764 17276 14816
rect 17316 14764 17368 14816
rect 18052 14764 18104 14816
rect 19156 14832 19208 14884
rect 19616 14832 19668 14884
rect 19432 14764 19484 14816
rect 19892 14764 19944 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 20904 14968 20956 15020
rect 21732 14968 21784 15020
rect 22192 14968 22244 15020
rect 20628 14832 20680 14884
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 21180 14900 21232 14952
rect 21640 14900 21692 14952
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 22836 14900 22888 14952
rect 23020 14900 23072 14952
rect 21272 14875 21324 14884
rect 21272 14841 21281 14875
rect 21281 14841 21315 14875
rect 21315 14841 21324 14875
rect 21272 14832 21324 14841
rect 22744 14832 22796 14884
rect 22928 14875 22980 14884
rect 22928 14841 22937 14875
rect 22937 14841 22971 14875
rect 22971 14841 22980 14875
rect 22928 14832 22980 14841
rect 23296 14943 23348 14952
rect 23296 14909 23305 14943
rect 23305 14909 23339 14943
rect 23339 14909 23348 14943
rect 23296 14900 23348 14909
rect 23756 14968 23808 15020
rect 23940 14968 23992 15020
rect 24308 14968 24360 15020
rect 24032 14900 24084 14952
rect 25136 14943 25188 14952
rect 25136 14909 25145 14943
rect 25145 14909 25179 14943
rect 25179 14909 25188 14943
rect 25136 14900 25188 14909
rect 25320 14943 25372 14952
rect 25320 14909 25329 14943
rect 25329 14909 25363 14943
rect 25363 14909 25372 14943
rect 25320 14900 25372 14909
rect 27528 15104 27580 15156
rect 28172 15104 28224 15156
rect 29368 15104 29420 15156
rect 30196 15104 30248 15156
rect 30840 15147 30892 15156
rect 30840 15113 30849 15147
rect 30849 15113 30883 15147
rect 30883 15113 30892 15147
rect 30840 15104 30892 15113
rect 25688 15036 25740 15088
rect 26608 14900 26660 14952
rect 27160 14968 27212 15020
rect 26884 14943 26936 14952
rect 26884 14909 26893 14943
rect 26893 14909 26927 14943
rect 26927 14909 26936 14943
rect 26884 14900 26936 14909
rect 26976 14943 27028 14952
rect 26976 14909 26985 14943
rect 26985 14909 27019 14943
rect 27019 14909 27028 14943
rect 27988 14968 28040 15020
rect 31116 14968 31168 15020
rect 26976 14900 27028 14909
rect 24216 14832 24268 14884
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 20352 14764 20404 14816
rect 20904 14764 20956 14816
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 28080 14875 28132 14884
rect 28080 14841 28089 14875
rect 28089 14841 28123 14875
rect 28123 14841 28132 14875
rect 28080 14832 28132 14841
rect 26792 14764 26844 14816
rect 26884 14764 26936 14816
rect 30472 14832 30524 14884
rect 28448 14764 28500 14816
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 15946 14662 15998 14714
rect 16010 14662 16062 14714
rect 16074 14662 16126 14714
rect 16138 14662 16190 14714
rect 16202 14662 16254 14714
rect 23720 14662 23772 14714
rect 23784 14662 23836 14714
rect 23848 14662 23900 14714
rect 23912 14662 23964 14714
rect 23976 14662 24028 14714
rect 31494 14662 31546 14714
rect 31558 14662 31610 14714
rect 31622 14662 31674 14714
rect 31686 14662 31738 14714
rect 31750 14662 31802 14714
rect 1216 14560 1268 14612
rect 2136 14560 2188 14612
rect 3976 14560 4028 14612
rect 4712 14560 4764 14612
rect 4804 14560 4856 14612
rect 5632 14560 5684 14612
rect 6092 14560 6144 14612
rect 7104 14560 7156 14612
rect 7932 14560 7984 14612
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 1768 14424 1820 14476
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 7564 14492 7616 14544
rect 2596 14424 2648 14476
rect 2780 14399 2832 14408
rect 2780 14365 2789 14399
rect 2789 14365 2823 14399
rect 2823 14365 2832 14399
rect 2780 14356 2832 14365
rect 5540 14424 5592 14476
rect 4160 14356 4212 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 6276 14424 6328 14476
rect 7104 14424 7156 14476
rect 7472 14424 7524 14476
rect 8392 14424 8444 14476
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 9220 14560 9272 14612
rect 9312 14560 9364 14612
rect 9496 14560 9548 14612
rect 10048 14560 10100 14612
rect 10324 14560 10376 14612
rect 9588 14492 9640 14544
rect 9036 14467 9088 14476
rect 9036 14433 9045 14467
rect 9045 14433 9079 14467
rect 9079 14433 9088 14467
rect 9036 14424 9088 14433
rect 3516 14220 3568 14272
rect 4528 14220 4580 14272
rect 7288 14356 7340 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 10048 14424 10100 14476
rect 11152 14467 11204 14476
rect 11152 14433 11161 14467
rect 11161 14433 11195 14467
rect 11195 14433 11204 14467
rect 11152 14424 11204 14433
rect 11244 14424 11296 14476
rect 13636 14560 13688 14612
rect 15476 14560 15528 14612
rect 11980 14492 12032 14544
rect 12532 14492 12584 14544
rect 14556 14492 14608 14544
rect 9772 14356 9824 14408
rect 9864 14356 9916 14408
rect 9404 14288 9456 14340
rect 7012 14220 7064 14272
rect 7472 14220 7524 14272
rect 8484 14220 8536 14272
rect 9128 14220 9180 14272
rect 9220 14220 9272 14272
rect 9680 14220 9732 14272
rect 10140 14288 10192 14340
rect 10324 14356 10376 14408
rect 11060 14356 11112 14408
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 12808 14424 12860 14476
rect 11980 14288 12032 14340
rect 10232 14220 10284 14272
rect 11612 14220 11664 14272
rect 13452 14356 13504 14408
rect 13912 14424 13964 14476
rect 14648 14467 14700 14476
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 14832 14492 14884 14544
rect 15384 14492 15436 14544
rect 16304 14560 16356 14612
rect 16580 14560 16632 14612
rect 17224 14560 17276 14612
rect 17408 14560 17460 14612
rect 18052 14560 18104 14612
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 19524 14560 19576 14612
rect 20996 14560 21048 14612
rect 21272 14560 21324 14612
rect 21916 14603 21968 14612
rect 21916 14569 21925 14603
rect 21925 14569 21959 14603
rect 21959 14569 21968 14603
rect 21916 14560 21968 14569
rect 22376 14560 22428 14612
rect 15016 14467 15068 14476
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 15476 14424 15528 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 17040 14492 17092 14544
rect 19984 14492 20036 14544
rect 23480 14492 23532 14544
rect 13452 14220 13504 14272
rect 14372 14356 14424 14408
rect 18052 14467 18104 14476
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 16580 14356 16632 14408
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 16488 14288 16540 14340
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 16396 14220 16448 14272
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 17316 14356 17368 14408
rect 18236 14356 18288 14408
rect 18420 14356 18472 14408
rect 17132 14220 17184 14272
rect 17960 14288 18012 14340
rect 18604 14424 18656 14476
rect 19248 14424 19300 14476
rect 19432 14424 19484 14476
rect 19800 14424 19852 14476
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 18972 14356 19024 14408
rect 19064 14399 19116 14408
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 19340 14356 19392 14408
rect 20444 14424 20496 14476
rect 22928 14424 22980 14476
rect 23388 14424 23440 14476
rect 23848 14424 23900 14476
rect 24676 14560 24728 14612
rect 20168 14356 20220 14408
rect 20352 14356 20404 14408
rect 21364 14356 21416 14408
rect 21548 14356 21600 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 20444 14288 20496 14340
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 22100 14356 22152 14365
rect 23020 14356 23072 14408
rect 24860 14492 24912 14544
rect 25780 14492 25832 14544
rect 24768 14467 24820 14476
rect 24768 14433 24777 14467
rect 24777 14433 24811 14467
rect 24811 14433 24820 14467
rect 24768 14424 24820 14433
rect 25228 14424 25280 14476
rect 25872 14467 25924 14476
rect 25872 14433 25881 14467
rect 25881 14433 25915 14467
rect 25915 14433 25924 14467
rect 25872 14424 25924 14433
rect 26240 14560 26292 14612
rect 26700 14560 26752 14612
rect 27160 14560 27212 14612
rect 27436 14492 27488 14544
rect 26608 14424 26660 14476
rect 26792 14467 26844 14476
rect 26792 14433 26801 14467
rect 26801 14433 26835 14467
rect 26835 14433 26844 14467
rect 26792 14424 26844 14433
rect 28264 14560 28316 14612
rect 29828 14560 29880 14612
rect 30104 14560 30156 14612
rect 30472 14560 30524 14612
rect 30932 14560 30984 14612
rect 31116 14560 31168 14612
rect 28540 14467 28592 14476
rect 22468 14288 22520 14340
rect 23940 14288 23992 14340
rect 24032 14288 24084 14340
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 28540 14424 28592 14433
rect 30380 14492 30432 14544
rect 28724 14424 28776 14476
rect 29092 14424 29144 14476
rect 29644 14424 29696 14476
rect 30012 14424 30064 14476
rect 30840 14424 30892 14476
rect 31024 14424 31076 14476
rect 25872 14288 25924 14340
rect 30104 14356 30156 14408
rect 19156 14220 19208 14272
rect 19248 14220 19300 14272
rect 20628 14220 20680 14272
rect 21180 14220 21232 14272
rect 22836 14220 22888 14272
rect 23204 14220 23256 14272
rect 24860 14220 24912 14272
rect 26884 14220 26936 14272
rect 27988 14220 28040 14272
rect 29828 14263 29880 14272
rect 29828 14229 29837 14263
rect 29837 14229 29871 14263
rect 29871 14229 29880 14263
rect 29828 14220 29880 14229
rect 30380 14220 30432 14272
rect 4285 14118 4337 14170
rect 4349 14118 4401 14170
rect 4413 14118 4465 14170
rect 4477 14118 4529 14170
rect 4541 14118 4593 14170
rect 12059 14118 12111 14170
rect 12123 14118 12175 14170
rect 12187 14118 12239 14170
rect 12251 14118 12303 14170
rect 12315 14118 12367 14170
rect 19833 14118 19885 14170
rect 19897 14118 19949 14170
rect 19961 14118 20013 14170
rect 20025 14118 20077 14170
rect 20089 14118 20141 14170
rect 27607 14118 27659 14170
rect 27671 14118 27723 14170
rect 27735 14118 27787 14170
rect 27799 14118 27851 14170
rect 27863 14118 27915 14170
rect 2780 14016 2832 14068
rect 3424 14016 3476 14068
rect 3516 14016 3568 14068
rect 4160 14016 4212 14068
rect 4896 14016 4948 14068
rect 5356 14016 5408 14068
rect 8300 13948 8352 14000
rect 9496 13948 9548 14000
rect 9864 13948 9916 14000
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 6368 13880 6420 13932
rect 7472 13880 7524 13932
rect 940 13812 992 13864
rect 1216 13855 1268 13864
rect 1216 13821 1225 13855
rect 1225 13821 1259 13855
rect 1259 13821 1268 13855
rect 1216 13812 1268 13821
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 5172 13812 5224 13864
rect 6920 13812 6972 13864
rect 2228 13744 2280 13796
rect 2780 13676 2832 13728
rect 3884 13676 3936 13728
rect 5816 13787 5868 13796
rect 5816 13753 5825 13787
rect 5825 13753 5859 13787
rect 5859 13753 5868 13787
rect 5816 13744 5868 13753
rect 4712 13676 4764 13728
rect 8944 13880 8996 13932
rect 9680 13880 9732 13932
rect 8576 13812 8628 13864
rect 9128 13812 9180 13864
rect 9404 13812 9456 13864
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 9588 13812 9640 13864
rect 9956 13812 10008 13864
rect 11152 14016 11204 14068
rect 11888 14016 11940 14068
rect 11980 14016 12032 14068
rect 13452 14016 13504 14068
rect 14188 14016 14240 14068
rect 14648 14016 14700 14068
rect 15660 14016 15712 14068
rect 16672 14016 16724 14068
rect 17592 14016 17644 14068
rect 17776 14016 17828 14068
rect 19340 14016 19392 14068
rect 20352 14016 20404 14068
rect 20444 14059 20496 14068
rect 20444 14025 20453 14059
rect 20453 14025 20487 14059
rect 20487 14025 20496 14059
rect 20444 14016 20496 14025
rect 20628 14059 20680 14068
rect 20628 14025 20637 14059
rect 20637 14025 20671 14059
rect 20671 14025 20680 14059
rect 20628 14016 20680 14025
rect 20720 14016 20772 14068
rect 21732 14016 21784 14068
rect 22744 14016 22796 14068
rect 23848 14016 23900 14068
rect 24400 14059 24452 14068
rect 24400 14025 24409 14059
rect 24409 14025 24443 14059
rect 24443 14025 24452 14059
rect 24400 14016 24452 14025
rect 11520 13880 11572 13932
rect 12992 13880 13044 13932
rect 17868 13948 17920 14000
rect 21548 13948 21600 14000
rect 24492 13948 24544 14000
rect 24584 13948 24636 14000
rect 24860 13948 24912 14000
rect 15384 13880 15436 13932
rect 10416 13812 10468 13864
rect 10784 13812 10836 13864
rect 13176 13812 13228 13864
rect 7380 13719 7432 13728
rect 7380 13685 7389 13719
rect 7389 13685 7423 13719
rect 7423 13685 7432 13719
rect 7380 13676 7432 13685
rect 7564 13676 7616 13728
rect 7932 13676 7984 13728
rect 9128 13676 9180 13728
rect 10324 13676 10376 13728
rect 10416 13676 10468 13728
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 10784 13676 10836 13728
rect 10968 13676 11020 13728
rect 11980 13744 12032 13796
rect 11244 13676 11296 13728
rect 14004 13812 14056 13864
rect 14188 13812 14240 13864
rect 15016 13812 15068 13864
rect 15660 13812 15712 13864
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17132 13880 17184 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 18972 13880 19024 13932
rect 22008 13880 22060 13932
rect 27436 14059 27488 14068
rect 27436 14025 27445 14059
rect 27445 14025 27479 14059
rect 27479 14025 27488 14059
rect 27436 14016 27488 14025
rect 30564 14016 30616 14068
rect 14464 13744 14516 13796
rect 15200 13744 15252 13796
rect 15476 13744 15528 13796
rect 17684 13812 17736 13864
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 19432 13812 19484 13864
rect 13820 13676 13872 13728
rect 14096 13676 14148 13728
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 15660 13719 15712 13728
rect 15660 13685 15669 13719
rect 15669 13685 15703 13719
rect 15703 13685 15712 13719
rect 15660 13676 15712 13685
rect 20168 13787 20220 13796
rect 20168 13753 20177 13787
rect 20177 13753 20211 13787
rect 20211 13753 20220 13787
rect 20168 13744 20220 13753
rect 21640 13812 21692 13864
rect 22652 13812 22704 13864
rect 22928 13812 22980 13864
rect 20996 13787 21048 13796
rect 20996 13753 21005 13787
rect 21005 13753 21039 13787
rect 21039 13753 21048 13787
rect 20996 13744 21048 13753
rect 21548 13744 21600 13796
rect 18512 13676 18564 13728
rect 20904 13676 20956 13728
rect 22744 13744 22796 13796
rect 23204 13744 23256 13796
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 24768 13812 24820 13864
rect 25412 13855 25464 13864
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 28264 13880 28316 13932
rect 28632 13880 28684 13932
rect 23572 13676 23624 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 24400 13744 24452 13796
rect 25228 13744 25280 13796
rect 24860 13676 24912 13728
rect 30196 13855 30248 13864
rect 30196 13821 30205 13855
rect 30205 13821 30239 13855
rect 30239 13821 30248 13855
rect 30196 13812 30248 13821
rect 30380 13812 30432 13864
rect 26516 13744 26568 13796
rect 26700 13744 26752 13796
rect 28356 13744 28408 13796
rect 27068 13676 27120 13728
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 15946 13574 15998 13626
rect 16010 13574 16062 13626
rect 16074 13574 16126 13626
rect 16138 13574 16190 13626
rect 16202 13574 16254 13626
rect 23720 13574 23772 13626
rect 23784 13574 23836 13626
rect 23848 13574 23900 13626
rect 23912 13574 23964 13626
rect 23976 13574 24028 13626
rect 31494 13574 31546 13626
rect 31558 13574 31610 13626
rect 31622 13574 31674 13626
rect 31686 13574 31738 13626
rect 31750 13574 31802 13626
rect 1216 13515 1268 13524
rect 1216 13481 1225 13515
rect 1225 13481 1259 13515
rect 1259 13481 1268 13515
rect 1216 13472 1268 13481
rect 2872 13472 2924 13524
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 2780 13404 2832 13456
rect 2136 13336 2188 13388
rect 2964 13336 3016 13388
rect 5540 13472 5592 13524
rect 5816 13472 5868 13524
rect 4712 13404 4764 13456
rect 2688 13268 2740 13320
rect 3700 13311 3752 13320
rect 3700 13277 3709 13311
rect 3709 13277 3743 13311
rect 3743 13277 3752 13311
rect 3700 13268 3752 13277
rect 940 13200 992 13252
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 8392 13472 8444 13524
rect 9772 13472 9824 13524
rect 10416 13472 10468 13524
rect 10692 13472 10744 13524
rect 12348 13472 12400 13524
rect 6920 13404 6972 13456
rect 8760 13404 8812 13456
rect 9128 13404 9180 13456
rect 9496 13447 9548 13456
rect 9496 13413 9505 13447
rect 9505 13413 9539 13447
rect 9539 13413 9548 13447
rect 9496 13404 9548 13413
rect 10508 13404 10560 13456
rect 5632 13268 5684 13277
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 6368 13336 6420 13388
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 9036 13379 9088 13388
rect 9036 13345 9045 13379
rect 9045 13345 9079 13379
rect 9079 13345 9088 13379
rect 9036 13336 9088 13345
rect 9588 13379 9640 13388
rect 9588 13345 9597 13379
rect 9597 13345 9631 13379
rect 9631 13345 9640 13379
rect 9588 13336 9640 13345
rect 8668 13200 8720 13252
rect 9036 13200 9088 13252
rect 7380 13132 7432 13184
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 8484 13132 8536 13184
rect 8576 13132 8628 13184
rect 9220 13200 9272 13252
rect 10048 13379 10100 13388
rect 10048 13345 10062 13379
rect 10062 13345 10096 13379
rect 10096 13345 10100 13379
rect 10048 13336 10100 13345
rect 10232 13336 10284 13388
rect 10140 13268 10192 13320
rect 12072 13404 12124 13456
rect 12256 13404 12308 13456
rect 13452 13404 13504 13456
rect 15568 13404 15620 13456
rect 16856 13404 16908 13456
rect 17040 13404 17092 13456
rect 10692 13336 10744 13388
rect 11244 13379 11296 13388
rect 11244 13345 11253 13379
rect 11253 13345 11287 13379
rect 11287 13345 11296 13379
rect 11244 13336 11296 13345
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 13544 13336 13596 13388
rect 11520 13268 11572 13320
rect 10232 13175 10284 13184
rect 10232 13141 10241 13175
rect 10241 13141 10275 13175
rect 10275 13141 10284 13175
rect 10232 13132 10284 13141
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 11428 13132 11480 13184
rect 11520 13132 11572 13184
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12072 13268 12124 13320
rect 14372 13336 14424 13388
rect 15016 13379 15068 13388
rect 15016 13345 15025 13379
rect 15025 13345 15059 13379
rect 15059 13345 15068 13379
rect 15016 13336 15068 13345
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 15844 13336 15896 13388
rect 12992 13200 13044 13252
rect 16212 13268 16264 13320
rect 16580 13336 16632 13388
rect 18052 13404 18104 13456
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 14004 13200 14056 13252
rect 14924 13200 14976 13252
rect 15752 13200 15804 13252
rect 11980 13132 12032 13184
rect 16672 13200 16724 13252
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 18972 13472 19024 13524
rect 20536 13472 20588 13524
rect 21180 13472 21232 13524
rect 21640 13472 21692 13524
rect 21824 13515 21876 13524
rect 21824 13481 21833 13515
rect 21833 13481 21867 13515
rect 21867 13481 21876 13515
rect 21824 13472 21876 13481
rect 22192 13515 22244 13524
rect 22192 13481 22201 13515
rect 22201 13481 22235 13515
rect 22235 13481 22244 13515
rect 22192 13472 22244 13481
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 17960 13200 18012 13252
rect 17868 13132 17920 13184
rect 18328 13200 18380 13252
rect 18512 13243 18564 13252
rect 18512 13209 18521 13243
rect 18521 13209 18555 13243
rect 18555 13209 18564 13243
rect 18512 13200 18564 13209
rect 19616 13336 19668 13388
rect 20812 13404 20864 13456
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 20260 13336 20312 13345
rect 20444 13336 20496 13388
rect 20168 13200 20220 13252
rect 19064 13132 19116 13184
rect 19432 13132 19484 13184
rect 20720 13336 20772 13388
rect 21180 13336 21232 13388
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 22652 13404 22704 13456
rect 24952 13472 25004 13524
rect 25044 13472 25096 13524
rect 25780 13472 25832 13524
rect 25872 13515 25924 13524
rect 25872 13481 25881 13515
rect 25881 13481 25915 13515
rect 25915 13481 25924 13515
rect 25872 13472 25924 13481
rect 22100 13379 22152 13388
rect 22100 13345 22109 13379
rect 22109 13345 22143 13379
rect 22143 13345 22152 13379
rect 22100 13336 22152 13345
rect 22744 13379 22796 13388
rect 22744 13345 22753 13379
rect 22753 13345 22787 13379
rect 22787 13345 22796 13379
rect 22744 13336 22796 13345
rect 24308 13404 24360 13456
rect 23572 13336 23624 13388
rect 23664 13379 23716 13388
rect 23664 13345 23673 13379
rect 23673 13345 23707 13379
rect 23707 13345 23716 13379
rect 23664 13336 23716 13345
rect 24032 13355 24041 13388
rect 24041 13355 24075 13388
rect 24075 13355 24084 13388
rect 24032 13336 24084 13355
rect 24216 13379 24268 13388
rect 24216 13345 24225 13379
rect 24225 13345 24259 13379
rect 24259 13345 24268 13379
rect 24216 13336 24268 13345
rect 24676 13336 24728 13388
rect 23204 13268 23256 13320
rect 24400 13268 24452 13320
rect 25596 13336 25648 13388
rect 23296 13243 23348 13252
rect 23296 13209 23305 13243
rect 23305 13209 23339 13243
rect 23339 13209 23348 13243
rect 23296 13200 23348 13209
rect 26424 13379 26476 13388
rect 26424 13345 26433 13379
rect 26433 13345 26467 13379
rect 26467 13345 26476 13379
rect 26424 13336 26476 13345
rect 26332 13268 26384 13320
rect 26700 13379 26752 13388
rect 26700 13345 26709 13379
rect 26709 13345 26743 13379
rect 26743 13345 26752 13379
rect 26700 13336 26752 13345
rect 27436 13336 27488 13388
rect 27712 13404 27764 13456
rect 28080 13404 28132 13456
rect 28356 13404 28408 13456
rect 30472 13472 30524 13524
rect 30840 13472 30892 13524
rect 31024 13472 31076 13524
rect 26976 13268 27028 13320
rect 27068 13268 27120 13320
rect 27712 13311 27764 13320
rect 27712 13277 27721 13311
rect 27721 13277 27755 13311
rect 27755 13277 27764 13311
rect 27712 13268 27764 13277
rect 27252 13200 27304 13252
rect 20352 13132 20404 13184
rect 20996 13132 21048 13184
rect 21456 13132 21508 13184
rect 21548 13132 21600 13184
rect 21916 13132 21968 13184
rect 24308 13132 24360 13184
rect 25780 13132 25832 13184
rect 29092 13336 29144 13388
rect 29828 13336 29880 13388
rect 28632 13243 28684 13252
rect 28632 13209 28641 13243
rect 28641 13209 28675 13243
rect 28675 13209 28684 13243
rect 28632 13200 28684 13209
rect 29460 13132 29512 13184
rect 4285 13030 4337 13082
rect 4349 13030 4401 13082
rect 4413 13030 4465 13082
rect 4477 13030 4529 13082
rect 4541 13030 4593 13082
rect 12059 13030 12111 13082
rect 12123 13030 12175 13082
rect 12187 13030 12239 13082
rect 12251 13030 12303 13082
rect 12315 13030 12367 13082
rect 19833 13030 19885 13082
rect 19897 13030 19949 13082
rect 19961 13030 20013 13082
rect 20025 13030 20077 13082
rect 20089 13030 20141 13082
rect 27607 13030 27659 13082
rect 27671 13030 27723 13082
rect 27735 13030 27787 13082
rect 27799 13030 27851 13082
rect 27863 13030 27915 13082
rect 4160 12928 4212 12980
rect 6276 12928 6328 12980
rect 7656 12928 7708 12980
rect 7932 12928 7984 12980
rect 9220 12928 9272 12980
rect 9496 12928 9548 12980
rect 10968 12928 11020 12980
rect 11428 12928 11480 12980
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 5448 12860 5500 12912
rect 940 12792 992 12844
rect 3148 12792 3200 12844
rect 2320 12724 2372 12776
rect 3424 12724 3476 12776
rect 3608 12724 3660 12776
rect 1308 12699 1360 12708
rect 1308 12665 1317 12699
rect 1317 12665 1351 12699
rect 1351 12665 1360 12699
rect 1308 12656 1360 12665
rect 4252 12724 4304 12776
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 6920 12792 6972 12844
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 7748 12792 7800 12844
rect 8116 12792 8168 12844
rect 3884 12656 3936 12708
rect 3976 12699 4028 12708
rect 3976 12665 3985 12699
rect 3985 12665 4019 12699
rect 4019 12665 4028 12699
rect 3976 12656 4028 12665
rect 4528 12656 4580 12708
rect 5632 12724 5684 12776
rect 9128 12792 9180 12844
rect 8852 12767 8904 12776
rect 4896 12656 4948 12708
rect 4160 12588 4212 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5448 12656 5500 12708
rect 7104 12656 7156 12708
rect 6552 12588 6604 12640
rect 8300 12656 8352 12708
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 9588 12860 9640 12912
rect 9496 12767 9548 12776
rect 9496 12733 9503 12767
rect 9503 12733 9548 12767
rect 9496 12724 9548 12733
rect 10416 12860 10468 12912
rect 10784 12860 10836 12912
rect 11152 12792 11204 12844
rect 11980 12792 12032 12844
rect 15108 12928 15160 12980
rect 15200 12928 15252 12980
rect 16396 12928 16448 12980
rect 16764 12928 16816 12980
rect 13084 12903 13136 12912
rect 13084 12869 13093 12903
rect 13093 12869 13127 12903
rect 13127 12869 13136 12903
rect 13084 12860 13136 12869
rect 15752 12860 15804 12912
rect 17776 12928 17828 12980
rect 18328 12928 18380 12980
rect 18420 12971 18472 12980
rect 18420 12937 18429 12971
rect 18429 12937 18463 12971
rect 18463 12937 18472 12971
rect 18420 12928 18472 12937
rect 19248 12928 19300 12980
rect 20168 12928 20220 12980
rect 19156 12860 19208 12912
rect 19524 12860 19576 12912
rect 20076 12903 20128 12912
rect 20076 12869 20085 12903
rect 20085 12869 20119 12903
rect 20119 12869 20128 12903
rect 20076 12860 20128 12869
rect 10600 12724 10652 12776
rect 10048 12656 10100 12708
rect 10324 12656 10376 12708
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 7932 12588 7984 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 9036 12588 9088 12640
rect 9312 12588 9364 12640
rect 9956 12588 10008 12640
rect 11060 12588 11112 12640
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 11704 12656 11756 12708
rect 12348 12656 12400 12708
rect 13820 12656 13872 12708
rect 15200 12724 15252 12776
rect 18052 12724 18104 12776
rect 20536 12971 20588 12980
rect 20536 12937 20545 12971
rect 20545 12937 20579 12971
rect 20579 12937 20588 12971
rect 20536 12928 20588 12937
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 20812 12928 20864 12980
rect 21272 12928 21324 12980
rect 22100 12928 22152 12980
rect 22744 12928 22796 12980
rect 23664 12928 23716 12980
rect 24584 12928 24636 12980
rect 24860 12928 24912 12980
rect 25044 12928 25096 12980
rect 25596 12928 25648 12980
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 25872 12928 25924 12980
rect 20904 12860 20956 12912
rect 14464 12656 14516 12708
rect 14924 12656 14976 12708
rect 15476 12699 15528 12708
rect 15476 12665 15485 12699
rect 15485 12665 15519 12699
rect 15519 12665 15528 12699
rect 15476 12656 15528 12665
rect 14280 12588 14332 12640
rect 15200 12588 15252 12640
rect 15844 12588 15896 12640
rect 17316 12656 17368 12708
rect 17868 12656 17920 12708
rect 18420 12656 18472 12708
rect 16764 12588 16816 12640
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 17960 12588 18012 12640
rect 19432 12699 19484 12708
rect 19432 12665 19441 12699
rect 19441 12665 19475 12699
rect 19475 12665 19484 12699
rect 19432 12656 19484 12665
rect 20628 12724 20680 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 19064 12588 19116 12640
rect 20904 12656 20956 12708
rect 21272 12724 21324 12776
rect 22008 12792 22060 12844
rect 22928 12835 22980 12844
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 22468 12724 22520 12776
rect 24124 12792 24176 12844
rect 25136 12792 25188 12844
rect 23204 12656 23256 12708
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 21548 12588 21600 12640
rect 21640 12588 21692 12640
rect 23572 12588 23624 12640
rect 24400 12588 24452 12640
rect 24860 12724 24912 12776
rect 24768 12699 24820 12708
rect 24768 12665 24777 12699
rect 24777 12665 24811 12699
rect 24811 12665 24820 12699
rect 24768 12656 24820 12665
rect 24676 12588 24728 12640
rect 25412 12724 25464 12776
rect 27068 12724 27120 12776
rect 27344 12928 27396 12980
rect 27988 12928 28040 12980
rect 29828 12928 29880 12980
rect 30288 12971 30340 12980
rect 30288 12937 30297 12971
rect 30297 12937 30331 12971
rect 30331 12937 30340 12971
rect 30288 12928 30340 12937
rect 30656 12928 30708 12980
rect 28172 12860 28224 12912
rect 27528 12835 27580 12844
rect 27528 12801 27537 12835
rect 27537 12801 27571 12835
rect 27571 12801 27580 12835
rect 27528 12792 27580 12801
rect 25044 12656 25096 12708
rect 26332 12699 26384 12708
rect 26332 12665 26341 12699
rect 26341 12665 26375 12699
rect 26375 12665 26384 12699
rect 26332 12656 26384 12665
rect 26884 12699 26936 12708
rect 26884 12665 26893 12699
rect 26893 12665 26927 12699
rect 26927 12665 26936 12699
rect 26884 12656 26936 12665
rect 27436 12724 27488 12776
rect 28264 12724 28316 12776
rect 30380 12724 30432 12776
rect 26976 12588 27028 12640
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 15946 12486 15998 12538
rect 16010 12486 16062 12538
rect 16074 12486 16126 12538
rect 16138 12486 16190 12538
rect 16202 12486 16254 12538
rect 23720 12486 23772 12538
rect 23784 12486 23836 12538
rect 23848 12486 23900 12538
rect 23912 12486 23964 12538
rect 23976 12486 24028 12538
rect 31494 12486 31546 12538
rect 31558 12486 31610 12538
rect 31622 12486 31674 12538
rect 31686 12486 31738 12538
rect 31750 12486 31802 12538
rect 1308 12384 1360 12436
rect 2780 12384 2832 12436
rect 3884 12384 3936 12436
rect 5356 12384 5408 12436
rect 6276 12384 6328 12436
rect 8760 12384 8812 12436
rect 9404 12384 9456 12436
rect 9680 12384 9732 12436
rect 3976 12359 4028 12368
rect 3976 12325 3985 12359
rect 3985 12325 4019 12359
rect 4019 12325 4028 12359
rect 3976 12316 4028 12325
rect 4068 12359 4120 12368
rect 4068 12325 4077 12359
rect 4077 12325 4111 12359
rect 4111 12325 4120 12359
rect 4068 12316 4120 12325
rect 4528 12316 4580 12368
rect 4620 12316 4672 12368
rect 6368 12316 6420 12368
rect 8484 12316 8536 12368
rect 9128 12316 9180 12368
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 4252 12248 4304 12300
rect 5080 12248 5132 12300
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 4804 12180 4856 12232
rect 7380 12248 7432 12300
rect 2136 12044 2188 12096
rect 3332 12044 3384 12096
rect 4620 12044 4672 12096
rect 5356 12044 5408 12096
rect 6000 12044 6052 12096
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 9312 12248 9364 12300
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9588 12316 9640 12368
rect 9956 12316 10008 12368
rect 9772 12248 9824 12300
rect 10232 12384 10284 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 14648 12384 14700 12436
rect 15476 12384 15528 12436
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 13452 12316 13504 12368
rect 15016 12316 15068 12368
rect 15752 12359 15804 12368
rect 16212 12384 16264 12436
rect 15752 12325 15793 12359
rect 15793 12325 15804 12359
rect 15752 12316 15804 12325
rect 10508 12180 10560 12232
rect 10048 12112 10100 12164
rect 10140 12112 10192 12164
rect 11060 12180 11112 12232
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 11796 12180 11848 12232
rect 11888 12180 11940 12232
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 10692 12112 10744 12164
rect 11152 12112 11204 12164
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 13820 12291 13872 12300
rect 13820 12257 13826 12291
rect 13826 12257 13872 12291
rect 13820 12248 13872 12257
rect 14096 12248 14148 12300
rect 15292 12248 15344 12300
rect 15936 12248 15988 12300
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 16948 12384 17000 12436
rect 18144 12384 18196 12436
rect 18236 12384 18288 12436
rect 18512 12384 18564 12436
rect 16212 12248 16264 12300
rect 16396 12248 16448 12300
rect 17040 12316 17092 12368
rect 16856 12248 16908 12300
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 19156 12384 19208 12436
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 12532 12044 12584 12096
rect 13084 12044 13136 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 14188 12044 14240 12096
rect 14740 12155 14792 12164
rect 14740 12121 14749 12155
rect 14749 12121 14783 12155
rect 14783 12121 14792 12155
rect 14740 12112 14792 12121
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 17868 12248 17920 12300
rect 17960 12248 18012 12300
rect 17684 12180 17736 12232
rect 18236 12291 18288 12300
rect 18236 12257 18245 12291
rect 18245 12257 18279 12291
rect 18279 12257 18288 12291
rect 18236 12248 18288 12257
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18604 12180 18656 12232
rect 18788 12291 18840 12300
rect 18788 12257 18797 12291
rect 18797 12257 18831 12291
rect 18831 12257 18840 12291
rect 18788 12248 18840 12257
rect 18880 12291 18932 12300
rect 18880 12257 18889 12291
rect 18889 12257 18923 12291
rect 18923 12257 18932 12291
rect 18880 12248 18932 12257
rect 18972 12180 19024 12232
rect 19156 12180 19208 12232
rect 20168 12384 20220 12436
rect 20996 12384 21048 12436
rect 21916 12384 21968 12436
rect 22284 12384 22336 12436
rect 20168 12291 20220 12300
rect 20168 12257 20177 12291
rect 20177 12257 20211 12291
rect 20211 12257 20220 12291
rect 20168 12248 20220 12257
rect 20628 12316 20680 12368
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 16120 12112 16172 12164
rect 16396 12112 16448 12164
rect 16856 12112 16908 12164
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 18052 12112 18104 12164
rect 18696 12112 18748 12164
rect 20536 12180 20588 12232
rect 20904 12180 20956 12232
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 22192 12316 22244 12368
rect 21916 12248 21968 12300
rect 24124 12384 24176 12436
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 27252 12384 27304 12436
rect 22652 12248 22704 12300
rect 23756 12291 23808 12300
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 20168 12112 20220 12164
rect 20260 12155 20312 12164
rect 20260 12121 20269 12155
rect 20269 12121 20303 12155
rect 20303 12121 20312 12155
rect 20260 12112 20312 12121
rect 20628 12112 20680 12164
rect 21088 12112 21140 12164
rect 22560 12112 22612 12164
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 23756 12257 23765 12291
rect 23765 12257 23799 12291
rect 23799 12257 23808 12291
rect 23756 12248 23808 12257
rect 24032 12248 24084 12300
rect 24492 12291 24544 12300
rect 24492 12257 24501 12291
rect 24501 12257 24535 12291
rect 24535 12257 24544 12291
rect 24492 12248 24544 12257
rect 25228 12316 25280 12368
rect 25688 12316 25740 12368
rect 24124 12223 24176 12232
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24216 12223 24268 12232
rect 24216 12189 24225 12223
rect 24225 12189 24259 12223
rect 24259 12189 24268 12223
rect 24216 12180 24268 12189
rect 26424 12180 26476 12232
rect 26884 12180 26936 12232
rect 19800 12044 19852 12096
rect 21732 12044 21784 12096
rect 22100 12044 22152 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 23756 12112 23808 12164
rect 23572 12087 23624 12096
rect 23572 12053 23581 12087
rect 23581 12053 23615 12087
rect 23615 12053 23624 12087
rect 23572 12044 23624 12053
rect 25044 12112 25096 12164
rect 26976 12087 27028 12096
rect 26976 12053 26985 12087
rect 26985 12053 27019 12087
rect 27019 12053 27028 12087
rect 26976 12044 27028 12053
rect 4285 11942 4337 11994
rect 4349 11942 4401 11994
rect 4413 11942 4465 11994
rect 4477 11942 4529 11994
rect 4541 11942 4593 11994
rect 12059 11942 12111 11994
rect 12123 11942 12175 11994
rect 12187 11942 12239 11994
rect 12251 11942 12303 11994
rect 12315 11942 12367 11994
rect 19833 11942 19885 11994
rect 19897 11942 19949 11994
rect 19961 11942 20013 11994
rect 20025 11942 20077 11994
rect 20089 11942 20141 11994
rect 27607 11942 27659 11994
rect 27671 11942 27723 11994
rect 27735 11942 27787 11994
rect 27799 11942 27851 11994
rect 27863 11942 27915 11994
rect 2964 11840 3016 11892
rect 3424 11840 3476 11892
rect 3608 11840 3660 11892
rect 4528 11840 4580 11892
rect 4804 11840 4856 11892
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 848 11679 900 11688
rect 848 11645 857 11679
rect 857 11645 891 11679
rect 891 11645 900 11679
rect 848 11636 900 11645
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 4436 11772 4488 11824
rect 7380 11772 7432 11824
rect 10784 11840 10836 11892
rect 10968 11883 11020 11892
rect 10968 11849 10977 11883
rect 10977 11849 11011 11883
rect 11011 11849 11020 11883
rect 10968 11840 11020 11849
rect 11612 11840 11664 11892
rect 11888 11840 11940 11892
rect 12992 11840 13044 11892
rect 10140 11772 10192 11824
rect 3516 11704 3568 11756
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6368 11704 6420 11756
rect 9036 11704 9088 11756
rect 1124 11611 1176 11620
rect 1124 11577 1133 11611
rect 1133 11577 1167 11611
rect 1167 11577 1176 11611
rect 1124 11568 1176 11577
rect 1768 11568 1820 11620
rect 2964 11568 3016 11620
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 8852 11636 8904 11688
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 6552 11568 6604 11620
rect 4896 11500 4948 11552
rect 5816 11500 5868 11552
rect 6828 11500 6880 11552
rect 8760 11611 8812 11620
rect 8760 11577 8769 11611
rect 8769 11577 8803 11611
rect 8803 11577 8812 11611
rect 9312 11636 9364 11688
rect 9588 11679 9640 11688
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10600 11772 10652 11824
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 10692 11636 10744 11688
rect 11244 11704 11296 11756
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 10968 11636 11020 11688
rect 11336 11636 11388 11688
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 11888 11679 11940 11688
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 12716 11704 12768 11756
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 8760 11568 8812 11577
rect 9036 11500 9088 11552
rect 9220 11500 9272 11552
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13084 11772 13136 11824
rect 14924 11840 14976 11892
rect 15568 11840 15620 11892
rect 13544 11772 13596 11824
rect 14188 11704 14240 11756
rect 16212 11772 16264 11824
rect 17776 11840 17828 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18144 11840 18196 11892
rect 20260 11840 20312 11892
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 15292 11636 15344 11688
rect 9956 11500 10008 11552
rect 11520 11500 11572 11552
rect 13820 11568 13872 11620
rect 15568 11568 15620 11620
rect 16120 11636 16172 11688
rect 16672 11704 16724 11756
rect 16856 11704 16908 11756
rect 20168 11772 20220 11824
rect 20444 11772 20496 11824
rect 20720 11772 20772 11824
rect 20812 11772 20864 11824
rect 21364 11840 21416 11892
rect 21456 11883 21508 11892
rect 21456 11849 21465 11883
rect 21465 11849 21499 11883
rect 21499 11849 21508 11883
rect 21456 11840 21508 11849
rect 22560 11840 22612 11892
rect 23480 11840 23532 11892
rect 23572 11840 23624 11892
rect 24032 11840 24084 11892
rect 26884 11840 26936 11892
rect 26976 11840 27028 11892
rect 22284 11772 22336 11824
rect 16764 11636 16816 11688
rect 18052 11704 18104 11756
rect 16856 11568 16908 11620
rect 18328 11636 18380 11688
rect 18788 11704 18840 11756
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 18880 11636 18932 11688
rect 19524 11704 19576 11756
rect 15384 11500 15436 11552
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 15936 11500 15988 11552
rect 16488 11500 16540 11552
rect 16948 11500 17000 11552
rect 18696 11568 18748 11620
rect 18420 11500 18472 11552
rect 19340 11568 19392 11620
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 20444 11636 20496 11688
rect 22192 11704 22244 11756
rect 20996 11679 21048 11688
rect 20996 11645 21027 11679
rect 21027 11645 21048 11679
rect 20996 11636 21048 11645
rect 21088 11636 21140 11688
rect 21456 11636 21508 11688
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 24860 11636 24912 11688
rect 26792 11636 26844 11688
rect 23296 11568 23348 11620
rect 24308 11568 24360 11620
rect 26332 11568 26384 11620
rect 20904 11500 20956 11552
rect 23388 11500 23440 11552
rect 24768 11500 24820 11552
rect 27528 11500 27580 11552
rect 28632 11543 28684 11552
rect 28632 11509 28641 11543
rect 28641 11509 28675 11543
rect 28675 11509 28684 11543
rect 28632 11500 28684 11509
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 15946 11398 15998 11450
rect 16010 11398 16062 11450
rect 16074 11398 16126 11450
rect 16138 11398 16190 11450
rect 16202 11398 16254 11450
rect 23720 11398 23772 11450
rect 23784 11398 23836 11450
rect 23848 11398 23900 11450
rect 23912 11398 23964 11450
rect 23976 11398 24028 11450
rect 31494 11398 31546 11450
rect 31558 11398 31610 11450
rect 31622 11398 31674 11450
rect 31686 11398 31738 11450
rect 31750 11398 31802 11450
rect 1124 11296 1176 11348
rect 2872 11296 2924 11348
rect 4436 11296 4488 11348
rect 4620 11296 4672 11348
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 2596 11160 2648 11212
rect 5172 11271 5224 11280
rect 5172 11237 5181 11271
rect 5181 11237 5215 11271
rect 5215 11237 5224 11271
rect 5172 11228 5224 11237
rect 5356 11228 5408 11280
rect 6552 11228 6604 11280
rect 4896 11203 4948 11212
rect 4896 11169 4906 11203
rect 4906 11169 4940 11203
rect 4940 11169 4948 11203
rect 4896 11160 4948 11169
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3424 11092 3476 11144
rect 3884 11135 3936 11144
rect 3884 11101 3893 11135
rect 3893 11101 3927 11135
rect 3927 11101 3936 11135
rect 3884 11092 3936 11101
rect 4896 11024 4948 11076
rect 3976 10956 4028 11008
rect 5632 11160 5684 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6184 11092 6236 11144
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 7840 11203 7892 11212
rect 7840 11169 7847 11203
rect 7847 11169 7892 11203
rect 7840 11160 7892 11169
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 8944 11160 8996 11212
rect 9128 11160 9180 11212
rect 9588 11160 9640 11212
rect 9956 11228 10008 11280
rect 5816 11024 5868 11076
rect 7196 11024 7248 11076
rect 7380 11024 7432 11076
rect 5540 10956 5592 11008
rect 6828 10956 6880 11008
rect 9864 11092 9916 11144
rect 8576 11024 8628 11076
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 9220 11024 9272 11076
rect 9680 11024 9732 11076
rect 10140 11203 10192 11212
rect 10140 11169 10150 11203
rect 10150 11169 10184 11203
rect 10184 11169 10192 11203
rect 10140 11160 10192 11169
rect 10692 11160 10744 11212
rect 12992 11296 13044 11348
rect 13268 11296 13320 11348
rect 11060 11228 11112 11280
rect 11244 11271 11296 11280
rect 11244 11237 11253 11271
rect 11253 11237 11287 11271
rect 11287 11237 11296 11271
rect 11244 11228 11296 11237
rect 11336 11271 11388 11280
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 11888 11228 11940 11280
rect 12164 11228 12216 11280
rect 12532 11228 12584 11280
rect 12716 11228 12768 11280
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 15476 11296 15528 11348
rect 15568 11296 15620 11348
rect 14096 11271 14148 11280
rect 11428 11160 11480 11212
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 10968 11092 11020 11144
rect 11336 11092 11388 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 12256 11092 12308 11144
rect 14096 11237 14123 11271
rect 14123 11237 14148 11271
rect 14096 11228 14148 11237
rect 14280 11271 14332 11280
rect 14280 11237 14289 11271
rect 14289 11237 14323 11271
rect 14323 11237 14332 11271
rect 14280 11228 14332 11237
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 10600 11024 10652 11076
rect 11612 11024 11664 11076
rect 14832 11160 14884 11212
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 15568 11160 15620 11169
rect 17776 11296 17828 11348
rect 16580 11228 16632 11280
rect 16396 11160 16448 11212
rect 14924 11092 14976 11144
rect 7840 10956 7892 11008
rect 9128 10956 9180 11008
rect 10784 10956 10836 11008
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 13268 11024 13320 11076
rect 14648 11024 14700 11076
rect 15016 11024 15068 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 13544 10956 13596 11008
rect 15844 10956 15896 11008
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 17684 11228 17736 11280
rect 18512 11296 18564 11348
rect 20536 11296 20588 11348
rect 20812 11296 20864 11348
rect 21456 11296 21508 11348
rect 29736 11339 29788 11348
rect 29736 11305 29745 11339
rect 29745 11305 29779 11339
rect 29779 11305 29788 11339
rect 29736 11296 29788 11305
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 17776 11203 17828 11212
rect 17776 11169 17785 11203
rect 17785 11169 17819 11203
rect 17819 11169 17828 11203
rect 17776 11160 17828 11169
rect 19800 11228 19852 11280
rect 20904 11228 20956 11280
rect 21364 11228 21416 11280
rect 18236 11160 18288 11212
rect 17224 11092 17276 11144
rect 17132 11024 17184 11076
rect 18052 11092 18104 11144
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 18972 11203 19024 11212
rect 18972 11169 18981 11203
rect 18981 11169 19015 11203
rect 19015 11169 19024 11203
rect 18972 11160 19024 11169
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 20352 11160 20404 11212
rect 20628 11203 20680 11212
rect 20628 11169 20637 11203
rect 20637 11169 20671 11203
rect 20671 11169 20680 11203
rect 20628 11160 20680 11169
rect 18328 11024 18380 11076
rect 19708 11092 19760 11144
rect 20536 11092 20588 11144
rect 21916 11160 21968 11212
rect 24676 11228 24728 11280
rect 26332 11228 26384 11280
rect 26608 11271 26660 11280
rect 26608 11237 26617 11271
rect 26617 11237 26651 11271
rect 26651 11237 26660 11271
rect 26608 11228 26660 11237
rect 22100 11092 22152 11144
rect 23020 11092 23072 11144
rect 24124 11092 24176 11144
rect 18052 10956 18104 11008
rect 19156 10956 19208 11008
rect 19340 10956 19392 11008
rect 20444 10956 20496 11008
rect 20720 10999 20772 11008
rect 20720 10965 20729 10999
rect 20729 10965 20763 10999
rect 20763 10965 20772 10999
rect 20720 10956 20772 10965
rect 21732 11024 21784 11076
rect 26608 11092 26660 11144
rect 26884 11160 26936 11212
rect 27068 11203 27120 11212
rect 27068 11169 27077 11203
rect 27077 11169 27111 11203
rect 27111 11169 27120 11203
rect 27068 11160 27120 11169
rect 28632 11160 28684 11212
rect 29920 11203 29972 11212
rect 29920 11169 29929 11203
rect 29929 11169 29963 11203
rect 29963 11169 29972 11203
rect 29920 11160 29972 11169
rect 26792 11024 26844 11076
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 22192 10956 22244 11008
rect 22928 10956 22980 11008
rect 24676 10956 24728 11008
rect 24952 10956 25004 11008
rect 29552 10999 29604 11008
rect 29552 10965 29561 10999
rect 29561 10965 29595 10999
rect 29595 10965 29604 10999
rect 29552 10956 29604 10965
rect 30196 10999 30248 11008
rect 30196 10965 30205 10999
rect 30205 10965 30239 10999
rect 30239 10965 30248 10999
rect 30196 10956 30248 10965
rect 4285 10854 4337 10906
rect 4349 10854 4401 10906
rect 4413 10854 4465 10906
rect 4477 10854 4529 10906
rect 4541 10854 4593 10906
rect 12059 10854 12111 10906
rect 12123 10854 12175 10906
rect 12187 10854 12239 10906
rect 12251 10854 12303 10906
rect 12315 10854 12367 10906
rect 19833 10854 19885 10906
rect 19897 10854 19949 10906
rect 19961 10854 20013 10906
rect 20025 10854 20077 10906
rect 20089 10854 20141 10906
rect 27607 10854 27659 10906
rect 27671 10854 27723 10906
rect 27735 10854 27787 10906
rect 27799 10854 27851 10906
rect 27863 10854 27915 10906
rect 2596 10752 2648 10804
rect 2136 10684 2188 10736
rect 3516 10684 3568 10736
rect 848 10659 900 10668
rect 848 10625 857 10659
rect 857 10625 891 10659
rect 891 10625 900 10659
rect 848 10616 900 10625
rect 2320 10616 2372 10668
rect 4068 10752 4120 10804
rect 4896 10752 4948 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 5908 10752 5960 10804
rect 7472 10752 7524 10804
rect 10048 10752 10100 10804
rect 10140 10752 10192 10804
rect 7748 10684 7800 10736
rect 9772 10684 9824 10736
rect 1768 10480 1820 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 4068 10548 4120 10600
rect 4160 10548 4212 10600
rect 3332 10480 3384 10532
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 6184 10616 6236 10668
rect 6276 10659 6328 10668
rect 6276 10625 6285 10659
rect 6285 10625 6319 10659
rect 6319 10625 6328 10659
rect 6276 10616 6328 10625
rect 6920 10616 6972 10668
rect 9312 10616 9364 10668
rect 4804 10412 4856 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5356 10412 5408 10464
rect 6828 10548 6880 10600
rect 7656 10548 7708 10600
rect 8024 10480 8076 10532
rect 7564 10412 7616 10464
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 8944 10548 8996 10600
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 9588 10523 9640 10532
rect 9588 10489 9597 10523
rect 9597 10489 9631 10523
rect 9631 10489 9640 10523
rect 9588 10480 9640 10489
rect 10508 10616 10560 10668
rect 11612 10616 11664 10668
rect 13176 10795 13228 10804
rect 13176 10761 13185 10795
rect 13185 10761 13219 10795
rect 13219 10761 13228 10795
rect 13176 10752 13228 10761
rect 13544 10752 13596 10804
rect 13728 10752 13780 10804
rect 15108 10752 15160 10804
rect 16948 10752 17000 10804
rect 18236 10752 18288 10804
rect 18696 10752 18748 10804
rect 19156 10752 19208 10804
rect 12440 10616 12492 10668
rect 14464 10684 14516 10736
rect 13268 10616 13320 10668
rect 14740 10616 14792 10668
rect 19340 10684 19392 10736
rect 14832 10548 14884 10600
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 17960 10616 18012 10668
rect 20352 10752 20404 10804
rect 21456 10752 21508 10804
rect 24400 10752 24452 10804
rect 24584 10795 24636 10804
rect 24584 10761 24593 10795
rect 24593 10761 24627 10795
rect 24627 10761 24636 10795
rect 24584 10752 24636 10761
rect 26516 10727 26568 10736
rect 26516 10693 26525 10727
rect 26525 10693 26559 10727
rect 26559 10693 26568 10727
rect 26516 10684 26568 10693
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 11336 10480 11388 10532
rect 8760 10412 8812 10464
rect 9128 10412 9180 10464
rect 9496 10412 9548 10464
rect 10968 10412 11020 10464
rect 11796 10412 11848 10464
rect 13544 10523 13596 10532
rect 13544 10489 13553 10523
rect 13553 10489 13587 10523
rect 13587 10489 13596 10523
rect 13544 10480 13596 10489
rect 15660 10480 15712 10532
rect 15752 10480 15804 10532
rect 19064 10548 19116 10600
rect 14924 10412 14976 10464
rect 16396 10412 16448 10464
rect 16580 10412 16632 10464
rect 17316 10412 17368 10464
rect 18972 10412 19024 10464
rect 23020 10616 23072 10668
rect 23388 10616 23440 10668
rect 26792 10616 26844 10668
rect 20168 10480 20220 10532
rect 19524 10412 19576 10464
rect 20628 10412 20680 10464
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 21640 10591 21692 10600
rect 21640 10557 21649 10591
rect 21649 10557 21683 10591
rect 21683 10557 21692 10591
rect 21640 10548 21692 10557
rect 28816 10548 28868 10600
rect 29092 10548 29144 10600
rect 22928 10480 22980 10532
rect 23112 10412 23164 10464
rect 23480 10480 23532 10532
rect 25780 10480 25832 10532
rect 26056 10523 26108 10532
rect 26056 10489 26065 10523
rect 26065 10489 26099 10523
rect 26099 10489 26108 10523
rect 26056 10480 26108 10489
rect 27528 10480 27580 10532
rect 25688 10412 25740 10464
rect 27712 10480 27764 10532
rect 29000 10523 29052 10532
rect 29000 10489 29009 10523
rect 29009 10489 29043 10523
rect 29043 10489 29052 10523
rect 29000 10480 29052 10489
rect 30196 10548 30248 10600
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 15946 10310 15998 10362
rect 16010 10310 16062 10362
rect 16074 10310 16126 10362
rect 16138 10310 16190 10362
rect 16202 10310 16254 10362
rect 23720 10310 23772 10362
rect 23784 10310 23836 10362
rect 23848 10310 23900 10362
rect 23912 10310 23964 10362
rect 23976 10310 24028 10362
rect 31494 10310 31546 10362
rect 31558 10310 31610 10362
rect 31622 10310 31674 10362
rect 31686 10310 31738 10362
rect 31750 10310 31802 10362
rect 2596 10208 2648 10260
rect 2780 10208 2832 10260
rect 3700 10208 3752 10260
rect 4988 10208 5040 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 7012 10208 7064 10260
rect 7564 10208 7616 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 9036 10208 9088 10260
rect 2320 10140 2372 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 10416 10208 10468 10260
rect 11796 10208 11848 10260
rect 11888 10208 11940 10260
rect 10508 10140 10560 10192
rect 2780 10004 2832 10056
rect 3424 10004 3476 10056
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 5356 10072 5408 10124
rect 7012 10072 7064 10124
rect 7472 10004 7524 10056
rect 8668 10072 8720 10124
rect 10140 10072 10192 10124
rect 7932 10004 7984 10056
rect 8760 10004 8812 10056
rect 4896 9936 4948 9988
rect 1768 9868 1820 9920
rect 3516 9868 3568 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7380 9868 7432 9920
rect 9956 9868 10008 9920
rect 10876 10004 10928 10056
rect 11060 10072 11112 10124
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 11520 10072 11572 10124
rect 12624 10140 12676 10192
rect 14648 10208 14700 10260
rect 14832 10208 14884 10260
rect 15200 10208 15252 10260
rect 13820 10140 13872 10192
rect 12348 10072 12400 10124
rect 14096 10072 14148 10124
rect 15752 10140 15804 10192
rect 16304 10140 16356 10192
rect 16396 10140 16448 10192
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 17868 10208 17920 10260
rect 18420 10208 18472 10260
rect 18512 10208 18564 10260
rect 18604 10208 18656 10260
rect 19156 10208 19208 10260
rect 19432 10208 19484 10260
rect 19708 10208 19760 10260
rect 15568 10072 15620 10124
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11612 10004 11664 10056
rect 12532 10004 12584 10056
rect 13728 10004 13780 10056
rect 14464 10004 14516 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 11888 9936 11940 9988
rect 12348 9936 12400 9988
rect 17224 10072 17276 10124
rect 17316 10072 17368 10124
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 18052 10115 18104 10124
rect 18052 10081 18061 10115
rect 18061 10081 18095 10115
rect 18095 10081 18104 10115
rect 18052 10072 18104 10081
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 18880 10072 18932 10124
rect 20536 10140 20588 10192
rect 20996 10140 21048 10192
rect 21640 10208 21692 10260
rect 22652 10208 22704 10260
rect 22928 10140 22980 10192
rect 24584 10208 24636 10260
rect 25688 10251 25740 10260
rect 25688 10217 25697 10251
rect 25697 10217 25731 10251
rect 25731 10217 25740 10251
rect 25688 10208 25740 10217
rect 26056 10208 26108 10260
rect 26516 10208 26568 10260
rect 11060 9868 11112 9920
rect 11152 9868 11204 9920
rect 12716 9868 12768 9920
rect 15568 9868 15620 9920
rect 17684 9979 17736 9988
rect 17684 9945 17693 9979
rect 17693 9945 17727 9979
rect 17727 9945 17736 9979
rect 17684 9936 17736 9945
rect 19340 10004 19392 10056
rect 18144 9868 18196 9920
rect 18972 9868 19024 9920
rect 19248 9868 19300 9920
rect 23388 10072 23440 10124
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 21640 10004 21692 10056
rect 22468 10004 22520 10056
rect 22652 10004 22704 10056
rect 23296 9936 23348 9988
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23848 10072 23900 10124
rect 23940 10072 23992 10124
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 24768 10072 24820 10124
rect 25412 10072 25464 10124
rect 27712 10208 27764 10260
rect 29000 10208 29052 10260
rect 28816 10140 28868 10192
rect 29552 10140 29604 10192
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25228 10004 25280 10056
rect 26056 10004 26108 10056
rect 26608 10004 26660 10056
rect 26700 10047 26752 10056
rect 26700 10013 26709 10047
rect 26709 10013 26743 10047
rect 26743 10013 26752 10047
rect 26700 10004 26752 10013
rect 27620 10047 27672 10056
rect 27620 10013 27629 10047
rect 27629 10013 27663 10047
rect 27663 10013 27672 10047
rect 27620 10004 27672 10013
rect 23756 9936 23808 9988
rect 25412 9936 25464 9988
rect 23940 9868 23992 9920
rect 24952 9868 25004 9920
rect 25872 9868 25924 9920
rect 4285 9766 4337 9818
rect 4349 9766 4401 9818
rect 4413 9766 4465 9818
rect 4477 9766 4529 9818
rect 4541 9766 4593 9818
rect 12059 9766 12111 9818
rect 12123 9766 12175 9818
rect 12187 9766 12239 9818
rect 12251 9766 12303 9818
rect 12315 9766 12367 9818
rect 19833 9766 19885 9818
rect 19897 9766 19949 9818
rect 19961 9766 20013 9818
rect 20025 9766 20077 9818
rect 20089 9766 20141 9818
rect 27607 9766 27659 9818
rect 27671 9766 27723 9818
rect 27735 9766 27787 9818
rect 27799 9766 27851 9818
rect 27863 9766 27915 9818
rect 3884 9664 3936 9716
rect 6276 9664 6328 9716
rect 7012 9664 7064 9716
rect 8024 9664 8076 9716
rect 8944 9664 8996 9716
rect 2504 9596 2556 9648
rect 2136 9460 2188 9512
rect 1768 9392 1820 9444
rect 4988 9596 5040 9648
rect 6460 9596 6512 9648
rect 6552 9639 6604 9648
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4528 9460 4580 9469
rect 4712 9503 4764 9512
rect 4712 9469 4719 9503
rect 4719 9469 4764 9503
rect 4712 9460 4764 9469
rect 4160 9392 4212 9444
rect 5172 9460 5224 9512
rect 7564 9596 7616 9648
rect 8852 9596 8904 9648
rect 11520 9664 11572 9716
rect 11612 9664 11664 9716
rect 11796 9664 11848 9716
rect 11980 9664 12032 9716
rect 6460 9460 6512 9512
rect 7012 9503 7064 9512
rect 7012 9469 7019 9503
rect 7019 9469 7064 9503
rect 7012 9460 7064 9469
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 7380 9460 7432 9512
rect 7932 9528 7984 9580
rect 5448 9392 5500 9444
rect 4712 9324 4764 9376
rect 5264 9324 5316 9376
rect 7564 9324 7616 9376
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9772 9571 9824 9580
rect 9036 9528 9088 9537
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 8300 9460 8352 9512
rect 8024 9324 8076 9376
rect 8668 9324 8720 9376
rect 8852 9435 8904 9444
rect 8852 9401 8861 9435
rect 8861 9401 8895 9435
rect 8895 9401 8904 9435
rect 8852 9392 8904 9401
rect 9404 9435 9456 9444
rect 9404 9401 9413 9435
rect 9413 9401 9447 9435
rect 9447 9401 9456 9435
rect 9404 9392 9456 9401
rect 9864 9392 9916 9444
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 11612 9528 11664 9580
rect 12532 9596 12584 9648
rect 12716 9664 12768 9716
rect 13636 9664 13688 9716
rect 13728 9664 13780 9716
rect 17408 9664 17460 9716
rect 17684 9664 17736 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 13084 9596 13136 9648
rect 12900 9528 12952 9580
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 10048 9460 10100 9469
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 12532 9460 12584 9512
rect 8944 9324 8996 9376
rect 10140 9324 10192 9376
rect 10508 9324 10560 9376
rect 11520 9392 11572 9444
rect 11704 9392 11756 9444
rect 11980 9324 12032 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 12808 9324 12860 9376
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 13176 9392 13228 9444
rect 14004 9528 14056 9580
rect 15384 9528 15436 9580
rect 16396 9596 16448 9648
rect 15844 9528 15896 9580
rect 16764 9639 16816 9648
rect 16764 9605 16773 9639
rect 16773 9605 16807 9639
rect 16807 9605 16816 9639
rect 16764 9596 16816 9605
rect 17592 9528 17644 9580
rect 15476 9460 15528 9512
rect 16580 9460 16632 9512
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 17684 9503 17736 9512
rect 17684 9469 17693 9503
rect 17693 9469 17727 9503
rect 17727 9469 17736 9503
rect 17684 9460 17736 9469
rect 21180 9707 21232 9716
rect 21180 9673 21189 9707
rect 21189 9673 21223 9707
rect 21223 9673 21232 9707
rect 21180 9664 21232 9673
rect 21732 9707 21784 9716
rect 21732 9673 21741 9707
rect 21741 9673 21775 9707
rect 21775 9673 21784 9707
rect 21732 9664 21784 9673
rect 23388 9664 23440 9716
rect 30196 9664 30248 9716
rect 20996 9596 21048 9648
rect 21824 9596 21876 9648
rect 23480 9596 23532 9648
rect 23572 9596 23624 9648
rect 18604 9460 18656 9512
rect 13820 9392 13872 9444
rect 16304 9435 16356 9444
rect 16304 9401 16313 9435
rect 16313 9401 16347 9435
rect 16347 9401 16356 9435
rect 16304 9392 16356 9401
rect 16396 9392 16448 9444
rect 19156 9503 19208 9512
rect 19156 9469 19165 9503
rect 19165 9469 19199 9503
rect 19199 9469 19208 9503
rect 19156 9460 19208 9469
rect 19248 9460 19300 9512
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 23388 9460 23440 9512
rect 24124 9460 24176 9512
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 24952 9596 25004 9648
rect 24308 9460 24360 9512
rect 25688 9503 25740 9512
rect 25688 9469 25697 9503
rect 25697 9469 25731 9503
rect 25731 9469 25740 9503
rect 25688 9460 25740 9469
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 16580 9324 16632 9376
rect 17316 9324 17368 9376
rect 17776 9324 17828 9376
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 17868 9324 17920 9333
rect 18512 9324 18564 9376
rect 19616 9392 19668 9444
rect 19984 9392 20036 9444
rect 20996 9392 21048 9444
rect 22008 9392 22060 9444
rect 19340 9324 19392 9376
rect 20536 9324 20588 9376
rect 20628 9324 20680 9376
rect 21732 9324 21784 9376
rect 22560 9324 22612 9376
rect 23296 9324 23348 9376
rect 25136 9392 25188 9444
rect 25320 9392 25372 9444
rect 25412 9435 25464 9444
rect 25412 9401 25421 9435
rect 25421 9401 25455 9435
rect 25455 9401 25464 9435
rect 25412 9392 25464 9401
rect 24400 9324 24452 9376
rect 25872 9392 25924 9444
rect 28172 9528 28224 9580
rect 28908 9528 28960 9580
rect 26700 9460 26752 9512
rect 26056 9324 26108 9376
rect 26332 9324 26384 9376
rect 26424 9367 26476 9376
rect 26424 9333 26433 9367
rect 26433 9333 26467 9367
rect 26467 9333 26476 9367
rect 26424 9324 26476 9333
rect 26792 9367 26844 9376
rect 26792 9333 26801 9367
rect 26801 9333 26835 9367
rect 26835 9333 26844 9367
rect 26792 9324 26844 9333
rect 27160 9392 27212 9444
rect 27528 9324 27580 9376
rect 27804 9367 27856 9376
rect 27804 9333 27813 9367
rect 27813 9333 27847 9367
rect 27847 9333 27856 9367
rect 27804 9324 27856 9333
rect 28356 9324 28408 9376
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 15946 9222 15998 9274
rect 16010 9222 16062 9274
rect 16074 9222 16126 9274
rect 16138 9222 16190 9274
rect 16202 9222 16254 9274
rect 23720 9222 23772 9274
rect 23784 9222 23836 9274
rect 23848 9222 23900 9274
rect 23912 9222 23964 9274
rect 23976 9222 24028 9274
rect 31494 9222 31546 9274
rect 31558 9222 31610 9274
rect 31622 9222 31674 9274
rect 31686 9222 31738 9274
rect 31750 9222 31802 9274
rect 2044 9120 2096 9172
rect 2596 9120 2648 9172
rect 4528 9120 4580 9172
rect 3884 9052 3936 9104
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 3516 8984 3568 9036
rect 5540 9120 5592 9172
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 4160 8916 4212 8968
rect 4804 8916 4856 8968
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5172 8984 5224 9036
rect 7656 9120 7708 9172
rect 8484 9120 8536 9172
rect 3608 8848 3660 8900
rect 5632 8916 5684 8968
rect 6368 9052 6420 9104
rect 6460 8984 6512 9036
rect 8576 9052 8628 9104
rect 9036 9052 9088 9104
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 10508 9163 10560 9172
rect 10508 9129 10517 9163
rect 10517 9129 10551 9163
rect 10551 9129 10560 9163
rect 10508 9120 10560 9129
rect 10784 9120 10836 9172
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 12716 9163 12768 9172
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 7012 9027 7064 9036
rect 7012 8993 7019 9027
rect 7019 8993 7064 9027
rect 7012 8984 7064 8993
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 7288 9027 7340 9036
rect 7288 8993 7302 9027
rect 7302 8993 7336 9027
rect 7336 8993 7340 9027
rect 7288 8984 7340 8993
rect 7472 8984 7524 9036
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 10232 9052 10284 9104
rect 14096 9052 14148 9104
rect 15568 9052 15620 9104
rect 10324 8984 10376 9036
rect 11152 8984 11204 9036
rect 11980 8984 12032 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 12256 8984 12308 9036
rect 12992 8984 13044 9036
rect 13084 8984 13136 9036
rect 3148 8780 3200 8832
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 4620 8780 4672 8832
rect 4804 8780 4856 8832
rect 4988 8780 5040 8832
rect 5172 8780 5224 8832
rect 6828 8848 6880 8900
rect 7104 8848 7156 8900
rect 8024 8848 8076 8900
rect 8116 8891 8168 8900
rect 8116 8857 8125 8891
rect 8125 8857 8159 8891
rect 8159 8857 8168 8891
rect 8116 8848 8168 8857
rect 8576 8848 8628 8900
rect 8760 8848 8812 8900
rect 8944 8848 8996 8900
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 11060 8916 11112 8968
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 13544 8916 13596 8968
rect 13912 8916 13964 8968
rect 15384 8916 15436 8968
rect 16396 9120 16448 9172
rect 17776 9120 17828 9172
rect 17040 9052 17092 9104
rect 16304 8984 16356 9036
rect 18420 8984 18472 9036
rect 12716 8848 12768 8900
rect 13084 8848 13136 8900
rect 18604 8916 18656 8968
rect 19248 8916 19300 8968
rect 18420 8848 18472 8900
rect 18696 8848 18748 8900
rect 19708 8916 19760 8968
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 20260 9120 20312 9172
rect 21364 9120 21416 9172
rect 21732 9163 21784 9172
rect 21732 9129 21741 9163
rect 21741 9129 21775 9163
rect 21775 9129 21784 9163
rect 21732 9120 21784 9129
rect 24124 9120 24176 9172
rect 25964 9120 26016 9172
rect 26424 9120 26476 9172
rect 28356 9120 28408 9172
rect 21180 9052 21232 9104
rect 22560 9052 22612 9104
rect 22376 8984 22428 9036
rect 22744 8984 22796 9036
rect 23112 9095 23164 9104
rect 23112 9061 23121 9095
rect 23121 9061 23155 9095
rect 23155 9061 23164 9095
rect 23112 9052 23164 9061
rect 24492 9052 24544 9104
rect 24860 9052 24912 9104
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 22192 8916 22244 8968
rect 23756 8916 23808 8968
rect 25872 8984 25924 9036
rect 27436 9052 27488 9104
rect 29092 9052 29144 9104
rect 26148 8916 26200 8968
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 8392 8780 8444 8832
rect 9496 8780 9548 8832
rect 9680 8780 9732 8832
rect 9956 8780 10008 8832
rect 10692 8780 10744 8832
rect 11336 8780 11388 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 16764 8780 16816 8832
rect 16856 8780 16908 8832
rect 20720 8780 20772 8832
rect 24768 8780 24820 8832
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 26608 8848 26660 8900
rect 26792 8780 26844 8832
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 4285 8678 4337 8730
rect 4349 8678 4401 8730
rect 4413 8678 4465 8730
rect 4477 8678 4529 8730
rect 4541 8678 4593 8730
rect 12059 8678 12111 8730
rect 12123 8678 12175 8730
rect 12187 8678 12239 8730
rect 12251 8678 12303 8730
rect 12315 8678 12367 8730
rect 19833 8678 19885 8730
rect 19897 8678 19949 8730
rect 19961 8678 20013 8730
rect 20025 8678 20077 8730
rect 20089 8678 20141 8730
rect 27607 8678 27659 8730
rect 27671 8678 27723 8730
rect 27735 8678 27787 8730
rect 27799 8678 27851 8730
rect 27863 8678 27915 8730
rect 2412 8576 2464 8628
rect 2504 8508 2556 8560
rect 848 8415 900 8424
rect 848 8381 857 8415
rect 857 8381 891 8415
rect 891 8381 900 8415
rect 848 8372 900 8381
rect 3976 8576 4028 8628
rect 4160 8576 4212 8628
rect 4252 8576 4304 8628
rect 4896 8576 4948 8628
rect 5172 8576 5224 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7104 8576 7156 8628
rect 7564 8576 7616 8628
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 8024 8576 8076 8628
rect 8392 8576 8444 8628
rect 9036 8576 9088 8628
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 10232 8576 10284 8628
rect 10324 8576 10376 8628
rect 8392 8440 8444 8492
rect 8668 8440 8720 8492
rect 1216 8304 1268 8356
rect 2964 8304 3016 8356
rect 3056 8304 3108 8356
rect 4252 8347 4304 8356
rect 4252 8313 4261 8347
rect 4261 8313 4295 8347
rect 4295 8313 4304 8347
rect 4252 8304 4304 8313
rect 6920 8372 6972 8424
rect 7656 8372 7708 8424
rect 3148 8236 3200 8288
rect 3424 8236 3476 8288
rect 4712 8304 4764 8356
rect 5540 8304 5592 8356
rect 7012 8304 7064 8356
rect 8392 8304 8444 8356
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 5172 8236 5224 8288
rect 5356 8236 5408 8288
rect 6736 8236 6788 8288
rect 7656 8236 7708 8288
rect 8484 8236 8536 8288
rect 10692 8508 10744 8560
rect 11336 8576 11388 8628
rect 11520 8576 11572 8628
rect 12348 8576 12400 8628
rect 13268 8576 13320 8628
rect 9588 8372 9640 8424
rect 9772 8372 9824 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 10508 8440 10560 8492
rect 11980 8440 12032 8492
rect 12072 8440 12124 8492
rect 13452 8508 13504 8560
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13084 8440 13136 8492
rect 9956 8372 10008 8381
rect 13360 8372 13412 8424
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 14832 8372 14884 8424
rect 15108 8576 15160 8628
rect 15752 8576 15804 8628
rect 16488 8619 16540 8628
rect 16488 8585 16497 8619
rect 16497 8585 16531 8619
rect 16531 8585 16540 8619
rect 16488 8576 16540 8585
rect 16580 8576 16632 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17684 8576 17736 8628
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 20352 8576 20404 8628
rect 21364 8576 21416 8628
rect 23112 8576 23164 8628
rect 23572 8576 23624 8628
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 24308 8619 24360 8628
rect 24308 8585 24317 8619
rect 24317 8585 24351 8619
rect 24351 8585 24360 8619
rect 24308 8576 24360 8585
rect 24860 8576 24912 8628
rect 26148 8619 26200 8628
rect 26148 8585 26157 8619
rect 26157 8585 26191 8619
rect 26191 8585 26200 8619
rect 26148 8576 26200 8585
rect 26240 8576 26292 8628
rect 15200 8508 15252 8560
rect 15292 8440 15344 8492
rect 16672 8508 16724 8560
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 9312 8236 9364 8288
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 10140 8236 10192 8288
rect 10324 8304 10376 8356
rect 10508 8304 10560 8356
rect 11336 8347 11388 8356
rect 11336 8313 11345 8347
rect 11345 8313 11379 8347
rect 11379 8313 11388 8347
rect 11336 8304 11388 8313
rect 12716 8304 12768 8356
rect 12900 8347 12952 8356
rect 12900 8313 12909 8347
rect 12909 8313 12943 8347
rect 12943 8313 12952 8347
rect 12900 8304 12952 8313
rect 10784 8236 10836 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 14188 8304 14240 8356
rect 13636 8236 13688 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 15200 8279 15252 8288
rect 15200 8245 15209 8279
rect 15209 8245 15243 8279
rect 15243 8245 15252 8279
rect 15200 8236 15252 8245
rect 15476 8347 15528 8356
rect 15476 8313 15485 8347
rect 15485 8313 15519 8347
rect 15519 8313 15528 8347
rect 15476 8304 15528 8313
rect 15568 8236 15620 8288
rect 16396 8236 16448 8288
rect 16764 8372 16816 8424
rect 16580 8304 16632 8356
rect 17960 8372 18012 8424
rect 18052 8372 18104 8424
rect 17960 8236 18012 8288
rect 18420 8304 18472 8356
rect 19248 8508 19300 8560
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20444 8440 20496 8492
rect 22560 8440 22612 8492
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23204 8483 23256 8492
rect 23204 8449 23213 8483
rect 23213 8449 23247 8483
rect 23247 8449 23256 8483
rect 23204 8440 23256 8449
rect 23296 8440 23348 8492
rect 23756 8440 23808 8492
rect 24676 8440 24728 8492
rect 27528 8576 27580 8628
rect 28632 8576 28684 8628
rect 27436 8551 27488 8560
rect 27436 8517 27445 8551
rect 27445 8517 27479 8551
rect 27479 8517 27488 8551
rect 27436 8508 27488 8517
rect 22008 8372 22060 8424
rect 22468 8372 22520 8424
rect 20260 8304 20312 8356
rect 23940 8304 23992 8356
rect 25780 8372 25832 8424
rect 24768 8304 24820 8356
rect 26700 8304 26752 8356
rect 28172 8372 28224 8424
rect 19524 8236 19576 8288
rect 21732 8236 21784 8288
rect 23388 8236 23440 8288
rect 23572 8236 23624 8288
rect 25320 8236 25372 8288
rect 27988 8236 28040 8288
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 15946 8134 15998 8186
rect 16010 8134 16062 8186
rect 16074 8134 16126 8186
rect 16138 8134 16190 8186
rect 16202 8134 16254 8186
rect 23720 8134 23772 8186
rect 23784 8134 23836 8186
rect 23848 8134 23900 8186
rect 23912 8134 23964 8186
rect 23976 8134 24028 8186
rect 31494 8134 31546 8186
rect 31558 8134 31610 8186
rect 31622 8134 31674 8186
rect 31686 8134 31738 8186
rect 31750 8134 31802 8186
rect 1584 8032 1636 8084
rect 3700 8032 3752 8084
rect 7012 8032 7064 8084
rect 7564 8032 7616 8084
rect 8852 8032 8904 8084
rect 1768 7964 1820 8016
rect 1124 7896 1176 7948
rect 1492 7896 1544 7948
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 7656 7964 7708 8016
rect 8300 7964 8352 8016
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2228 7828 2280 7880
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 5448 7896 5500 7948
rect 3516 7828 3568 7880
rect 5724 7896 5776 7948
rect 5816 7896 5868 7948
rect 1676 7760 1728 7812
rect 1768 7692 1820 7744
rect 3976 7760 4028 7812
rect 5264 7760 5316 7812
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4712 7692 4764 7744
rect 4896 7692 4948 7744
rect 5448 7692 5500 7744
rect 5724 7692 5776 7744
rect 7380 7828 7432 7880
rect 7472 7828 7524 7880
rect 8024 7896 8076 7948
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 8668 7896 8720 7948
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 8576 7828 8628 7880
rect 10048 8032 10100 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11060 8032 11112 8084
rect 12072 8032 12124 8084
rect 12992 8032 13044 8084
rect 13176 8032 13228 8084
rect 14372 8032 14424 8084
rect 15568 8032 15620 8084
rect 16580 8032 16632 8084
rect 16764 8032 16816 8084
rect 24124 8032 24176 8084
rect 24492 8032 24544 8084
rect 24676 8032 24728 8084
rect 7012 7760 7064 7812
rect 7932 7760 7984 7812
rect 8668 7760 8720 7812
rect 9312 7896 9364 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9864 7828 9916 7880
rect 9956 7828 10008 7880
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 10324 7828 10376 7880
rect 10692 7828 10744 7880
rect 12808 7964 12860 8016
rect 11796 7828 11848 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 11060 7760 11112 7812
rect 12992 7896 13044 7948
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 13360 7896 13412 7948
rect 15660 8007 15712 8016
rect 15660 7973 15669 8007
rect 15669 7973 15703 8007
rect 15703 7973 15712 8007
rect 15660 7964 15712 7973
rect 16672 7964 16724 8016
rect 17040 7964 17092 8016
rect 15292 7828 15344 7880
rect 17040 7828 17092 7880
rect 17592 7828 17644 7880
rect 17684 7828 17736 7880
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 18972 7964 19024 8016
rect 19708 8007 19760 8016
rect 19708 7973 19733 8007
rect 19733 7973 19760 8007
rect 19708 7964 19760 7973
rect 20444 8007 20496 8016
rect 18604 7896 18656 7948
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 20444 7973 20453 8007
rect 20453 7973 20487 8007
rect 20487 7973 20496 8007
rect 20444 7964 20496 7973
rect 20536 7964 20588 8016
rect 22744 7964 22796 8016
rect 23572 7964 23624 8016
rect 24952 7964 25004 8016
rect 25688 8032 25740 8084
rect 25780 8032 25832 8084
rect 28264 8032 28316 8084
rect 29092 8032 29144 8084
rect 21180 7896 21232 7948
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 19064 7828 19116 7880
rect 19156 7828 19208 7880
rect 20168 7760 20220 7812
rect 20628 7828 20680 7880
rect 20996 7828 21048 7880
rect 21916 7828 21968 7880
rect 22928 7828 22980 7880
rect 6644 7692 6696 7744
rect 7104 7692 7156 7744
rect 7380 7735 7432 7744
rect 7380 7701 7389 7735
rect 7389 7701 7423 7735
rect 7423 7701 7432 7735
rect 7380 7692 7432 7701
rect 8116 7692 8168 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9312 7692 9364 7744
rect 9864 7692 9916 7744
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11980 7692 12032 7744
rect 13452 7692 13504 7744
rect 14004 7692 14056 7744
rect 16488 7692 16540 7744
rect 20720 7692 20772 7744
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 23848 7828 23900 7880
rect 24400 7828 24452 7880
rect 25412 7939 25464 7948
rect 25412 7905 25421 7939
rect 25421 7905 25455 7939
rect 25455 7905 25464 7939
rect 25412 7896 25464 7905
rect 25872 7939 25924 7948
rect 25872 7905 25881 7939
rect 25881 7905 25915 7939
rect 25915 7905 25924 7939
rect 25872 7896 25924 7905
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 28724 7939 28776 7948
rect 28724 7905 28733 7939
rect 28733 7905 28767 7939
rect 28767 7905 28776 7939
rect 28724 7896 28776 7905
rect 25504 7828 25556 7880
rect 23112 7692 23164 7744
rect 23572 7692 23624 7744
rect 25136 7760 25188 7812
rect 25228 7692 25280 7744
rect 28080 7828 28132 7880
rect 28356 7760 28408 7812
rect 28540 7692 28592 7744
rect 4285 7590 4337 7642
rect 4349 7590 4401 7642
rect 4413 7590 4465 7642
rect 4477 7590 4529 7642
rect 4541 7590 4593 7642
rect 12059 7590 12111 7642
rect 12123 7590 12175 7642
rect 12187 7590 12239 7642
rect 12251 7590 12303 7642
rect 12315 7590 12367 7642
rect 19833 7590 19885 7642
rect 19897 7590 19949 7642
rect 19961 7590 20013 7642
rect 20025 7590 20077 7642
rect 20089 7590 20141 7642
rect 27607 7590 27659 7642
rect 27671 7590 27723 7642
rect 27735 7590 27787 7642
rect 27799 7590 27851 7642
rect 27863 7590 27915 7642
rect 3792 7488 3844 7540
rect 4896 7488 4948 7540
rect 1216 7352 1268 7404
rect 2780 7420 2832 7472
rect 2964 7420 3016 7472
rect 4804 7420 4856 7472
rect 5908 7488 5960 7540
rect 6736 7488 6788 7540
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 9312 7488 9364 7540
rect 848 7327 900 7336
rect 848 7293 857 7327
rect 857 7293 891 7327
rect 891 7293 900 7327
rect 848 7284 900 7293
rect 2228 7284 2280 7336
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 3792 7352 3844 7361
rect 4160 7284 4212 7336
rect 4804 7284 4856 7336
rect 5448 7352 5500 7404
rect 940 7148 992 7200
rect 2780 7216 2832 7268
rect 2596 7148 2648 7200
rect 3884 7148 3936 7200
rect 4528 7216 4580 7268
rect 4896 7216 4948 7268
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 4712 7148 4764 7200
rect 5632 7216 5684 7268
rect 6644 7420 6696 7472
rect 7840 7420 7892 7472
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7288 7352 7340 7404
rect 8208 7420 8260 7472
rect 8852 7420 8904 7472
rect 7564 7284 7616 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8024 7327 8076 7336
rect 8024 7293 8069 7327
rect 8069 7293 8076 7327
rect 8024 7284 8076 7293
rect 8300 7284 8352 7336
rect 6552 7148 6604 7200
rect 7472 7216 7524 7268
rect 7196 7148 7248 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 7656 7148 7708 7200
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9220 7352 9272 7404
rect 9036 7327 9088 7336
rect 9036 7293 9043 7327
rect 9043 7293 9088 7327
rect 9036 7284 9088 7293
rect 10232 7488 10284 7540
rect 10968 7488 11020 7540
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 11612 7488 11664 7540
rect 9772 7420 9824 7472
rect 11704 7420 11756 7472
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 10048 7284 10100 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11428 7352 11480 7404
rect 10876 7216 10928 7268
rect 8576 7148 8628 7200
rect 9036 7148 9088 7200
rect 9312 7148 9364 7200
rect 9956 7148 10008 7200
rect 10968 7148 11020 7200
rect 11152 7148 11204 7200
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 12440 7352 12492 7404
rect 13360 7420 13412 7472
rect 13452 7352 13504 7404
rect 15568 7463 15620 7472
rect 15568 7429 15577 7463
rect 15577 7429 15611 7463
rect 15611 7429 15620 7463
rect 15568 7420 15620 7429
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14464 7352 14516 7404
rect 12900 7216 12952 7268
rect 13360 7216 13412 7268
rect 15200 7284 15252 7336
rect 14096 7259 14148 7268
rect 14096 7225 14105 7259
rect 14105 7225 14139 7259
rect 14139 7225 14148 7259
rect 14096 7216 14148 7225
rect 15108 7148 15160 7200
rect 18052 7488 18104 7540
rect 19616 7488 19668 7540
rect 23204 7488 23256 7540
rect 23664 7488 23716 7540
rect 23756 7488 23808 7540
rect 24400 7488 24452 7540
rect 15936 7352 15988 7404
rect 16488 7420 16540 7472
rect 20812 7420 20864 7472
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 16856 7352 16908 7404
rect 17868 7352 17920 7404
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 18972 7352 19024 7404
rect 17684 7284 17736 7336
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 18512 7284 18564 7336
rect 20076 7284 20128 7336
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 16948 7148 17000 7200
rect 21548 7352 21600 7404
rect 21272 7284 21324 7336
rect 23020 7420 23072 7472
rect 21916 7327 21968 7336
rect 21916 7293 21925 7327
rect 21925 7293 21959 7327
rect 21959 7293 21968 7327
rect 21916 7284 21968 7293
rect 21640 7216 21692 7268
rect 22284 7284 22336 7336
rect 22284 7191 22336 7200
rect 22284 7157 22293 7191
rect 22293 7157 22327 7191
rect 22327 7157 22336 7191
rect 22284 7148 22336 7157
rect 22468 7284 22520 7336
rect 22652 7259 22704 7268
rect 22652 7225 22661 7259
rect 22661 7225 22695 7259
rect 22695 7225 22704 7259
rect 22652 7216 22704 7225
rect 22560 7148 22612 7200
rect 23204 7284 23256 7336
rect 23756 7284 23808 7336
rect 23848 7284 23900 7336
rect 24216 7420 24268 7472
rect 25780 7420 25832 7472
rect 29000 7488 29052 7540
rect 26332 7420 26384 7472
rect 28264 7420 28316 7472
rect 24676 7284 24728 7336
rect 25504 7395 25556 7404
rect 25504 7361 25513 7395
rect 25513 7361 25547 7395
rect 25547 7361 25556 7395
rect 25504 7352 25556 7361
rect 26516 7352 26568 7404
rect 26792 7395 26844 7404
rect 26792 7361 26801 7395
rect 26801 7361 26835 7395
rect 26835 7361 26844 7395
rect 26792 7352 26844 7361
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 23480 7148 23532 7200
rect 24124 7148 24176 7200
rect 25320 7216 25372 7268
rect 25228 7148 25280 7200
rect 26240 7284 26292 7336
rect 26700 7216 26752 7268
rect 25596 7191 25648 7200
rect 25596 7157 25605 7191
rect 25605 7157 25639 7191
rect 25639 7157 25648 7191
rect 25596 7148 25648 7157
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 26148 7148 26200 7200
rect 26884 7148 26936 7200
rect 28816 7259 28868 7268
rect 28816 7225 28825 7259
rect 28825 7225 28859 7259
rect 28859 7225 28868 7259
rect 28816 7216 28868 7225
rect 27988 7148 28040 7200
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 15946 7046 15998 7098
rect 16010 7046 16062 7098
rect 16074 7046 16126 7098
rect 16138 7046 16190 7098
rect 16202 7046 16254 7098
rect 23720 7046 23772 7098
rect 23784 7046 23836 7098
rect 23848 7046 23900 7098
rect 23912 7046 23964 7098
rect 23976 7046 24028 7098
rect 31494 7046 31546 7098
rect 31558 7046 31610 7098
rect 31622 7046 31674 7098
rect 31686 7046 31738 7098
rect 31750 7046 31802 7098
rect 1676 6944 1728 6996
rect 3424 6944 3476 6996
rect 1032 6851 1084 6860
rect 1032 6817 1041 6851
rect 1041 6817 1075 6851
rect 1075 6817 1084 6851
rect 1032 6808 1084 6817
rect 2504 6876 2556 6928
rect 3976 6944 4028 6996
rect 5264 6944 5316 6996
rect 5540 6944 5592 6996
rect 6552 6944 6604 6996
rect 7288 6944 7340 6996
rect 7472 6944 7524 6996
rect 7564 6944 7616 6996
rect 10048 6944 10100 6996
rect 10416 6944 10468 6996
rect 11244 6944 11296 6996
rect 11428 6944 11480 6996
rect 11612 6987 11664 6996
rect 11612 6953 11621 6987
rect 11621 6953 11655 6987
rect 11655 6953 11664 6987
rect 11612 6944 11664 6953
rect 11796 6944 11848 6996
rect 11980 6944 12032 6996
rect 12440 6944 12492 6996
rect 1400 6808 1452 6860
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 2780 6808 2832 6860
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 1676 6715 1728 6724
rect 1676 6681 1685 6715
rect 1685 6681 1719 6715
rect 1719 6681 1728 6715
rect 1676 6672 1728 6681
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3148 6740 3200 6792
rect 1032 6604 1084 6656
rect 3608 6672 3660 6724
rect 4528 6740 4580 6792
rect 4988 6808 5040 6860
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5816 6876 5868 6928
rect 8116 6876 8168 6928
rect 5540 6740 5592 6792
rect 5816 6740 5868 6792
rect 4804 6672 4856 6724
rect 5448 6672 5500 6724
rect 5724 6672 5776 6724
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 6920 6740 6972 6792
rect 9128 6808 9180 6860
rect 7564 6740 7616 6792
rect 8760 6740 8812 6792
rect 9036 6740 9088 6792
rect 9772 6808 9824 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 9680 6740 9732 6792
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 13452 6944 13504 6996
rect 13636 6944 13688 6996
rect 14188 6876 14240 6928
rect 15108 6876 15160 6928
rect 19432 6944 19484 6996
rect 20260 6944 20312 6996
rect 4068 6604 4120 6656
rect 5080 6604 5132 6656
rect 5264 6604 5316 6656
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7748 6604 7800 6656
rect 9496 6604 9548 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10140 6604 10192 6656
rect 11336 6740 11388 6792
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 11704 6740 11756 6792
rect 12440 6740 12492 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 12900 6740 12952 6792
rect 11428 6604 11480 6656
rect 11520 6604 11572 6656
rect 12624 6604 12676 6656
rect 13452 6604 13504 6656
rect 14188 6604 14240 6656
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14556 6740 14608 6792
rect 17500 6876 17552 6928
rect 18328 6876 18380 6928
rect 21916 6876 21968 6928
rect 14924 6740 14976 6792
rect 16488 6740 16540 6792
rect 15016 6672 15068 6724
rect 17684 6808 17736 6860
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18144 6740 18196 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18420 6740 18472 6792
rect 19800 6808 19852 6860
rect 20168 6851 20220 6860
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 20260 6808 20312 6860
rect 20536 6808 20588 6860
rect 21640 6808 21692 6860
rect 25596 6944 25648 6996
rect 22468 6876 22520 6928
rect 22928 6876 22980 6928
rect 23296 6876 23348 6928
rect 24952 6876 25004 6928
rect 17960 6672 18012 6724
rect 18880 6672 18932 6724
rect 18972 6715 19024 6724
rect 18972 6681 18981 6715
rect 18981 6681 19015 6715
rect 19015 6681 19024 6715
rect 18972 6672 19024 6681
rect 20444 6672 20496 6724
rect 21180 6672 21232 6724
rect 15200 6604 15252 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 19800 6604 19852 6656
rect 20168 6604 20220 6656
rect 22192 6672 22244 6724
rect 23572 6851 23624 6860
rect 23572 6817 23581 6851
rect 23581 6817 23615 6851
rect 23615 6817 23624 6851
rect 23572 6808 23624 6817
rect 24124 6851 24176 6860
rect 24124 6817 24133 6851
rect 24133 6817 24167 6851
rect 24167 6817 24176 6851
rect 24124 6808 24176 6817
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 24308 6808 24360 6860
rect 24492 6808 24544 6860
rect 25412 6876 25464 6928
rect 26332 6944 26384 6996
rect 26640 6987 26692 6996
rect 26640 6953 26651 6987
rect 26651 6953 26692 6987
rect 26640 6944 26692 6953
rect 28080 6944 28132 6996
rect 29000 6944 29052 6996
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 23480 6672 23532 6724
rect 26148 6808 26200 6860
rect 26240 6808 26292 6860
rect 28540 6876 28592 6928
rect 26792 6808 26844 6860
rect 28264 6808 28316 6860
rect 25136 6740 25188 6792
rect 25504 6740 25556 6792
rect 25872 6740 25924 6792
rect 26332 6740 26384 6792
rect 24768 6672 24820 6724
rect 24676 6604 24728 6656
rect 26148 6604 26200 6656
rect 26240 6647 26292 6656
rect 26240 6613 26249 6647
rect 26249 6613 26283 6647
rect 26283 6613 26292 6647
rect 26240 6604 26292 6613
rect 26332 6604 26384 6656
rect 27160 6604 27212 6656
rect 28632 6647 28684 6656
rect 28632 6613 28641 6647
rect 28641 6613 28675 6647
rect 28675 6613 28684 6647
rect 28632 6604 28684 6613
rect 4285 6502 4337 6554
rect 4349 6502 4401 6554
rect 4413 6502 4465 6554
rect 4477 6502 4529 6554
rect 4541 6502 4593 6554
rect 12059 6502 12111 6554
rect 12123 6502 12175 6554
rect 12187 6502 12239 6554
rect 12251 6502 12303 6554
rect 12315 6502 12367 6554
rect 19833 6502 19885 6554
rect 19897 6502 19949 6554
rect 19961 6502 20013 6554
rect 20025 6502 20077 6554
rect 20089 6502 20141 6554
rect 27607 6502 27659 6554
rect 27671 6502 27723 6554
rect 27735 6502 27787 6554
rect 27799 6502 27851 6554
rect 27863 6502 27915 6554
rect 1400 6400 1452 6452
rect 2964 6400 3016 6452
rect 4252 6400 4304 6452
rect 5356 6400 5408 6452
rect 5540 6400 5592 6452
rect 848 6307 900 6316
rect 848 6273 857 6307
rect 857 6273 891 6307
rect 891 6273 900 6307
rect 4068 6332 4120 6384
rect 7288 6400 7340 6452
rect 8484 6400 8536 6452
rect 8576 6400 8628 6452
rect 9496 6400 9548 6452
rect 9864 6400 9916 6452
rect 8852 6332 8904 6384
rect 848 6264 900 6273
rect 1216 6239 1268 6248
rect 1216 6205 1225 6239
rect 1225 6205 1259 6239
rect 1259 6205 1268 6239
rect 1216 6196 1268 6205
rect 2044 6196 2096 6248
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 6920 6264 6972 6316
rect 2228 6128 2280 6180
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 2872 6060 2924 6112
rect 3976 6128 4028 6180
rect 4620 6196 4672 6248
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 5172 6196 5224 6248
rect 5632 6196 5684 6248
rect 7196 6196 7248 6248
rect 4160 6060 4212 6112
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 7564 6264 7616 6316
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 8024 6239 8076 6248
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 8576 6264 8628 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9680 6264 9732 6316
rect 9220 6196 9272 6248
rect 10232 6264 10284 6316
rect 11520 6400 11572 6452
rect 11980 6400 12032 6452
rect 12992 6400 13044 6452
rect 14096 6400 14148 6452
rect 14372 6400 14424 6452
rect 14740 6443 14792 6452
rect 14740 6409 14749 6443
rect 14749 6409 14783 6443
rect 14783 6409 14792 6443
rect 14740 6400 14792 6409
rect 15752 6400 15804 6452
rect 11888 6332 11940 6384
rect 17684 6400 17736 6452
rect 17776 6400 17828 6452
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 18052 6400 18104 6452
rect 18604 6400 18656 6452
rect 11244 6264 11296 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 14188 6264 14240 6316
rect 14556 6264 14608 6316
rect 15016 6264 15068 6316
rect 16672 6264 16724 6316
rect 13084 6196 13136 6248
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 8024 6060 8076 6112
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 9496 6060 9548 6112
rect 10692 6128 10744 6180
rect 11336 6128 11388 6180
rect 12624 6128 12676 6180
rect 14004 6196 14056 6248
rect 14280 6196 14332 6248
rect 15108 6196 15160 6248
rect 15384 6171 15436 6180
rect 15384 6137 15393 6171
rect 15393 6137 15427 6171
rect 15427 6137 15436 6171
rect 15384 6128 15436 6137
rect 15568 6171 15620 6180
rect 15568 6137 15577 6171
rect 15577 6137 15611 6171
rect 15611 6137 15620 6171
rect 15568 6128 15620 6137
rect 18144 6332 18196 6384
rect 19708 6332 19760 6384
rect 21180 6400 21232 6452
rect 21272 6332 21324 6384
rect 21364 6332 21416 6384
rect 25872 6400 25924 6452
rect 26240 6400 26292 6452
rect 28172 6400 28224 6452
rect 28356 6400 28408 6452
rect 28632 6400 28684 6452
rect 17040 6128 17092 6180
rect 13636 6060 13688 6112
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 16304 6060 16356 6112
rect 16488 6060 16540 6112
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 18512 6196 18564 6248
rect 18236 6171 18288 6180
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 18236 6128 18288 6137
rect 18328 6128 18380 6180
rect 19248 6128 19300 6180
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 19800 6239 19852 6248
rect 19800 6205 19809 6239
rect 19809 6205 19843 6239
rect 19843 6205 19852 6239
rect 19800 6196 19852 6205
rect 20260 6264 20312 6316
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 21732 6264 21784 6316
rect 22468 6264 22520 6316
rect 19984 6196 20036 6205
rect 21088 6196 21140 6248
rect 25136 6332 25188 6384
rect 25964 6332 26016 6384
rect 20076 6128 20128 6180
rect 20536 6128 20588 6180
rect 21824 6239 21876 6248
rect 21824 6205 21833 6239
rect 21833 6205 21867 6239
rect 21867 6205 21876 6239
rect 21824 6196 21876 6205
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22100 6196 22152 6248
rect 24032 6239 24084 6248
rect 21640 6128 21692 6180
rect 22836 6128 22888 6180
rect 22192 6060 22244 6112
rect 22468 6060 22520 6112
rect 24032 6205 24036 6239
rect 24036 6205 24070 6239
rect 24070 6205 24084 6239
rect 24032 6196 24084 6205
rect 24400 6239 24452 6248
rect 24400 6205 24408 6239
rect 24408 6205 24442 6239
rect 24442 6205 24452 6239
rect 24400 6196 24452 6205
rect 24768 6264 24820 6316
rect 24676 6196 24728 6248
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 24124 6171 24176 6180
rect 24124 6137 24133 6171
rect 24133 6137 24167 6171
rect 24167 6137 24176 6171
rect 24124 6128 24176 6137
rect 25136 6196 25188 6248
rect 25320 6196 25372 6248
rect 25596 6239 25648 6248
rect 25596 6205 25605 6239
rect 25605 6205 25639 6239
rect 25639 6205 25648 6239
rect 25596 6196 25648 6205
rect 25688 6239 25740 6248
rect 25688 6205 25697 6239
rect 25697 6205 25731 6239
rect 25731 6205 25740 6239
rect 25688 6196 25740 6205
rect 25780 6239 25832 6248
rect 25780 6205 25789 6239
rect 25789 6205 25823 6239
rect 25823 6205 25832 6239
rect 25780 6196 25832 6205
rect 25136 6060 25188 6112
rect 25320 6103 25372 6112
rect 25320 6069 25329 6103
rect 25329 6069 25363 6103
rect 25363 6069 25372 6103
rect 25320 6060 25372 6069
rect 25596 6060 25648 6112
rect 26700 6239 26752 6248
rect 26700 6205 26709 6239
rect 26709 6205 26743 6239
rect 26743 6205 26752 6239
rect 26700 6196 26752 6205
rect 27160 6239 27212 6248
rect 27160 6205 27169 6239
rect 27169 6205 27203 6239
rect 27203 6205 27212 6239
rect 27160 6196 27212 6205
rect 27344 6196 27396 6248
rect 28080 6239 28132 6248
rect 28080 6205 28089 6239
rect 28089 6205 28123 6239
rect 28123 6205 28132 6239
rect 28080 6196 28132 6205
rect 27620 6128 27672 6180
rect 27988 6171 28040 6180
rect 27988 6137 27997 6171
rect 27997 6137 28031 6171
rect 28031 6137 28040 6171
rect 27988 6128 28040 6137
rect 28356 6171 28408 6180
rect 28356 6137 28365 6171
rect 28365 6137 28399 6171
rect 28399 6137 28408 6171
rect 28356 6128 28408 6137
rect 28724 6196 28776 6248
rect 29368 6239 29420 6248
rect 29368 6205 29377 6239
rect 29377 6205 29411 6239
rect 29411 6205 29420 6239
rect 29368 6196 29420 6205
rect 26240 6060 26292 6112
rect 26608 6060 26660 6112
rect 26976 6060 27028 6112
rect 29000 6060 29052 6112
rect 29644 6060 29696 6112
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 15946 5958 15998 6010
rect 16010 5958 16062 6010
rect 16074 5958 16126 6010
rect 16138 5958 16190 6010
rect 16202 5958 16254 6010
rect 23720 5958 23772 6010
rect 23784 5958 23836 6010
rect 23848 5958 23900 6010
rect 23912 5958 23964 6010
rect 23976 5958 24028 6010
rect 31494 5958 31546 6010
rect 31558 5958 31610 6010
rect 31622 5958 31674 6010
rect 31686 5958 31738 6010
rect 31750 5958 31802 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 756 5788 808 5840
rect 1952 5856 2004 5908
rect 1860 5831 1912 5840
rect 1860 5797 1869 5831
rect 1869 5797 1903 5831
rect 1903 5797 1912 5831
rect 1860 5788 1912 5797
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2872 5856 2924 5908
rect 3792 5856 3844 5908
rect 4804 5856 4856 5908
rect 5172 5856 5224 5908
rect 6000 5856 6052 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 6920 5856 6972 5908
rect 7380 5856 7432 5908
rect 7656 5856 7708 5908
rect 8576 5856 8628 5908
rect 8760 5856 8812 5908
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 13636 5856 13688 5908
rect 2044 5652 2096 5704
rect 2688 5720 2740 5772
rect 4068 5720 4120 5772
rect 4252 5720 4304 5772
rect 4620 5720 4672 5772
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6000 5720 6052 5772
rect 2780 5652 2832 5704
rect 3884 5652 3936 5704
rect 6184 5720 6236 5772
rect 7012 5763 7064 5772
rect 7012 5729 7021 5763
rect 7021 5729 7055 5763
rect 7055 5729 7064 5763
rect 7012 5720 7064 5729
rect 9404 5788 9456 5840
rect 8760 5720 8812 5772
rect 10232 5720 10284 5772
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 10692 5788 10744 5840
rect 12900 5788 12952 5840
rect 10876 5720 10928 5772
rect 1124 5584 1176 5636
rect 4988 5584 5040 5636
rect 6092 5584 6144 5636
rect 7472 5652 7524 5704
rect 12992 5720 13044 5772
rect 11336 5652 11388 5704
rect 13452 5652 13504 5704
rect 14372 5720 14424 5772
rect 14464 5720 14516 5772
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 14924 5856 14976 5908
rect 18236 5856 18288 5908
rect 15844 5788 15896 5840
rect 17040 5720 17092 5772
rect 16120 5695 16172 5704
rect 3792 5516 3844 5568
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 4896 5559 4948 5568
rect 4896 5525 4905 5559
rect 4905 5525 4939 5559
rect 4939 5525 4948 5559
rect 4896 5516 4948 5525
rect 7748 5516 7800 5568
rect 7932 5516 7984 5568
rect 8576 5516 8628 5568
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 10968 5584 11020 5636
rect 12808 5584 12860 5636
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16304 5652 16356 5704
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 18052 5652 18104 5704
rect 18236 5720 18288 5772
rect 18880 5788 18932 5840
rect 19800 5856 19852 5908
rect 19984 5788 20036 5840
rect 21180 5856 21232 5908
rect 22376 5856 22428 5908
rect 22928 5899 22980 5908
rect 22928 5865 22937 5899
rect 22937 5865 22971 5899
rect 22971 5865 22980 5899
rect 22928 5856 22980 5865
rect 23204 5856 23256 5908
rect 20536 5831 20588 5840
rect 20536 5797 20545 5831
rect 20545 5797 20579 5831
rect 20579 5797 20588 5831
rect 20536 5788 20588 5797
rect 19524 5763 19576 5772
rect 19524 5729 19566 5763
rect 19566 5729 19576 5763
rect 19524 5720 19576 5729
rect 20076 5763 20128 5772
rect 20076 5729 20085 5763
rect 20085 5729 20119 5763
rect 20119 5729 20128 5763
rect 20076 5720 20128 5729
rect 20260 5720 20312 5772
rect 20628 5720 20680 5772
rect 20904 5720 20956 5772
rect 19708 5652 19760 5704
rect 21088 5652 21140 5704
rect 21640 5763 21692 5772
rect 21640 5729 21649 5763
rect 21649 5729 21683 5763
rect 21683 5729 21692 5763
rect 21640 5720 21692 5729
rect 21732 5720 21784 5772
rect 21824 5720 21876 5772
rect 24124 5788 24176 5840
rect 22560 5720 22612 5772
rect 22836 5720 22888 5772
rect 23480 5720 23532 5772
rect 23572 5720 23624 5772
rect 24492 5856 24544 5908
rect 25136 5856 25188 5908
rect 25228 5856 25280 5908
rect 14280 5516 14332 5568
rect 14556 5516 14608 5568
rect 15016 5516 15068 5568
rect 18972 5584 19024 5636
rect 19432 5559 19484 5568
rect 19432 5525 19441 5559
rect 19441 5525 19475 5559
rect 19475 5525 19484 5559
rect 19432 5516 19484 5525
rect 21916 5627 21968 5636
rect 21916 5593 21925 5627
rect 21925 5593 21959 5627
rect 21959 5593 21968 5627
rect 21916 5584 21968 5593
rect 20260 5516 20312 5568
rect 20536 5516 20588 5568
rect 22284 5584 22336 5636
rect 23204 5652 23256 5704
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 24308 5695 24360 5704
rect 24308 5661 24317 5695
rect 24317 5661 24351 5695
rect 24351 5661 24360 5695
rect 24308 5652 24360 5661
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24860 5763 24912 5772
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 24952 5652 25004 5704
rect 25228 5720 25280 5772
rect 25596 5720 25648 5772
rect 26240 5856 26292 5908
rect 26424 5856 26476 5908
rect 25964 5720 26016 5772
rect 26148 5720 26200 5772
rect 26976 5720 27028 5772
rect 28080 5788 28132 5840
rect 28816 5856 28868 5908
rect 29368 5856 29420 5908
rect 28448 5720 28500 5772
rect 22836 5516 22888 5568
rect 23112 5559 23164 5568
rect 23112 5525 23121 5559
rect 23121 5525 23155 5559
rect 23155 5525 23164 5559
rect 23112 5516 23164 5525
rect 23572 5516 23624 5568
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 25044 5516 25096 5568
rect 25504 5516 25556 5568
rect 26516 5652 26568 5704
rect 27068 5652 27120 5704
rect 26608 5584 26660 5636
rect 26700 5584 26752 5636
rect 29000 5652 29052 5704
rect 29092 5584 29144 5636
rect 25964 5516 26016 5568
rect 26056 5516 26108 5568
rect 26516 5516 26568 5568
rect 28448 5516 28500 5568
rect 28632 5516 28684 5568
rect 29644 5763 29696 5772
rect 29644 5729 29653 5763
rect 29653 5729 29687 5763
rect 29687 5729 29696 5763
rect 29644 5720 29696 5729
rect 29552 5559 29604 5568
rect 29552 5525 29561 5559
rect 29561 5525 29595 5559
rect 29595 5525 29604 5559
rect 29552 5516 29604 5525
rect 4285 5414 4337 5466
rect 4349 5414 4401 5466
rect 4413 5414 4465 5466
rect 4477 5414 4529 5466
rect 4541 5414 4593 5466
rect 12059 5414 12111 5466
rect 12123 5414 12175 5466
rect 12187 5414 12239 5466
rect 12251 5414 12303 5466
rect 12315 5414 12367 5466
rect 19833 5414 19885 5466
rect 19897 5414 19949 5466
rect 19961 5414 20013 5466
rect 20025 5414 20077 5466
rect 20089 5414 20141 5466
rect 27607 5414 27659 5466
rect 27671 5414 27723 5466
rect 27735 5414 27787 5466
rect 27799 5414 27851 5466
rect 27863 5414 27915 5466
rect 848 5219 900 5228
rect 848 5185 857 5219
rect 857 5185 891 5219
rect 891 5185 900 5219
rect 848 5176 900 5185
rect 2320 5176 2372 5228
rect 2412 5108 2464 5160
rect 4804 5312 4856 5364
rect 6828 5312 6880 5364
rect 2872 5244 2924 5296
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4160 5176 4212 5228
rect 7564 5312 7616 5364
rect 7840 5312 7892 5364
rect 9496 5312 9548 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 16764 5312 16816 5364
rect 10968 5244 11020 5296
rect 4804 5176 4856 5228
rect 9220 5176 9272 5228
rect 1124 5083 1176 5092
rect 1124 5049 1133 5083
rect 1133 5049 1167 5083
rect 1167 5049 1176 5083
rect 1124 5040 1176 5049
rect 2412 4972 2464 5024
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 6000 5108 6052 5160
rect 4712 5083 4764 5092
rect 4712 5049 4721 5083
rect 4721 5049 4755 5083
rect 4755 5049 4764 5083
rect 4712 5040 4764 5049
rect 3332 4972 3384 5024
rect 4068 4972 4120 5024
rect 6184 5040 6236 5092
rect 7196 5040 7248 5092
rect 7840 5040 7892 5092
rect 8024 5040 8076 5092
rect 8852 5083 8904 5092
rect 8852 5049 8861 5083
rect 8861 5049 8895 5083
rect 8895 5049 8904 5083
rect 8852 5040 8904 5049
rect 10324 5040 10376 5092
rect 11520 5176 11572 5228
rect 13360 5287 13412 5296
rect 13360 5253 13369 5287
rect 13369 5253 13403 5287
rect 13403 5253 13412 5287
rect 13360 5244 13412 5253
rect 14188 5287 14240 5296
rect 14188 5253 14197 5287
rect 14197 5253 14231 5287
rect 14231 5253 14240 5287
rect 14188 5244 14240 5253
rect 12532 5176 12584 5228
rect 12900 5108 12952 5160
rect 11796 5040 11848 5092
rect 11152 4972 11204 5024
rect 14648 5244 14700 5296
rect 16120 5244 16172 5296
rect 16856 5244 16908 5296
rect 14096 5151 14148 5160
rect 14096 5117 14105 5151
rect 14105 5117 14139 5151
rect 14139 5117 14148 5151
rect 14096 5108 14148 5117
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 14924 5108 14976 5160
rect 15292 5176 15344 5228
rect 15752 5108 15804 5160
rect 14004 4972 14056 5024
rect 15384 4972 15436 5024
rect 16212 5108 16264 5160
rect 17132 5176 17184 5228
rect 17040 5108 17092 5160
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 18420 5176 18472 5228
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 19616 5355 19668 5364
rect 19616 5321 19625 5355
rect 19625 5321 19659 5355
rect 19659 5321 19668 5355
rect 19616 5312 19668 5321
rect 21732 5312 21784 5364
rect 22284 5312 22336 5364
rect 19708 5244 19760 5296
rect 19432 5176 19484 5228
rect 21088 5244 21140 5296
rect 21640 5244 21692 5296
rect 16488 4972 16540 5024
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 19340 5040 19392 5092
rect 19248 4972 19300 5024
rect 19708 5108 19760 5160
rect 22100 5176 22152 5228
rect 24216 5312 24268 5364
rect 24952 5312 25004 5364
rect 25780 5312 25832 5364
rect 25964 5312 26016 5364
rect 26516 5312 26568 5364
rect 26700 5312 26752 5364
rect 23020 5244 23072 5296
rect 20260 5040 20312 5092
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 23296 5176 23348 5228
rect 24400 5244 24452 5296
rect 24768 5287 24820 5296
rect 24768 5253 24777 5287
rect 24777 5253 24811 5287
rect 24811 5253 24820 5287
rect 24768 5244 24820 5253
rect 22376 5108 22428 5117
rect 20444 4972 20496 5024
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 21732 4972 21784 5024
rect 21824 4972 21876 5024
rect 22468 5015 22520 5024
rect 22468 4981 22477 5015
rect 22477 4981 22511 5015
rect 22511 4981 22520 5015
rect 22468 4972 22520 4981
rect 22836 5108 22888 5160
rect 22928 5108 22980 5160
rect 23204 5040 23256 5092
rect 23388 5040 23440 5092
rect 23848 5083 23900 5092
rect 23848 5049 23857 5083
rect 23857 5049 23891 5083
rect 23891 5049 23900 5083
rect 23848 5040 23900 5049
rect 24400 5083 24452 5092
rect 24400 5049 24409 5083
rect 24409 5049 24443 5083
rect 24443 5049 24452 5083
rect 24400 5040 24452 5049
rect 28632 5312 28684 5364
rect 25412 5151 25464 5160
rect 25412 5117 25421 5151
rect 25421 5117 25455 5151
rect 25455 5117 25464 5151
rect 25412 5108 25464 5117
rect 26608 5151 26660 5160
rect 26608 5117 26617 5151
rect 26617 5117 26651 5151
rect 26651 5117 26660 5151
rect 26608 5108 26660 5117
rect 23940 4972 23992 5024
rect 25964 5083 26016 5092
rect 25964 5049 25973 5083
rect 25973 5049 26007 5083
rect 26007 5049 26016 5083
rect 25964 5040 26016 5049
rect 26700 5040 26752 5092
rect 27344 5040 27396 5092
rect 28080 5176 28132 5228
rect 28356 5108 28408 5160
rect 28080 5083 28132 5092
rect 28080 5049 28089 5083
rect 28089 5049 28123 5083
rect 28123 5049 28132 5083
rect 28080 5040 28132 5049
rect 29092 5108 29144 5160
rect 29552 5108 29604 5160
rect 26976 4972 27028 5024
rect 27160 4972 27212 5024
rect 27620 5015 27672 5024
rect 27620 4981 27629 5015
rect 27629 4981 27663 5015
rect 27663 4981 27672 5015
rect 27620 4972 27672 4981
rect 28264 4972 28316 5024
rect 29644 5015 29696 5024
rect 29644 4981 29653 5015
rect 29653 4981 29687 5015
rect 29687 4981 29696 5015
rect 29644 4972 29696 4981
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 15946 4870 15998 4922
rect 16010 4870 16062 4922
rect 16074 4870 16126 4922
rect 16138 4870 16190 4922
rect 16202 4870 16254 4922
rect 23720 4870 23772 4922
rect 23784 4870 23836 4922
rect 23848 4870 23900 4922
rect 23912 4870 23964 4922
rect 23976 4870 24028 4922
rect 31494 4870 31546 4922
rect 31558 4870 31610 4922
rect 31622 4870 31674 4922
rect 31686 4870 31738 4922
rect 31750 4870 31802 4922
rect 1032 4768 1084 4820
rect 1216 4768 1268 4820
rect 1676 4768 1728 4820
rect 2596 4768 2648 4820
rect 2872 4768 2924 4820
rect 4620 4768 4672 4820
rect 2136 4700 2188 4752
rect 2412 4632 2464 4684
rect 2688 4700 2740 4752
rect 4068 4700 4120 4752
rect 5264 4811 5316 4820
rect 5264 4777 5273 4811
rect 5273 4777 5307 4811
rect 5307 4777 5316 4811
rect 5264 4768 5316 4777
rect 940 4496 992 4548
rect 1032 4496 1084 4548
rect 3332 4564 3384 4616
rect 6000 4700 6052 4752
rect 5816 4632 5868 4684
rect 7472 4768 7524 4820
rect 7564 4768 7616 4820
rect 8944 4768 8996 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 10968 4768 11020 4820
rect 11888 4768 11940 4820
rect 6552 4700 6604 4752
rect 7196 4700 7248 4752
rect 9220 4700 9272 4752
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 10784 4632 10836 4684
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 12624 4632 12676 4684
rect 14096 4768 14148 4820
rect 14740 4768 14792 4820
rect 13912 4743 13964 4752
rect 13912 4709 13921 4743
rect 13921 4709 13955 4743
rect 13955 4709 13964 4743
rect 13912 4700 13964 4709
rect 15200 4768 15252 4820
rect 15292 4768 15344 4820
rect 15384 4768 15436 4820
rect 15476 4768 15528 4820
rect 14464 4675 14516 4684
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 3884 4496 3936 4548
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7012 4564 7064 4616
rect 8760 4496 8812 4548
rect 12992 4539 13044 4548
rect 12992 4505 13001 4539
rect 13001 4505 13035 4539
rect 13035 4505 13044 4539
rect 12992 4496 13044 4505
rect 13084 4539 13136 4548
rect 13084 4505 13093 4539
rect 13093 4505 13127 4539
rect 13127 4505 13136 4539
rect 13084 4496 13136 4505
rect 13176 4496 13228 4548
rect 2596 4428 2648 4480
rect 4620 4428 4672 4480
rect 6184 4428 6236 4480
rect 7012 4428 7064 4480
rect 9404 4428 9456 4480
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16764 4768 16816 4820
rect 16856 4768 16908 4820
rect 17132 4768 17184 4820
rect 17776 4768 17828 4820
rect 18052 4768 18104 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18328 4768 18380 4820
rect 21824 4768 21876 4820
rect 21916 4768 21968 4820
rect 17224 4700 17276 4752
rect 15108 4564 15160 4616
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 15568 4496 15620 4548
rect 15660 4496 15712 4548
rect 18144 4496 18196 4548
rect 16580 4428 16632 4480
rect 16672 4471 16724 4480
rect 16672 4437 16681 4471
rect 16681 4437 16715 4471
rect 16715 4437 16724 4471
rect 16672 4428 16724 4437
rect 17040 4428 17092 4480
rect 17776 4471 17828 4480
rect 17776 4437 17785 4471
rect 17785 4437 17819 4471
rect 17819 4437 17828 4471
rect 17776 4428 17828 4437
rect 18788 4428 18840 4480
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 19340 4632 19392 4684
rect 20444 4675 20496 4684
rect 20444 4641 20448 4675
rect 20448 4641 20482 4675
rect 20482 4641 20496 4675
rect 20444 4632 20496 4641
rect 21180 4700 21232 4752
rect 21732 4743 21784 4752
rect 21732 4709 21741 4743
rect 21741 4709 21775 4743
rect 21775 4709 21784 4743
rect 21732 4700 21784 4709
rect 20812 4675 20864 4684
rect 20812 4641 20820 4675
rect 20820 4641 20854 4675
rect 20854 4641 20864 4675
rect 20812 4632 20864 4641
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 19156 4496 19208 4548
rect 19432 4428 19484 4480
rect 21364 4496 21416 4548
rect 21824 4496 21876 4548
rect 22284 4632 22336 4684
rect 23020 4768 23072 4820
rect 23112 4768 23164 4820
rect 23572 4768 23624 4820
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 24400 4768 24452 4820
rect 25136 4768 25188 4820
rect 22560 4700 22612 4752
rect 22836 4632 22888 4684
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 22928 4632 22980 4641
rect 25228 4700 25280 4752
rect 25780 4768 25832 4820
rect 26332 4768 26384 4820
rect 24492 4632 24544 4684
rect 25136 4632 25188 4684
rect 26516 4700 26568 4752
rect 26884 4700 26936 4752
rect 25320 4564 25372 4616
rect 25688 4675 25740 4684
rect 25688 4641 25697 4675
rect 25697 4641 25731 4675
rect 25731 4641 25740 4675
rect 25688 4632 25740 4641
rect 26332 4632 26384 4684
rect 26792 4632 26844 4684
rect 23204 4496 23256 4548
rect 25596 4496 25648 4548
rect 26332 4496 26384 4548
rect 26516 4496 26568 4548
rect 27528 4496 27580 4548
rect 23388 4428 23440 4480
rect 23848 4428 23900 4480
rect 25412 4471 25464 4480
rect 25412 4437 25421 4471
rect 25421 4437 25455 4471
rect 25455 4437 25464 4471
rect 25412 4428 25464 4437
rect 25504 4428 25556 4480
rect 26240 4428 26292 4480
rect 26700 4428 26752 4480
rect 26976 4428 27028 4480
rect 29644 4428 29696 4480
rect 4285 4326 4337 4378
rect 4349 4326 4401 4378
rect 4413 4326 4465 4378
rect 4477 4326 4529 4378
rect 4541 4326 4593 4378
rect 12059 4326 12111 4378
rect 12123 4326 12175 4378
rect 12187 4326 12239 4378
rect 12251 4326 12303 4378
rect 12315 4326 12367 4378
rect 19833 4326 19885 4378
rect 19897 4326 19949 4378
rect 19961 4326 20013 4378
rect 20025 4326 20077 4378
rect 20089 4326 20141 4378
rect 27607 4326 27659 4378
rect 27671 4326 27723 4378
rect 27735 4326 27787 4378
rect 27799 4326 27851 4378
rect 27863 4326 27915 4378
rect 1124 4224 1176 4276
rect 4620 4224 4672 4276
rect 6736 4224 6788 4276
rect 7196 4224 7248 4276
rect 7472 4224 7524 4276
rect 8852 4224 8904 4276
rect 9588 4224 9640 4276
rect 10416 4224 10468 4276
rect 10968 4224 11020 4276
rect 14280 4224 14332 4276
rect 15660 4267 15712 4276
rect 15660 4233 15669 4267
rect 15669 4233 15703 4267
rect 15703 4233 15712 4267
rect 15660 4224 15712 4233
rect 16028 4224 16080 4276
rect 19708 4224 19760 4276
rect 2780 4156 2832 4208
rect 3884 4156 3936 4208
rect 1032 4088 1084 4140
rect 2044 4088 2096 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3240 4088 3292 4140
rect 2412 4020 2464 4072
rect 1400 3995 1452 4004
rect 1400 3961 1409 3995
rect 1409 3961 1443 3995
rect 1443 3961 1452 3995
rect 1400 3952 1452 3961
rect 2780 4020 2832 4072
rect 3056 4020 3108 4072
rect 6092 4088 6144 4140
rect 4068 4020 4120 4072
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5908 4020 5960 4072
rect 7564 4088 7616 4140
rect 7104 4020 7156 4072
rect 8576 4088 8628 4140
rect 9312 4156 9364 4208
rect 14004 4156 14056 4208
rect 9220 4088 9272 4140
rect 10600 4088 10652 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12992 4088 13044 4140
rect 13544 4088 13596 4140
rect 4896 3952 4948 4004
rect 6184 3952 6236 4004
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 3332 3884 3384 3936
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 8760 3952 8812 4004
rect 9036 3995 9088 4004
rect 9036 3961 9045 3995
rect 9045 3961 9079 3995
rect 9079 3961 9088 3995
rect 9036 3952 9088 3961
rect 9772 3995 9824 4004
rect 9772 3961 9781 3995
rect 9781 3961 9815 3995
rect 9815 3961 9824 3995
rect 9772 3952 9824 3961
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9496 3884 9548 3936
rect 15016 4156 15068 4208
rect 18236 4156 18288 4208
rect 10508 3952 10560 4004
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 11612 3952 11664 4004
rect 13820 3952 13872 4004
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 15200 3995 15252 4004
rect 15200 3961 15209 3995
rect 15209 3961 15243 3995
rect 15243 3961 15252 3995
rect 15200 3952 15252 3961
rect 13544 3884 13596 3936
rect 14464 3884 14516 3936
rect 15108 3884 15160 3936
rect 16304 4088 16356 4140
rect 16672 4088 16724 4140
rect 16028 4020 16080 4072
rect 16212 3952 16264 4004
rect 17316 4020 17368 4072
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 18788 4020 18840 4072
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 20536 4156 20588 4208
rect 19616 4088 19668 4140
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 19708 4020 19760 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 20260 4020 20312 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 20444 4063 20496 4072
rect 20444 4029 20453 4063
rect 20453 4029 20487 4063
rect 20487 4029 20496 4063
rect 20444 4020 20496 4029
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 21272 4063 21324 4072
rect 21272 4029 21286 4063
rect 21286 4029 21320 4063
rect 21320 4029 21324 4063
rect 21272 4020 21324 4029
rect 21824 4020 21876 4072
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 22928 4224 22980 4276
rect 22468 4156 22520 4208
rect 23204 4156 23256 4208
rect 23480 4199 23532 4208
rect 23480 4165 23489 4199
rect 23489 4165 23523 4199
rect 23523 4165 23532 4199
rect 23480 4156 23532 4165
rect 24124 4267 24176 4276
rect 24124 4233 24133 4267
rect 24133 4233 24167 4267
rect 24167 4233 24176 4267
rect 24124 4224 24176 4233
rect 25872 4267 25924 4276
rect 25872 4233 25881 4267
rect 25881 4233 25915 4267
rect 25915 4233 25924 4267
rect 25872 4224 25924 4233
rect 16672 3884 16724 3936
rect 17132 3884 17184 3936
rect 19432 3884 19484 3936
rect 19708 3884 19760 3936
rect 20260 3884 20312 3936
rect 21456 3927 21508 3936
rect 21456 3893 21465 3927
rect 21465 3893 21499 3927
rect 21499 3893 21508 3927
rect 21456 3884 21508 3893
rect 21548 3927 21600 3936
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 21824 3884 21876 3936
rect 22284 3884 22336 3936
rect 23020 3884 23072 3936
rect 23296 4020 23348 4072
rect 24676 4156 24728 4208
rect 25320 4088 25372 4140
rect 24860 4020 24912 4072
rect 25136 4020 25188 4072
rect 25504 4063 25556 4072
rect 25504 4029 25513 4063
rect 25513 4029 25547 4063
rect 25547 4029 25556 4063
rect 25504 4020 25556 4029
rect 26424 4088 26476 4140
rect 26516 4063 26568 4072
rect 23572 3884 23624 3936
rect 23756 3884 23808 3936
rect 25596 3995 25648 4004
rect 25596 3961 25605 3995
rect 25605 3961 25639 3995
rect 25639 3961 25648 3995
rect 25596 3952 25648 3961
rect 24768 3927 24820 3936
rect 24768 3893 24777 3927
rect 24777 3893 24811 3927
rect 24811 3893 24820 3927
rect 24768 3884 24820 3893
rect 26516 4029 26520 4063
rect 26520 4029 26554 4063
rect 26554 4029 26568 4063
rect 26516 4020 26568 4029
rect 26884 4063 26936 4072
rect 26884 4029 26892 4063
rect 26892 4029 26926 4063
rect 26926 4029 26936 4063
rect 26884 4020 26936 4029
rect 26976 4063 27028 4072
rect 26976 4029 26985 4063
rect 26985 4029 27019 4063
rect 27019 4029 27028 4063
rect 26976 4020 27028 4029
rect 27068 4063 27120 4072
rect 27068 4029 27077 4063
rect 27077 4029 27111 4063
rect 27111 4029 27120 4063
rect 27068 4020 27120 4029
rect 27160 4063 27212 4072
rect 27160 4029 27169 4063
rect 27169 4029 27203 4063
rect 27203 4029 27212 4063
rect 27160 4020 27212 4029
rect 27252 4020 27304 4072
rect 26700 3995 26752 4004
rect 26700 3961 26709 3995
rect 26709 3961 26743 3995
rect 26743 3961 26752 3995
rect 26700 3952 26752 3961
rect 27528 3952 27580 4004
rect 27988 4020 28040 4072
rect 28080 3952 28132 4004
rect 28172 3995 28224 4004
rect 28172 3961 28181 3995
rect 28181 3961 28215 3995
rect 28215 3961 28224 3995
rect 28172 3952 28224 3961
rect 26884 3884 26936 3936
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 15946 3782 15998 3834
rect 16010 3782 16062 3834
rect 16074 3782 16126 3834
rect 16138 3782 16190 3834
rect 16202 3782 16254 3834
rect 23720 3782 23772 3834
rect 23784 3782 23836 3834
rect 23848 3782 23900 3834
rect 23912 3782 23964 3834
rect 23976 3782 24028 3834
rect 31494 3782 31546 3834
rect 31558 3782 31610 3834
rect 31622 3782 31674 3834
rect 31686 3782 31738 3834
rect 31750 3782 31802 3834
rect 2044 3680 2096 3732
rect 4528 3680 4580 3732
rect 4804 3680 4856 3732
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 4068 3612 4120 3664
rect 4252 3612 4304 3664
rect 5908 3612 5960 3664
rect 6184 3612 6236 3664
rect 3884 3587 3936 3596
rect 3884 3553 3893 3587
rect 3893 3553 3927 3587
rect 3927 3553 3936 3587
rect 3884 3544 3936 3553
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 6828 3680 6880 3732
rect 9220 3680 9272 3732
rect 9312 3680 9364 3732
rect 7012 3612 7064 3664
rect 8392 3655 8444 3664
rect 8392 3621 8401 3655
rect 8401 3621 8435 3655
rect 8435 3621 8444 3655
rect 8392 3612 8444 3621
rect 8484 3612 8536 3664
rect 9128 3612 9180 3664
rect 11428 3680 11480 3732
rect 11980 3680 12032 3732
rect 14832 3680 14884 3732
rect 15200 3680 15252 3732
rect 15292 3680 15344 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 18144 3723 18196 3732
rect 18144 3689 18153 3723
rect 18153 3689 18187 3723
rect 18187 3689 18196 3723
rect 18144 3680 18196 3689
rect 19064 3680 19116 3732
rect 20260 3680 20312 3732
rect 20352 3680 20404 3732
rect 20996 3680 21048 3732
rect 21456 3680 21508 3732
rect 12624 3612 12676 3664
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 13820 3612 13872 3621
rect 14004 3612 14056 3664
rect 21732 3680 21784 3732
rect 21824 3680 21876 3732
rect 22008 3680 22060 3732
rect 8024 3476 8076 3528
rect 8852 3476 8904 3528
rect 9404 3476 9456 3528
rect 11152 3544 11204 3596
rect 11244 3544 11296 3596
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 9956 3476 10008 3528
rect 10416 3476 10468 3528
rect 1400 3408 1452 3460
rect 11612 3476 11664 3528
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 15384 3544 15436 3596
rect 17408 3544 17460 3596
rect 17868 3544 17920 3596
rect 19064 3587 19116 3596
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 20168 3544 20220 3596
rect 20260 3544 20312 3596
rect 20996 3587 21048 3596
rect 20996 3553 21005 3587
rect 21005 3553 21039 3587
rect 21039 3553 21048 3587
rect 20996 3544 21048 3553
rect 21456 3587 21508 3596
rect 21456 3553 21463 3587
rect 21463 3553 21508 3587
rect 21456 3544 21508 3553
rect 17132 3476 17184 3485
rect 20904 3476 20956 3528
rect 17500 3408 17552 3460
rect 19616 3408 19668 3460
rect 20076 3408 20128 3460
rect 21916 3544 21968 3596
rect 23204 3680 23256 3732
rect 23848 3680 23900 3732
rect 26056 3680 26108 3732
rect 26700 3680 26752 3732
rect 28172 3680 28224 3732
rect 24400 3655 24452 3664
rect 24400 3621 24409 3655
rect 24409 3621 24443 3655
rect 24443 3621 24452 3655
rect 24400 3612 24452 3621
rect 24860 3612 24912 3664
rect 22928 3544 22980 3596
rect 24032 3544 24084 3596
rect 21824 3476 21876 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23296 3476 23348 3485
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 6644 3340 6696 3392
rect 8760 3340 8812 3392
rect 9036 3340 9088 3392
rect 11428 3340 11480 3392
rect 15476 3340 15528 3392
rect 16672 3340 16724 3392
rect 16856 3340 16908 3392
rect 20536 3340 20588 3392
rect 20812 3340 20864 3392
rect 23112 3383 23164 3392
rect 23112 3349 23121 3383
rect 23121 3349 23155 3383
rect 23155 3349 23164 3383
rect 23112 3340 23164 3349
rect 23664 3476 23716 3528
rect 24676 3587 24728 3596
rect 24676 3553 24685 3587
rect 24685 3553 24719 3587
rect 24719 3553 24728 3587
rect 24676 3544 24728 3553
rect 25136 3544 25188 3596
rect 25688 3544 25740 3596
rect 25872 3544 25924 3596
rect 25688 3408 25740 3460
rect 26516 3544 26568 3596
rect 27436 3587 27488 3596
rect 27436 3553 27445 3587
rect 27445 3553 27479 3587
rect 27479 3553 27488 3587
rect 27436 3544 27488 3553
rect 26792 3476 26844 3528
rect 27160 3476 27212 3528
rect 26884 3408 26936 3460
rect 23572 3340 23624 3392
rect 24492 3340 24544 3392
rect 24952 3383 25004 3392
rect 24952 3349 24961 3383
rect 24961 3349 24995 3383
rect 24995 3349 25004 3383
rect 24952 3340 25004 3349
rect 4285 3238 4337 3290
rect 4349 3238 4401 3290
rect 4413 3238 4465 3290
rect 4477 3238 4529 3290
rect 4541 3238 4593 3290
rect 12059 3238 12111 3290
rect 12123 3238 12175 3290
rect 12187 3238 12239 3290
rect 12251 3238 12303 3290
rect 12315 3238 12367 3290
rect 19833 3238 19885 3290
rect 19897 3238 19949 3290
rect 19961 3238 20013 3290
rect 20025 3238 20077 3290
rect 20089 3238 20141 3290
rect 27607 3238 27659 3290
rect 27671 3238 27723 3290
rect 27735 3238 27787 3290
rect 27799 3238 27851 3290
rect 27863 3238 27915 3290
rect 1676 3136 1728 3188
rect 2320 3136 2372 3188
rect 3240 3136 3292 3188
rect 3700 3136 3752 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6828 3136 6880 3188
rect 7840 3136 7892 3188
rect 8392 3136 8444 3188
rect 8576 3136 8628 3188
rect 2780 3000 2832 3052
rect 2872 3000 2924 3052
rect 3792 3000 3844 3052
rect 6736 3000 6788 3052
rect 2504 2864 2556 2916
rect 7104 2932 7156 2984
rect 7748 3000 7800 3052
rect 8484 3000 8536 3052
rect 7932 2932 7984 2984
rect 8852 3068 8904 3120
rect 11152 3136 11204 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 15384 3136 15436 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 11428 3068 11480 3120
rect 11796 3068 11848 3120
rect 9036 2932 9088 2984
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 10416 2864 10468 2916
rect 11520 3000 11572 3052
rect 13912 3000 13964 3052
rect 15292 3000 15344 3052
rect 15568 3000 15620 3052
rect 16856 3136 16908 3188
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 18604 3136 18656 3188
rect 11980 2932 12032 2984
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 16764 2932 16816 2984
rect 20444 3179 20496 3188
rect 20444 3145 20453 3179
rect 20453 3145 20487 3179
rect 20487 3145 20496 3179
rect 20444 3136 20496 3145
rect 20536 3136 20588 3188
rect 22100 3136 22152 3188
rect 23020 3136 23072 3188
rect 23112 3136 23164 3188
rect 23296 3179 23348 3188
rect 23296 3145 23305 3179
rect 23305 3145 23339 3179
rect 23339 3145 23348 3179
rect 23296 3136 23348 3145
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 10324 2796 10376 2848
rect 13544 2864 13596 2916
rect 16396 2864 16448 2916
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 17408 2932 17460 2984
rect 19616 3000 19668 3052
rect 19708 3000 19760 3052
rect 20720 3068 20772 3120
rect 21824 3068 21876 3120
rect 10784 2796 10836 2848
rect 16580 2796 16632 2848
rect 17592 2864 17644 2916
rect 19800 2932 19852 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 20260 2932 20312 2984
rect 21732 3000 21784 3052
rect 21548 2932 21600 2984
rect 18420 2864 18472 2916
rect 18696 2907 18748 2916
rect 18696 2873 18705 2907
rect 18705 2873 18739 2907
rect 18739 2873 18748 2907
rect 18696 2864 18748 2873
rect 21272 2864 21324 2916
rect 17684 2839 17736 2848
rect 17684 2805 17693 2839
rect 17693 2805 17727 2839
rect 17727 2805 17736 2839
rect 17684 2796 17736 2805
rect 18880 2839 18932 2848
rect 18880 2805 18905 2839
rect 18905 2805 18932 2839
rect 18880 2796 18932 2805
rect 19064 2839 19116 2848
rect 19064 2805 19073 2839
rect 19073 2805 19107 2839
rect 19107 2805 19116 2839
rect 19064 2796 19116 2805
rect 19340 2796 19392 2848
rect 19984 2796 20036 2848
rect 20076 2796 20128 2848
rect 22100 2864 22152 2916
rect 22376 2907 22428 2916
rect 22376 2873 22385 2907
rect 22385 2873 22419 2907
rect 22419 2873 22428 2907
rect 22376 2864 22428 2873
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 23204 2975 23256 2984
rect 23204 2941 23213 2975
rect 23213 2941 23247 2975
rect 23247 2941 23256 2975
rect 23204 2932 23256 2941
rect 23388 2932 23440 2984
rect 24124 3136 24176 3188
rect 24860 3136 24912 3188
rect 24952 3136 25004 3188
rect 23756 3068 23808 3120
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 24216 3000 24268 3052
rect 24676 3000 24728 3052
rect 23940 2864 23992 2916
rect 24216 2864 24268 2916
rect 24124 2839 24176 2848
rect 24124 2805 24133 2839
rect 24133 2805 24167 2839
rect 24167 2805 24176 2839
rect 24124 2796 24176 2805
rect 24952 2932 25004 2984
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 27160 3179 27212 3188
rect 27160 3145 27169 3179
rect 27169 3145 27203 3179
rect 27203 3145 27212 3179
rect 27160 3136 27212 3145
rect 26976 3068 27028 3120
rect 24676 2907 24728 2916
rect 24676 2873 24685 2907
rect 24685 2873 24719 2907
rect 24719 2873 24728 2907
rect 24676 2864 24728 2873
rect 25044 2864 25096 2916
rect 25320 2864 25372 2916
rect 25596 2932 25648 2984
rect 27436 3000 27488 3052
rect 26424 2839 26476 2848
rect 26424 2805 26433 2839
rect 26433 2805 26467 2839
rect 26467 2805 26476 2839
rect 26424 2796 26476 2805
rect 27344 2839 27396 2848
rect 27344 2805 27353 2839
rect 27353 2805 27387 2839
rect 27387 2805 27396 2839
rect 27344 2796 27396 2805
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 15946 2694 15998 2746
rect 16010 2694 16062 2746
rect 16074 2694 16126 2746
rect 16138 2694 16190 2746
rect 16202 2694 16254 2746
rect 23720 2694 23772 2746
rect 23784 2694 23836 2746
rect 23848 2694 23900 2746
rect 23912 2694 23964 2746
rect 23976 2694 24028 2746
rect 31494 2694 31546 2746
rect 31558 2694 31610 2746
rect 31622 2694 31674 2746
rect 31686 2694 31738 2746
rect 31750 2694 31802 2746
rect 7472 2592 7524 2644
rect 9220 2592 9272 2644
rect 15660 2592 15712 2644
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 17592 2592 17644 2644
rect 17684 2592 17736 2644
rect 13544 2567 13596 2576
rect 13544 2533 13553 2567
rect 13553 2533 13587 2567
rect 13587 2533 13596 2567
rect 13544 2524 13596 2533
rect 15844 2524 15896 2576
rect 18236 2635 18288 2644
rect 18236 2601 18245 2635
rect 18245 2601 18279 2635
rect 18279 2601 18288 2635
rect 18236 2592 18288 2601
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 18880 2592 18932 2644
rect 21364 2635 21416 2644
rect 8668 2456 8720 2508
rect 9680 2456 9732 2508
rect 14004 2499 14056 2508
rect 14004 2465 14013 2499
rect 14013 2465 14047 2499
rect 14047 2465 14056 2499
rect 14004 2456 14056 2465
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 15200 2499 15252 2508
rect 15200 2465 15209 2499
rect 15209 2465 15243 2499
rect 15243 2465 15252 2499
rect 15200 2456 15252 2465
rect 15384 2499 15436 2508
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 17684 2456 17736 2508
rect 15752 2388 15804 2440
rect 16580 2388 16632 2440
rect 17960 2456 18012 2508
rect 18512 2456 18564 2508
rect 18604 2499 18656 2508
rect 18604 2465 18613 2499
rect 18613 2465 18647 2499
rect 18647 2465 18656 2499
rect 18604 2456 18656 2465
rect 18144 2320 18196 2372
rect 19064 2499 19116 2508
rect 19064 2465 19073 2499
rect 19073 2465 19107 2499
rect 19107 2465 19116 2499
rect 19064 2456 19116 2465
rect 19248 2456 19300 2508
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 18788 2388 18840 2440
rect 18972 2388 19024 2440
rect 20904 2524 20956 2576
rect 21916 2592 21968 2644
rect 22376 2592 22428 2644
rect 23388 2592 23440 2644
rect 19616 2456 19668 2508
rect 19984 2456 20036 2508
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 20996 2499 21048 2508
rect 20996 2465 21005 2499
rect 21005 2465 21039 2499
rect 21039 2465 21048 2499
rect 20996 2456 21048 2465
rect 21548 2567 21600 2576
rect 21548 2533 21557 2567
rect 21557 2533 21591 2567
rect 21591 2533 21600 2567
rect 21548 2524 21600 2533
rect 21272 2499 21324 2508
rect 21272 2465 21281 2499
rect 21281 2465 21315 2499
rect 21315 2465 21324 2499
rect 21272 2456 21324 2465
rect 20352 2388 20404 2440
rect 21456 2388 21508 2440
rect 19800 2320 19852 2372
rect 22008 2499 22060 2508
rect 22008 2465 22017 2499
rect 22017 2465 22051 2499
rect 22051 2465 22060 2499
rect 22008 2456 22060 2465
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 22192 2456 22244 2465
rect 23572 2499 23624 2508
rect 23572 2465 23581 2499
rect 23581 2465 23615 2499
rect 23615 2465 23624 2499
rect 23572 2456 23624 2465
rect 25412 2592 25464 2644
rect 24768 2524 24820 2576
rect 24952 2524 25004 2576
rect 18972 2252 19024 2304
rect 22100 2320 22152 2372
rect 21824 2252 21876 2304
rect 22284 2252 22336 2304
rect 24032 2388 24084 2440
rect 24308 2456 24360 2508
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 25228 2456 25280 2508
rect 25504 2499 25556 2508
rect 25504 2465 25513 2499
rect 25513 2465 25547 2499
rect 25547 2465 25556 2499
rect 25504 2456 25556 2465
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 26608 2592 26660 2644
rect 26424 2499 26476 2508
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 24768 2388 24820 2440
rect 25596 2388 25648 2440
rect 26148 2388 26200 2440
rect 23480 2320 23532 2372
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 24216 2320 24268 2372
rect 26516 2363 26568 2372
rect 26516 2329 26525 2363
rect 26525 2329 26559 2363
rect 26559 2329 26568 2363
rect 26516 2320 26568 2329
rect 27344 2320 27396 2372
rect 24308 2252 24360 2304
rect 24676 2252 24728 2304
rect 4285 2150 4337 2202
rect 4349 2150 4401 2202
rect 4413 2150 4465 2202
rect 4477 2150 4529 2202
rect 4541 2150 4593 2202
rect 12059 2150 12111 2202
rect 12123 2150 12175 2202
rect 12187 2150 12239 2202
rect 12251 2150 12303 2202
rect 12315 2150 12367 2202
rect 19833 2150 19885 2202
rect 19897 2150 19949 2202
rect 19961 2150 20013 2202
rect 20025 2150 20077 2202
rect 20089 2150 20141 2202
rect 27607 2150 27659 2202
rect 27671 2150 27723 2202
rect 27735 2150 27787 2202
rect 27799 2150 27851 2202
rect 27863 2150 27915 2202
rect 15292 2048 15344 2100
rect 15844 2048 15896 2100
rect 17132 2048 17184 2100
rect 17500 1980 17552 2032
rect 18144 2091 18196 2100
rect 18144 2057 18153 2091
rect 18153 2057 18187 2091
rect 18187 2057 18196 2091
rect 18144 2048 18196 2057
rect 18880 2091 18932 2100
rect 18880 2057 18889 2091
rect 18889 2057 18923 2091
rect 18923 2057 18932 2091
rect 18880 2048 18932 2057
rect 19340 2091 19392 2100
rect 19340 2057 19349 2091
rect 19349 2057 19383 2091
rect 19383 2057 19392 2091
rect 19340 2048 19392 2057
rect 19616 1980 19668 2032
rect 16580 1844 16632 1896
rect 19064 1912 19116 1964
rect 19708 1887 19760 1896
rect 19708 1853 19717 1887
rect 19717 1853 19751 1887
rect 19751 1853 19760 1887
rect 20352 1887 20404 1896
rect 19708 1844 19760 1853
rect 20352 1853 20361 1887
rect 20361 1853 20395 1887
rect 20395 1853 20404 1887
rect 20352 1844 20404 1853
rect 20904 2048 20956 2100
rect 21272 2048 21324 2100
rect 22284 2091 22336 2100
rect 22284 2057 22293 2091
rect 22293 2057 22327 2091
rect 22327 2057 22336 2091
rect 22284 2048 22336 2057
rect 23756 2048 23808 2100
rect 24400 2091 24452 2100
rect 24400 2057 24409 2091
rect 24409 2057 24443 2091
rect 24443 2057 24452 2091
rect 24400 2048 24452 2057
rect 20812 1887 20864 1896
rect 20812 1853 20821 1887
rect 20821 1853 20855 1887
rect 20855 1853 20864 1887
rect 20812 1844 20864 1853
rect 23480 1980 23532 2032
rect 21916 1955 21968 1964
rect 21916 1921 21925 1955
rect 21925 1921 21959 1955
rect 21959 1921 21968 1955
rect 24584 2048 24636 2100
rect 25320 2048 25372 2100
rect 25504 2048 25556 2100
rect 21916 1912 21968 1921
rect 20444 1776 20496 1828
rect 21548 1844 21600 1896
rect 21732 1776 21784 1828
rect 24860 1955 24912 1964
rect 24860 1921 24869 1955
rect 24869 1921 24903 1955
rect 24903 1921 24912 1955
rect 24860 1912 24912 1921
rect 24768 1853 24777 1886
rect 24777 1853 24811 1886
rect 24811 1853 24820 1886
rect 24768 1834 24820 1853
rect 25688 1980 25740 2032
rect 25964 2048 26016 2100
rect 26608 2091 26660 2100
rect 26608 2057 26617 2091
rect 26617 2057 26651 2091
rect 26651 2057 26660 2091
rect 26608 2048 26660 2057
rect 26148 1980 26200 2032
rect 26240 1912 26292 1964
rect 27988 1912 28040 1964
rect 24860 1776 24912 1828
rect 26516 1776 26568 1828
rect 15752 1708 15804 1760
rect 18972 1708 19024 1760
rect 19156 1708 19208 1760
rect 20812 1708 20864 1760
rect 8172 1606 8224 1658
rect 8236 1606 8288 1658
rect 8300 1606 8352 1658
rect 8364 1606 8416 1658
rect 8428 1606 8480 1658
rect 15946 1606 15998 1658
rect 16010 1606 16062 1658
rect 16074 1606 16126 1658
rect 16138 1606 16190 1658
rect 16202 1606 16254 1658
rect 23720 1606 23772 1658
rect 23784 1606 23836 1658
rect 23848 1606 23900 1658
rect 23912 1606 23964 1658
rect 23976 1606 24028 1658
rect 31494 1606 31546 1658
rect 31558 1606 31610 1658
rect 31622 1606 31674 1658
rect 31686 1606 31738 1658
rect 31750 1606 31802 1658
rect 19248 1504 19300 1556
rect 19340 1504 19392 1556
rect 14188 1436 14240 1488
rect 19156 1368 19208 1420
rect 19064 1343 19116 1352
rect 19064 1309 19073 1343
rect 19073 1309 19107 1343
rect 19107 1309 19116 1343
rect 19064 1300 19116 1309
rect 20444 1504 20496 1556
rect 21364 1504 21416 1556
rect 26240 1504 26292 1556
rect 21824 1436 21876 1488
rect 19708 1411 19760 1420
rect 19708 1377 19717 1411
rect 19717 1377 19751 1411
rect 19751 1377 19760 1411
rect 19708 1368 19760 1377
rect 4285 1062 4337 1114
rect 4349 1062 4401 1114
rect 4413 1062 4465 1114
rect 4477 1062 4529 1114
rect 4541 1062 4593 1114
rect 12059 1062 12111 1114
rect 12123 1062 12175 1114
rect 12187 1062 12239 1114
rect 12251 1062 12303 1114
rect 12315 1062 12367 1114
rect 19833 1062 19885 1114
rect 19897 1062 19949 1114
rect 19961 1062 20013 1114
rect 20025 1062 20077 1114
rect 20089 1062 20141 1114
rect 27607 1062 27659 1114
rect 27671 1062 27723 1114
rect 27735 1062 27787 1114
rect 27799 1062 27851 1114
rect 27863 1062 27915 1114
rect 8172 518 8224 570
rect 8236 518 8288 570
rect 8300 518 8352 570
rect 8364 518 8416 570
rect 8428 518 8480 570
rect 15946 518 15998 570
rect 16010 518 16062 570
rect 16074 518 16126 570
rect 16138 518 16190 570
rect 16202 518 16254 570
rect 23720 518 23772 570
rect 23784 518 23836 570
rect 23848 518 23900 570
rect 23912 518 23964 570
rect 23976 518 24028 570
rect 31494 518 31546 570
rect 31558 518 31610 570
rect 31622 518 31674 570
rect 31686 518 31738 570
rect 31750 518 31802 570
<< metal2 >>
rect 13726 22128 13782 22137
rect 13648 22086 13726 22114
rect 5080 22024 5132 22030
rect 4526 21992 4582 22001
rect 4068 21956 4120 21962
rect 4582 21950 4752 21978
rect 5080 21966 5132 21972
rect 12530 21992 12586 22001
rect 4526 21927 4582 21936
rect 4068 21898 4120 21904
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 1308 21548 1360 21554
rect 1308 21490 1360 21496
rect 1320 21321 1348 21490
rect 3528 21486 3556 21830
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 1306 21312 1362 21321
rect 1306 21247 1362 21256
rect 2134 21176 2190 21185
rect 2134 21111 2136 21120
rect 2188 21111 2190 21120
rect 2136 21082 2188 21088
rect 1216 20936 1268 20942
rect 1216 20878 1268 20884
rect 940 20800 992 20806
rect 940 20742 992 20748
rect 952 19718 980 20742
rect 1124 20256 1176 20262
rect 1124 20198 1176 20204
rect 1136 20058 1164 20198
rect 1124 20052 1176 20058
rect 1124 19994 1176 20000
rect 940 19712 992 19718
rect 940 19654 992 19660
rect 952 19514 980 19654
rect 940 19508 992 19514
rect 940 19450 992 19456
rect 952 19334 980 19450
rect 952 19306 1072 19334
rect 1044 18290 1072 19306
rect 1124 19236 1176 19242
rect 1124 19178 1176 19184
rect 1136 18970 1164 19178
rect 1124 18964 1176 18970
rect 1124 18906 1176 18912
rect 1228 18630 1256 20878
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1596 20398 1624 20703
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 2056 18970 2084 20198
rect 2148 18970 2176 21082
rect 2240 21010 2268 21354
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 2240 19922 2268 20946
rect 2700 20602 2728 21422
rect 3608 21412 3660 21418
rect 3608 21354 3660 21360
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 2964 21344 3016 21350
rect 2884 21292 2964 21298
rect 2884 21286 3016 21292
rect 2884 21270 3004 21286
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2516 18873 2544 20402
rect 2884 20398 2912 21270
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3330 20768 3386 20777
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2608 19174 2636 20198
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2700 19718 2728 19858
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 18902 2636 19110
rect 2596 18896 2648 18902
rect 2502 18864 2558 18873
rect 2596 18838 2648 18844
rect 2502 18799 2558 18808
rect 2516 18766 2544 18799
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 1216 18624 1268 18630
rect 1216 18566 1268 18572
rect 2608 18426 2636 18702
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 1032 18284 1084 18290
rect 1032 18226 1084 18232
rect 2700 18154 2728 19246
rect 2792 18970 2820 20266
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2884 18698 2912 20334
rect 3252 20330 3280 20742
rect 3330 20703 3386 20712
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 3344 19990 3372 20703
rect 3620 20466 3648 21354
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3804 20942 3832 21286
rect 3896 21146 3924 21354
rect 3974 21176 4030 21185
rect 3884 21140 3936 21146
rect 4080 21146 4108 21898
rect 4285 21788 4593 21797
rect 4285 21786 4291 21788
rect 4347 21786 4371 21788
rect 4427 21786 4451 21788
rect 4507 21786 4531 21788
rect 4587 21786 4593 21788
rect 4347 21734 4349 21786
rect 4529 21734 4531 21786
rect 4285 21732 4291 21734
rect 4347 21732 4371 21734
rect 4427 21732 4451 21734
rect 4507 21732 4531 21734
rect 4587 21732 4593 21734
rect 4285 21723 4593 21732
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 3974 21111 3976 21120
rect 3884 21082 3936 21088
rect 4028 21111 4030 21120
rect 4068 21140 4120 21146
rect 3976 21082 4028 21088
rect 4068 21082 4120 21088
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3988 20754 4016 21082
rect 3988 20726 4200 20754
rect 4172 20466 4200 20726
rect 4285 20700 4593 20709
rect 4285 20698 4291 20700
rect 4347 20698 4371 20700
rect 4427 20698 4451 20700
rect 4507 20698 4531 20700
rect 4587 20698 4593 20700
rect 4347 20646 4349 20698
rect 4529 20646 4531 20698
rect 4285 20644 4291 20646
rect 4347 20644 4371 20646
rect 4427 20644 4451 20646
rect 4507 20644 4531 20646
rect 4587 20644 4593 20646
rect 4285 20635 4593 20644
rect 4632 20602 4660 21286
rect 4724 21078 4752 21950
rect 4988 21616 5040 21622
rect 4986 21584 4988 21593
rect 5040 21584 5042 21593
rect 4986 21519 5042 21528
rect 5000 21146 5028 21519
rect 5092 21146 5120 21966
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10324 21956 10376 21962
rect 12530 21927 12586 21936
rect 10324 21898 10376 21904
rect 7010 21856 7066 21865
rect 7010 21791 7066 21800
rect 8850 21856 8906 21865
rect 8850 21791 8906 21800
rect 7024 21690 7052 21791
rect 8864 21690 8892 21791
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 6276 21548 6328 21554
rect 6276 21490 6328 21496
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3620 19922 3648 20402
rect 4540 20262 4568 20470
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 19514 3096 19790
rect 3620 19786 3648 19858
rect 3608 19780 3660 19786
rect 3608 19722 3660 19728
rect 3988 19718 4016 19994
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3252 18970 3280 19178
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3068 18426 3096 18566
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2700 18057 2728 18090
rect 2686 18048 2742 18057
rect 2608 18006 2686 18034
rect 2608 17814 2636 18006
rect 2686 17983 2742 17992
rect 2792 17882 2820 18362
rect 3252 18358 3280 18906
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3344 18154 3372 19110
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 1124 17672 1176 17678
rect 1124 17614 1176 17620
rect 1136 17338 1164 17614
rect 1124 17332 1176 17338
rect 1124 17274 1176 17280
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 1124 16584 1176 16590
rect 1124 16526 1176 16532
rect 1136 16250 1164 16526
rect 1124 16244 1176 16250
rect 1124 16186 1176 16192
rect 1032 16176 1084 16182
rect 1032 16118 1084 16124
rect 1044 15706 1072 16118
rect 2148 16114 2176 17138
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1032 15700 1084 15706
rect 1032 15642 1084 15648
rect 940 15360 992 15366
rect 940 15302 992 15308
rect 756 15020 808 15026
rect 756 14962 808 14968
rect 768 5846 796 14962
rect 952 14958 980 15302
rect 940 14952 992 14958
rect 940 14894 992 14900
rect 1216 14952 1268 14958
rect 1216 14894 1268 14900
rect 952 13870 980 14894
rect 1228 14618 1256 14894
rect 2148 14618 2176 16050
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 1216 14612 1268 14618
rect 1216 14554 1268 14560
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 1216 13864 1268 13870
rect 1216 13806 1268 13812
rect 952 13258 980 13806
rect 1228 13530 1256 13806
rect 1216 13524 1268 13530
rect 1216 13466 1268 13472
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 952 12850 980 13194
rect 940 12844 992 12850
rect 940 12786 992 12792
rect 1308 12708 1360 12714
rect 1308 12650 1360 12656
rect 1320 12442 1348 12650
rect 1308 12436 1360 12442
rect 1780 12434 1808 14418
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 13394 2176 14350
rect 2240 13802 2268 14826
rect 2228 13796 2280 13802
rect 2280 13756 2360 13784
rect 2228 13738 2280 13744
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2332 12782 2360 13756
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 1780 12406 1900 12434
rect 1308 12378 1360 12384
rect 848 11688 900 11694
rect 848 11630 900 11636
rect 860 10674 888 11630
rect 1124 11620 1176 11626
rect 1124 11562 1176 11568
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 1136 11354 1164 11562
rect 1124 11348 1176 11354
rect 1124 11290 1176 11296
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 1780 10538 1808 11562
rect 1768 10532 1820 10538
rect 1768 10474 1820 10480
rect 1780 9926 1808 10474
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9450 1808 9862
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 860 7342 888 8366
rect 1216 8356 1268 8362
rect 1216 8298 1268 8304
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 1030 7440 1086 7449
rect 1030 7375 1086 7384
rect 848 7336 900 7342
rect 848 7278 900 7284
rect 860 6322 888 7278
rect 940 7200 992 7206
rect 940 7142 992 7148
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 756 5840 808 5846
rect 756 5782 808 5788
rect 860 5234 888 6258
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 952 4554 980 7142
rect 1044 6866 1072 7375
rect 1032 6860 1084 6866
rect 1032 6802 1084 6808
rect 1032 6656 1084 6662
rect 1032 6598 1084 6604
rect 1044 4826 1072 6598
rect 1136 5642 1164 7890
rect 1228 7410 1256 8298
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1596 7954 1624 8026
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1216 7404 1268 7410
rect 1216 7346 1268 7352
rect 1504 6866 1532 7890
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7002 1716 7754
rect 1780 7750 1808 7958
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1766 6896 1822 6905
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1584 6860 1636 6866
rect 1766 6831 1822 6840
rect 1584 6802 1636 6808
rect 1412 6458 1440 6802
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1216 6248 1268 6254
rect 1216 6190 1268 6196
rect 1124 5636 1176 5642
rect 1124 5578 1176 5584
rect 1124 5092 1176 5098
rect 1124 5034 1176 5040
rect 1032 4820 1084 4826
rect 1032 4762 1084 4768
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 1032 4548 1084 4554
rect 1032 4490 1084 4496
rect 1044 4146 1072 4490
rect 1136 4282 1164 5034
rect 1228 4826 1256 6190
rect 1492 5908 1544 5914
rect 1596 5896 1624 6802
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1544 5868 1624 5896
rect 1492 5850 1544 5856
rect 1688 4826 1716 6666
rect 1780 5778 1808 6831
rect 1872 5846 1900 12406
rect 2516 12238 2544 16934
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 16046 2636 16390
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2700 15502 2728 17682
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2976 17338 3004 17614
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2884 17134 2912 17206
rect 2872 17128 2924 17134
rect 3068 17082 3096 17478
rect 3436 17338 3464 18770
rect 3528 18426 3556 18770
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3620 18290 3648 19110
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3712 17542 3740 18838
rect 3790 18184 3846 18193
rect 3790 18119 3792 18128
rect 3844 18119 3846 18128
rect 3792 18090 3844 18096
rect 3804 17882 3832 18090
rect 3988 18057 4016 19654
rect 4172 19394 4200 20198
rect 5000 19990 5028 20266
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 4285 19612 4593 19621
rect 4285 19610 4291 19612
rect 4347 19610 4371 19612
rect 4427 19610 4451 19612
rect 4507 19610 4531 19612
rect 4587 19610 4593 19612
rect 4347 19558 4349 19610
rect 4529 19558 4531 19610
rect 4285 19556 4291 19558
rect 4347 19556 4371 19558
rect 4427 19556 4451 19558
rect 4507 19556 4531 19558
rect 4587 19556 4593 19558
rect 4285 19547 4593 19556
rect 4250 19408 4306 19417
rect 4172 19366 4250 19394
rect 4250 19343 4306 19352
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18970 4108 19110
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4356 18873 4384 19314
rect 4342 18864 4398 18873
rect 4342 18799 4398 18808
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4250 18728 4306 18737
rect 4080 18154 4108 18702
rect 4250 18663 4252 18672
rect 4304 18663 4306 18672
rect 4252 18634 4304 18640
rect 4285 18524 4593 18533
rect 4285 18522 4291 18524
rect 4347 18522 4371 18524
rect 4427 18522 4451 18524
rect 4507 18522 4531 18524
rect 4587 18522 4593 18524
rect 4347 18470 4349 18522
rect 4529 18470 4531 18522
rect 4285 18468 4291 18470
rect 4347 18468 4371 18470
rect 4427 18468 4451 18470
rect 4507 18468 4531 18470
rect 4587 18468 4593 18470
rect 4285 18459 4593 18468
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3974 18048 4030 18057
rect 3974 17983 4030 17992
rect 3988 17882 4016 17983
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2872 17070 2924 17076
rect 2884 16946 2912 17070
rect 2976 17066 3096 17082
rect 2964 17060 3096 17066
rect 3016 17054 3096 17060
rect 2964 17002 3016 17008
rect 3516 16992 3568 16998
rect 2884 16918 3096 16946
rect 3516 16934 3568 16940
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 15638 2820 16594
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14482 2636 14758
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2700 13326 2728 14962
rect 2792 14890 2820 15574
rect 2884 15366 2912 15982
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2792 14074 2820 14350
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2792 13462 2820 13670
rect 2884 13530 2912 13806
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12238 2728 13262
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2792 12442 2820 12854
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2136 12096 2188 12102
rect 2056 12044 2136 12050
rect 2056 12038 2188 12044
rect 2056 12022 2176 12038
rect 2056 11218 2084 12022
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2056 9178 2084 11154
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2148 10130 2176 10678
rect 2332 10674 2360 11086
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 10198 2360 10610
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2148 9518 2176 10066
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2148 9042 2176 9454
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8129 2084 8774
rect 2042 8120 2098 8129
rect 2042 8055 2098 8064
rect 1952 7880 2004 7886
rect 2004 7840 2084 7868
rect 1952 7822 2004 7828
rect 1950 6760 2006 6769
rect 1950 6695 2006 6704
rect 1964 5914 1992 6695
rect 2056 6254 2084 7840
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 2056 5710 2084 6190
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 2148 4758 2176 8978
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7342 2268 7822
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 6186 2268 7278
rect 2332 6798 2360 10134
rect 2516 9654 2544 12174
rect 2976 11898 3004 13330
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11218 2636 11494
rect 2884 11354 2912 11630
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2608 10266 2636 10746
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10266 2820 10406
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2424 8634 2452 8910
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2516 8566 2544 9590
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2516 6934 2544 8502
rect 2608 7206 2636 9114
rect 2792 7478 2820 9998
rect 2976 8362 3004 11562
rect 3068 8362 3096 16918
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3160 15094 3188 16050
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3160 8838 3188 12786
rect 3252 10554 3280 15846
rect 3344 15570 3372 15846
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3436 15162 3464 16526
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3528 15026 3556 16934
rect 3620 16046 3648 16934
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3620 14958 3648 15982
rect 3712 15162 3740 16730
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3804 16454 3832 16526
rect 3896 16454 3924 16934
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3608 14952 3660 14958
rect 3344 14900 3608 14906
rect 3804 14906 3832 15438
rect 3344 14894 3660 14900
rect 3344 14878 3648 14894
rect 3712 14878 3832 14906
rect 3344 12102 3372 14878
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 14074 3556 14214
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3436 13530 3464 14010
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3436 12782 3464 13466
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3528 12434 3556 14010
rect 3620 12782 3648 14758
rect 3712 13326 3740 14878
rect 3896 14362 3924 16390
rect 3988 14618 4016 17614
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4080 16182 4108 17138
rect 4172 17134 4200 18294
rect 4434 18184 4490 18193
rect 4632 18170 4660 19314
rect 5368 19310 5396 19654
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5460 19242 5488 20946
rect 5552 19922 5580 21490
rect 6184 21344 6236 21350
rect 6182 21312 6184 21321
rect 6236 21312 6238 21321
rect 6182 21247 6238 21256
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 19990 5672 20742
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 4816 18970 4844 19110
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4724 18850 4752 18906
rect 4724 18822 4844 18850
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4434 18119 4436 18128
rect 4488 18119 4490 18128
rect 4540 18142 4660 18170
rect 4436 18090 4488 18096
rect 4448 17746 4476 18090
rect 4540 17814 4568 18142
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4528 17808 4580 17814
rect 4528 17750 4580 17756
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4285 17436 4593 17445
rect 4285 17434 4291 17436
rect 4347 17434 4371 17436
rect 4427 17434 4451 17436
rect 4507 17434 4531 17436
rect 4587 17434 4593 17436
rect 4347 17382 4349 17434
rect 4529 17382 4531 17434
rect 4285 17380 4291 17382
rect 4347 17380 4371 17382
rect 4427 17380 4451 17382
rect 4507 17380 4531 17382
rect 4587 17380 4593 17382
rect 4285 17371 4593 17380
rect 4160 17128 4212 17134
rect 4632 17082 4660 18022
rect 4724 17542 4752 18702
rect 4816 18698 4844 18822
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4908 18426 4936 19110
rect 5276 18970 5304 19110
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5080 18828 5132 18834
rect 5132 18788 5304 18816
rect 5080 18770 5132 18776
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18426 5028 18566
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4988 18284 5040 18290
rect 5040 18244 5120 18272
rect 4988 18226 5040 18232
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 17270 4752 17478
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4160 17070 4212 17076
rect 4540 17066 4660 17082
rect 4528 17060 4660 17066
rect 4580 17054 4660 17060
rect 4528 17002 4580 17008
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4080 15502 4108 16118
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3804 14334 3924 14362
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3528 12406 3648 12434
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3620 11898 3648 12406
rect 3804 12306 3832 14334
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 12714 3924 13670
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3896 12442 3924 12650
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3988 12374 4016 12650
rect 4080 12374 4108 14758
rect 4172 14414 4200 16934
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4285 16348 4593 16357
rect 4285 16346 4291 16348
rect 4347 16346 4371 16348
rect 4427 16346 4451 16348
rect 4507 16346 4531 16348
rect 4587 16346 4593 16348
rect 4347 16294 4349 16346
rect 4529 16294 4531 16346
rect 4285 16292 4291 16294
rect 4347 16292 4371 16294
rect 4427 16292 4451 16294
rect 4507 16292 4531 16294
rect 4587 16292 4593 16294
rect 4285 16283 4593 16292
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4285 15260 4593 15269
rect 4285 15258 4291 15260
rect 4347 15258 4371 15260
rect 4427 15258 4451 15260
rect 4507 15258 4531 15260
rect 4587 15258 4593 15260
rect 4347 15206 4349 15258
rect 4529 15206 4531 15258
rect 4285 15204 4291 15206
rect 4347 15204 4371 15206
rect 4427 15204 4451 15206
rect 4507 15204 4531 15206
rect 4587 15204 4593 15206
rect 4285 15195 4593 15204
rect 4632 14822 4660 15846
rect 4724 15722 4752 16594
rect 4816 16454 4844 18022
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4724 15694 4844 15722
rect 4816 15570 4844 15694
rect 4804 15564 4856 15570
rect 4724 15524 4804 15552
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4264 14260 4292 14758
rect 4724 14618 4752 15524
rect 4804 15506 4856 15512
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14618 4844 14826
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4172 14232 4292 14260
rect 4528 14272 4580 14278
rect 4172 14074 4200 14232
rect 4580 14232 4660 14260
rect 4528 14214 4580 14220
rect 4285 14172 4593 14181
rect 4285 14170 4291 14172
rect 4347 14170 4371 14172
rect 4427 14170 4451 14172
rect 4507 14170 4531 14172
rect 4587 14170 4593 14172
rect 4347 14118 4349 14170
rect 4529 14118 4531 14170
rect 4285 14116 4291 14118
rect 4347 14116 4371 14118
rect 4427 14116 4451 14118
rect 4507 14116 4531 14118
rect 4587 14116 4593 14118
rect 4285 14107 4593 14116
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12986 4200 13262
rect 4285 13084 4593 13093
rect 4285 13082 4291 13084
rect 4347 13082 4371 13084
rect 4427 13082 4451 13084
rect 4507 13082 4531 13084
rect 4587 13082 4593 13084
rect 4347 13030 4349 13082
rect 4529 13030 4531 13082
rect 4285 13028 4291 13030
rect 4347 13028 4371 13030
rect 4427 13028 4451 13030
rect 4507 13028 4531 13030
rect 4587 13028 4593 13030
rect 4285 13019 4593 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4632 12850 4660 14232
rect 4724 13734 4752 14554
rect 4908 14498 4936 17478
rect 5092 17241 5120 18244
rect 5276 18086 5304 18788
rect 5368 18222 5396 19110
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5460 18426 5488 18702
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 18329 5488 18362
rect 5446 18320 5502 18329
rect 5446 18255 5502 18264
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5078 17232 5134 17241
rect 5078 17167 5134 17176
rect 5092 17134 5120 17167
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5184 16794 5212 17070
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5276 16522 5304 18022
rect 5460 17762 5488 18255
rect 5368 17734 5488 17762
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5184 16114 5212 16390
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5000 15366 5028 16050
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4816 14470 4936 14498
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13462 4752 13670
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4816 13308 4844 14470
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 14074 4936 14350
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4724 13280 4844 13308
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3436 11150 3464 11834
rect 3988 11778 4016 12310
rect 3516 11756 3568 11762
rect 3988 11750 4108 11778
rect 3516 11698 3568 11704
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3252 10538 3372 10554
rect 3252 10532 3384 10538
rect 3252 10526 3332 10532
rect 3332 10474 3384 10480
rect 3238 8936 3294 8945
rect 3238 8871 3294 8880
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3160 8294 3188 8774
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 2870 8120 2926 8129
rect 2870 8055 2926 8064
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2884 7342 2912 8055
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2228 6180 2280 6186
rect 2280 6140 2360 6168
rect 2228 6122 2280 6128
rect 2332 5234 2360 6140
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 1124 4276 1176 4282
rect 1124 4218 1176 4224
rect 1032 4140 1084 4146
rect 1032 4082 1084 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1400 4004 1452 4010
rect 1400 3946 1452 3952
rect 1412 3466 1440 3946
rect 2056 3738 2084 4082
rect 2332 4060 2360 5170
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2424 5030 2452 5102
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2424 4690 2452 4966
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2412 4072 2464 4078
rect 2332 4032 2412 4060
rect 2412 4014 2464 4020
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1688 3194 1716 3538
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2332 3194 2360 3470
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2516 2922 2544 6870
rect 2608 4826 2636 7142
rect 2792 6866 2820 7210
rect 2976 7188 3004 7414
rect 2884 7160 3004 7188
rect 2884 6866 2912 7160
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6118 2912 6802
rect 3160 6798 3188 8230
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2976 6458 3004 6734
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5556 2728 5714
rect 2792 5710 2820 6054
rect 2976 5930 3004 6394
rect 2884 5914 3004 5930
rect 2872 5908 3004 5914
rect 2924 5902 3004 5908
rect 2872 5850 2924 5856
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2700 5528 2912 5556
rect 2884 5302 2912 5528
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4826 2912 4966
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2608 4060 2636 4422
rect 2700 4162 2728 4694
rect 2780 4208 2832 4214
rect 2700 4156 2780 4162
rect 2700 4150 2832 4156
rect 2700 4134 2820 4150
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 4072 2832 4078
rect 2608 4032 2780 4060
rect 2780 4014 2832 4020
rect 2792 3058 2820 4014
rect 2884 3058 2912 4082
rect 3068 4078 3096 6734
rect 3252 4146 3280 8871
rect 3344 5030 3372 10474
rect 3436 10062 3464 11086
rect 3528 10742 3556 11698
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 10266 3740 10406
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9042 3556 9862
rect 3896 9722 3924 11086
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9674 4016 10950
rect 4080 10810 4108 11750
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 4080 10606 4108 10639
rect 4172 10606 4200 12582
rect 4264 12306 4292 12718
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12374 4568 12650
rect 4632 12374 4660 12786
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4632 12238 4660 12310
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4285 11996 4593 12005
rect 4285 11994 4291 11996
rect 4347 11994 4371 11996
rect 4427 11994 4451 11996
rect 4507 11994 4531 11996
rect 4587 11994 4593 11996
rect 4347 11942 4349 11994
rect 4529 11942 4531 11994
rect 4285 11940 4291 11942
rect 4347 11940 4371 11942
rect 4427 11940 4451 11942
rect 4507 11940 4531 11942
rect 4587 11940 4593 11942
rect 4285 11931 4593 11940
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4448 11354 4476 11766
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4540 11234 4568 11834
rect 4632 11354 4660 12038
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4540 11206 4660 11234
rect 4285 10908 4593 10917
rect 4285 10906 4291 10908
rect 4347 10906 4371 10908
rect 4427 10906 4451 10908
rect 4507 10906 4531 10908
rect 4587 10906 4593 10908
rect 4347 10854 4349 10906
rect 4529 10854 4531 10906
rect 4285 10852 4291 10854
rect 4347 10852 4371 10854
rect 4427 10852 4451 10854
rect 4507 10852 4531 10854
rect 4587 10852 4593 10854
rect 4285 10843 4593 10852
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4285 9820 4593 9829
rect 4285 9818 4291 9820
rect 4347 9818 4371 9820
rect 4427 9818 4451 9820
rect 4507 9818 4531 9820
rect 4587 9818 4593 9820
rect 4347 9766 4349 9818
rect 4529 9766 4531 9818
rect 4285 9764 4291 9766
rect 4347 9764 4371 9766
rect 4427 9764 4451 9766
rect 4507 9764 4531 9766
rect 4587 9764 4593 9766
rect 4285 9755 4593 9764
rect 3896 9110 3924 9658
rect 3988 9646 4200 9674
rect 4172 9450 4200 9646
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4540 9178 4568 9454
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7002 3464 8230
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3424 6860 3476 6866
rect 3528 6848 3556 7822
rect 3476 6820 3556 6848
rect 3424 6802 3476 6808
rect 3620 6730 3648 8842
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 8634 4016 8774
rect 4172 8634 4200 8910
rect 4632 8838 4660 11206
rect 4724 9518 4752 13280
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11898 4844 12174
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4816 10606 4844 11834
rect 4908 11558 4936 12650
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 11082 4936 11154
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9217 4752 9318
rect 4710 9208 4766 9217
rect 4710 9143 4766 9152
rect 4816 8974 4844 10406
rect 4908 10130 4936 10746
rect 5000 10266 5028 15302
rect 5184 13870 5212 15846
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5170 12880 5226 12889
rect 5170 12815 5226 12824
rect 5184 12646 5212 12815
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11132 5120 12242
rect 5172 11280 5224 11286
rect 5276 11268 5304 16458
rect 5368 16454 5396 17734
rect 5448 17672 5500 17678
rect 5446 17640 5448 17649
rect 5500 17640 5502 17649
rect 5446 17575 5502 17584
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5354 16144 5410 16153
rect 5552 16114 5580 19858
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5644 18426 5672 19110
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5736 18426 5764 18702
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5828 17882 5856 20946
rect 6288 20942 6316 21490
rect 6380 21350 6408 21626
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 19174 6040 19246
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 5906 18728 5962 18737
rect 5906 18663 5962 18672
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5644 17338 5672 17750
rect 5920 17626 5948 18663
rect 6012 18086 6040 19110
rect 6104 18222 6132 20742
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 18952 6224 19790
rect 6288 19378 6316 20878
rect 6380 20777 6408 21286
rect 6458 21176 6514 21185
rect 6656 21146 6684 21422
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 6458 21111 6460 21120
rect 6512 21111 6514 21120
rect 6644 21140 6696 21146
rect 6460 21082 6512 21088
rect 6644 21082 6696 21088
rect 6366 20768 6422 20777
rect 6366 20703 6422 20712
rect 6472 20262 6500 21082
rect 6932 21010 6960 21354
rect 7024 21078 7052 21354
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6932 20262 6960 20946
rect 7208 20466 7236 21286
rect 7300 20942 7328 21354
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19990 6960 20198
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6550 19544 6606 19553
rect 6550 19479 6606 19488
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6564 19174 6592 19479
rect 6656 19281 6684 19790
rect 6932 19718 6960 19926
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6642 19272 6698 19281
rect 6642 19207 6644 19216
rect 6696 19207 6698 19216
rect 6644 19178 6696 19184
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6276 18964 6328 18970
rect 6196 18924 6276 18952
rect 6196 18222 6224 18924
rect 6276 18906 6328 18912
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6184 18216 6236 18222
rect 6472 18193 6500 18566
rect 6184 18158 6236 18164
rect 6458 18184 6514 18193
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5736 17598 5948 17626
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16726 5672 16934
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5354 16079 5410 16088
rect 5540 16108 5592 16114
rect 5368 16046 5396 16079
rect 5540 16050 5592 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15706 5396 15982
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5552 15162 5580 16050
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5552 14482 5580 15098
rect 5644 14618 5672 15914
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5368 12442 5396 14010
rect 5552 13938 5580 14418
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5552 13530 5580 13874
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5460 12714 5488 12854
rect 5644 12782 5672 13262
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5354 12336 5410 12345
rect 5354 12271 5410 12280
rect 5368 12102 5396 12271
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5224 11240 5304 11268
rect 5356 11280 5408 11286
rect 5172 11222 5224 11228
rect 5356 11222 5408 11228
rect 5092 11104 5212 11132
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 9994 4936 10066
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4285 8732 4593 8741
rect 4285 8730 4291 8732
rect 4347 8730 4371 8732
rect 4427 8730 4451 8732
rect 4507 8730 4531 8732
rect 4587 8730 4593 8732
rect 4347 8678 4349 8730
rect 4529 8678 4531 8730
rect 4285 8676 4291 8678
rect 4347 8676 4371 8678
rect 4427 8676 4451 8678
rect 4507 8676 4531 8678
rect 4587 8676 4593 8678
rect 4285 8667 4593 8676
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3712 6322 3740 8026
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7546 3832 7686
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3792 7404 3844 7410
rect 3896 7392 3924 8434
rect 4264 8362 4292 8570
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3844 7364 3924 7392
rect 3792 7346 3844 7352
rect 3700 6316 3752 6322
rect 3804 6304 3832 7346
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3896 7041 3924 7142
rect 3882 7032 3938 7041
rect 3988 7002 4016 7754
rect 3882 6967 3938 6976
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4080 6662 4108 8055
rect 4285 7644 4593 7653
rect 4285 7642 4291 7644
rect 4347 7642 4371 7644
rect 4427 7642 4451 7644
rect 4507 7642 4531 7644
rect 4587 7642 4593 7644
rect 4347 7590 4349 7642
rect 4529 7590 4531 7642
rect 4285 7588 4291 7590
rect 4347 7588 4371 7590
rect 4427 7588 4451 7590
rect 4507 7588 4531 7590
rect 4587 7588 4593 7590
rect 4285 7579 4593 7588
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6390 4108 6598
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3884 6316 3936 6322
rect 3804 6276 3884 6304
rect 3700 6258 3752 6264
rect 3884 6258 3936 6264
rect 3712 5896 3740 6258
rect 3792 5908 3844 5914
rect 3712 5868 3792 5896
rect 3792 5850 3844 5856
rect 3896 5710 3924 6258
rect 3974 6216 4030 6225
rect 3974 6151 3976 6160
rect 4028 6151 4030 6160
rect 3976 6122 4028 6128
rect 4172 6118 4200 7278
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4540 6798 4568 7210
rect 4528 6792 4580 6798
rect 4526 6760 4528 6769
rect 4580 6760 4582 6769
rect 4526 6695 4582 6704
rect 4285 6556 4593 6565
rect 4285 6554 4291 6556
rect 4347 6554 4371 6556
rect 4427 6554 4451 6556
rect 4507 6554 4531 6556
rect 4587 6554 4593 6556
rect 4347 6502 4349 6554
rect 4529 6502 4531 6554
rect 4285 6500 4291 6502
rect 4347 6500 4371 6502
rect 4427 6500 4451 6502
rect 4507 6500 4531 6502
rect 4587 6500 4593 6502
rect 4285 6491 4593 6500
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4264 5778 4292 6394
rect 4632 6254 4660 8230
rect 4724 7750 4752 8298
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4816 7478 4844 8774
rect 4908 8634 4936 9930
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5000 9042 5028 9590
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7546 4936 7686
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3344 4622 3372 4966
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3344 3942 3372 4558
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3252 3194 3280 3878
rect 3712 3194 3740 3878
rect 3804 3534 3832 5510
rect 3896 5234 3924 5646
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4080 5030 4108 5714
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5234 4200 5510
rect 4285 5468 4593 5477
rect 4285 5466 4291 5468
rect 4347 5466 4371 5468
rect 4427 5466 4451 5468
rect 4507 5466 4531 5468
rect 4587 5466 4593 5468
rect 4347 5414 4349 5466
rect 4529 5414 4531 5466
rect 4285 5412 4291 5414
rect 4347 5412 4371 5414
rect 4427 5412 4451 5414
rect 4507 5412 4531 5414
rect 4587 5412 4593 5414
rect 4285 5403 4593 5412
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4758 4108 4966
rect 4632 4826 4660 5714
rect 4724 5098 4752 7142
rect 4816 6848 4844 7278
rect 4896 7268 4948 7274
rect 5000 7256 5028 8774
rect 4948 7228 5028 7256
rect 4896 7210 4948 7216
rect 4988 6860 5040 6866
rect 4816 6820 4936 6848
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6338 4844 6666
rect 4908 6440 4936 6820
rect 4988 6802 5040 6808
rect 5000 6633 5028 6802
rect 5092 6662 5120 10406
rect 5184 9625 5212 11104
rect 5262 11112 5318 11121
rect 5262 11047 5318 11056
rect 5276 10266 5304 11047
rect 5368 10470 5396 11222
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 10130 5396 10406
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5170 9616 5226 9625
rect 5170 9551 5226 9560
rect 5184 9518 5212 9551
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8945 5212 8978
rect 5170 8936 5226 8945
rect 5170 8871 5226 8880
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5080 6656 5132 6662
rect 4986 6624 5042 6633
rect 5080 6598 5132 6604
rect 4986 6559 5042 6568
rect 4908 6412 5028 6440
rect 4816 6310 4936 6338
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5914 4844 6190
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4908 5658 4936 6310
rect 4816 5630 4936 5658
rect 5000 5642 5028 6412
rect 5184 6254 5212 8230
rect 5276 7954 5304 9318
rect 5368 8294 5396 10066
rect 5460 9450 5488 12650
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10810 5580 10950
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5540 9172 5592 9178
rect 5644 9160 5672 11154
rect 5592 9132 5672 9160
rect 5540 9114 5592 9120
rect 5552 8362 5580 9114
rect 5736 9081 5764 17598
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17338 5948 17478
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6196 17202 6224 18158
rect 6458 18119 6514 18128
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6104 15706 6132 15914
rect 6196 15706 6224 17138
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5828 13530 5856 13738
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11762 6040 12038
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11218 5856 11494
rect 5816 11212 5868 11218
rect 5868 11172 5948 11200
rect 5816 11154 5868 11160
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5722 9072 5778 9081
rect 5722 9007 5778 9016
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8401 5672 8910
rect 5630 8392 5686 8401
rect 5540 8356 5592 8362
rect 5630 8327 5686 8336
rect 5540 8298 5592 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7002 5304 7754
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5276 6662 5304 6802
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5368 6458 5396 7890
rect 5460 7857 5488 7890
rect 5446 7848 5502 7857
rect 5446 7783 5502 7792
rect 5448 7744 5500 7750
rect 5446 7712 5448 7721
rect 5500 7712 5502 7721
rect 5446 7647 5502 7656
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 7177 5488 7346
rect 5446 7168 5502 7177
rect 5446 7103 5502 7112
rect 5460 6905 5488 7103
rect 5552 7002 5580 8298
rect 5736 7954 5764 9007
rect 5828 7954 5856 11018
rect 5920 10810 5948 11172
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6104 9489 6132 14554
rect 6288 14482 6316 14758
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6380 13394 6408 13874
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6288 12986 6316 13330
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6472 12866 6500 17614
rect 6564 15450 6592 19110
rect 6932 18766 6960 19654
rect 7392 19310 7420 21354
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 8956 21146 8984 21286
rect 9048 21146 9076 21490
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 7930 20632 7986 20641
rect 7930 20567 7986 20576
rect 8666 20632 8722 20641
rect 8666 20567 8668 20576
rect 7838 20496 7894 20505
rect 7838 20431 7840 20440
rect 7892 20431 7894 20440
rect 7840 20402 7892 20408
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7484 19174 7512 19926
rect 7852 19922 7880 20198
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7944 19446 7972 20567
rect 8720 20567 8722 20576
rect 8668 20538 8720 20544
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 8036 19310 8064 20470
rect 9048 20330 9076 20878
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6642 16688 6698 16697
rect 6642 16623 6698 16632
rect 6656 15706 6684 16623
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6748 15570 6776 17478
rect 6840 15570 6868 17818
rect 6932 17134 6960 18702
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7208 17814 7236 18022
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 7116 16590 7144 17614
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 7012 15564 7064 15570
rect 7116 15552 7144 16526
rect 7064 15524 7144 15552
rect 7012 15506 7064 15512
rect 6564 15422 6776 15450
rect 6288 12838 6500 12866
rect 6288 12442 6316 12838
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10674 6224 11086
rect 6288 10792 6316 12378
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6380 11762 6408 12310
rect 6368 11756 6420 11762
rect 6420 11716 6500 11744
rect 6368 11698 6420 11704
rect 6288 10764 6408 10792
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6288 9722 6316 10610
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6182 9616 6238 9625
rect 6182 9551 6238 9560
rect 6090 9480 6146 9489
rect 6012 9438 6090 9466
rect 5906 7984 5962 7993
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5816 7948 5868 7954
rect 5906 7919 5962 7928
rect 5816 7890 5868 7896
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 5540 6792 5592 6798
rect 5446 6760 5502 6769
rect 5540 6734 5592 6740
rect 5446 6695 5448 6704
rect 5500 6695 5502 6704
rect 5448 6666 5500 6672
rect 5552 6458 5580 6734
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 6254 5672 7210
rect 5736 6730 5764 7686
rect 5920 7546 5948 7919
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5828 6934 5856 7278
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5828 6497 5856 6734
rect 5814 6488 5870 6497
rect 5814 6423 5870 6432
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5914 5212 6054
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 4988 5636 5040 5642
rect 4816 5370 4844 5630
rect 4988 5578 5040 5584
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3896 4214 3924 4490
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3896 3602 3924 4150
rect 4080 4078 4108 4694
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4285 4380 4593 4389
rect 4285 4378 4291 4380
rect 4347 4378 4371 4380
rect 4427 4378 4451 4380
rect 4507 4378 4531 4380
rect 4587 4378 4593 4380
rect 4347 4326 4349 4378
rect 4529 4326 4531 4378
rect 4285 4324 4291 4326
rect 4347 4324 4371 4326
rect 4427 4324 4451 4326
rect 4507 4324 4531 4326
rect 4587 4324 4593 4326
rect 4285 4315 4593 4324
rect 4632 4282 4660 4422
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4080 3670 4108 4014
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 3670 4292 3878
rect 4540 3738 4568 4014
rect 4816 3738 4844 5170
rect 4908 4010 4936 5510
rect 5276 4826 5304 5714
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 5644 3534 5672 6190
rect 6012 5914 6040 9438
rect 6090 9415 6146 9424
rect 6090 8800 6146 8809
rect 6090 8735 6146 8744
rect 6104 7342 6132 8735
rect 6196 7342 6224 9551
rect 6380 9110 6408 10764
rect 6472 9654 6500 11716
rect 6564 11626 6592 12582
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6564 11286 6592 11562
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6550 10568 6606 10577
rect 6550 10503 6606 10512
rect 6564 9654 6592 10503
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6472 9042 6500 9454
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 7834 6408 8910
rect 6472 8129 6500 8978
rect 6748 8922 6776 15422
rect 6840 15026 6868 15506
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 13870 6960 14894
rect 7024 14278 7052 15506
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14618 7144 14758
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7116 14090 7144 14418
rect 7024 14062 7144 14090
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13462 6960 13806
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11014 6868 11494
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10606 6868 10950
rect 6932 10674 6960 12786
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6932 10033 6960 10610
rect 7024 10266 7052 14062
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7116 11665 7144 12650
rect 7102 11656 7158 11665
rect 7102 11591 7158 11600
rect 7208 11234 7236 17750
rect 7392 17728 7420 18566
rect 7484 18154 7512 19110
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7654 18320 7710 18329
rect 7654 18255 7710 18264
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7472 17740 7524 17746
rect 7392 17700 7472 17728
rect 7472 17682 7524 17688
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7300 16114 7328 17614
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7392 16046 7420 16662
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7392 14958 7420 15982
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7484 14482 7512 17682
rect 7668 17202 7696 18255
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7760 17882 7788 18090
rect 7852 18086 7880 18838
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7840 17536 7892 17542
rect 7838 17504 7840 17513
rect 7892 17504 7894 17513
rect 7838 17439 7894 17448
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7116 11206 7236 11234
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6656 8894 6776 8922
rect 6828 8900 6880 8906
rect 6458 8120 6514 8129
rect 6458 8055 6514 8064
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6288 7806 6408 7834
rect 6472 7834 6500 7890
rect 6656 7834 6684 8894
rect 6828 8842 6880 8848
rect 6840 8634 6868 8842
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6734 8528 6790 8537
rect 6734 8463 6790 8472
rect 6748 8294 6776 8463
rect 6932 8430 6960 9862
rect 7024 9722 7052 10066
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7012 9512 7064 9518
rect 7116 9500 7144 11206
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7208 9518 7236 11018
rect 7064 9472 7144 9500
rect 7196 9512 7248 9518
rect 7012 9454 7064 9460
rect 7196 9454 7248 9460
rect 7300 9364 7328 14350
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7576 13734 7604 14486
rect 7668 14414 7696 17138
rect 7944 17134 7972 19178
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 8392 18964 8444 18970
rect 8588 18952 8616 20198
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18970 8708 19110
rect 8444 18924 8616 18952
rect 8668 18964 8720 18970
rect 8392 18906 8444 18912
rect 8668 18906 8720 18912
rect 8404 18834 8432 18906
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8312 18136 8340 18294
rect 8404 18290 8432 18770
rect 8680 18630 8708 18770
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8036 18108 8340 18136
rect 8576 18148 8628 18154
rect 8036 17882 8064 18108
rect 8576 18090 8628 18096
rect 8588 18057 8616 18090
rect 8574 18048 8630 18057
rect 8172 17980 8480 17989
rect 8574 17983 8630 17992
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8300 17808 8352 17814
rect 8114 17776 8170 17785
rect 8300 17750 8352 17756
rect 8114 17711 8170 17720
rect 8128 17338 8156 17711
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 17338 8248 17478
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8312 17134 8340 17750
rect 8680 17660 8708 17818
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8588 17632 8708 17660
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 7932 17128 7984 17134
rect 8300 17128 8352 17134
rect 7932 17070 7984 17076
rect 8036 17088 8300 17116
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7760 16794 7788 16934
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7852 16658 7880 16934
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7668 13841 7696 14350
rect 7654 13832 7710 13841
rect 7654 13767 7710 13776
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7392 13190 7420 13670
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 11830 7420 12242
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7392 11082 7420 11766
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7484 10810 7512 12174
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7576 10470 7604 13670
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7668 12850 7696 12922
rect 7760 12850 7788 16050
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11898 7788 12174
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7852 11218 7880 16594
rect 7944 15638 7972 17070
rect 8036 16046 8064 17088
rect 8496 17105 8524 17546
rect 8300 17070 8352 17076
rect 8482 17096 8538 17105
rect 8588 17066 8616 17632
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8482 17031 8538 17040
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8482 16416 8538 16425
rect 8482 16351 8538 16360
rect 8496 16046 8524 16351
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8036 15570 8064 15982
rect 8588 15910 8616 16730
rect 8680 16182 8708 17478
rect 8772 17338 8800 17682
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8772 16590 8800 17002
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8772 16250 8800 16526
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 8588 15688 8616 15846
rect 8404 15660 8616 15688
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8404 15201 8432 15660
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8390 15192 8446 15201
rect 8390 15127 8446 15136
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14618 7972 14894
rect 8496 14890 8524 15506
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8574 15192 8630 15201
rect 8574 15127 8630 15136
rect 8588 15026 8616 15127
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 12986 7972 13670
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7944 12753 7972 12922
rect 7930 12744 7986 12753
rect 7930 12679 7986 12688
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 11694 7972 12582
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7668 10606 7696 11154
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7748 10736 7800 10742
rect 7746 10704 7748 10713
rect 7800 10704 7802 10713
rect 7746 10639 7802 10648
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9625 7420 9862
rect 7378 9616 7434 9625
rect 7378 9551 7434 9560
rect 7392 9518 7420 9551
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7116 9336 7328 9364
rect 7012 9036 7064 9042
rect 7116 9024 7144 9336
rect 7194 9208 7250 9217
rect 7194 9143 7250 9152
rect 7064 8996 7144 9024
rect 7012 8978 7064 8984
rect 7102 8936 7158 8945
rect 7102 8871 7104 8880
rect 7156 8871 7158 8880
rect 7104 8842 7156 8848
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6748 7954 6776 8230
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6472 7806 6592 7834
rect 6656 7806 6776 7834
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6288 7188 6316 7806
rect 6564 7290 6592 7806
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7478 6684 7686
rect 6748 7546 6776 7806
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6748 7313 6776 7482
rect 6734 7304 6790 7313
rect 6564 7262 6684 7290
rect 6196 7160 6316 7188
rect 6552 7200 6604 7206
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6012 5778 6040 5850
rect 6104 5817 6132 6598
rect 6090 5808 6146 5817
rect 6000 5772 6052 5778
rect 6196 5778 6224 7160
rect 6552 7142 6604 7148
rect 6564 7002 6592 7142
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 5914 6316 6598
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6090 5743 6146 5752
rect 6184 5772 6236 5778
rect 6000 5714 6052 5720
rect 6184 5714 6236 5720
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6012 4758 6040 5102
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3804 3058 3832 3470
rect 4285 3292 4593 3301
rect 4285 3290 4291 3292
rect 4347 3290 4371 3292
rect 4427 3290 4451 3292
rect 4507 3290 4531 3292
rect 4587 3290 4593 3292
rect 4347 3238 4349 3290
rect 4529 3238 4531 3290
rect 4285 3236 4291 3238
rect 4347 3236 4371 3238
rect 4427 3236 4451 3238
rect 4507 3236 4531 3238
rect 4587 3236 4593 3238
rect 4285 3227 4593 3236
rect 5828 3194 5856 4626
rect 6104 4146 6132 5578
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6196 4486 6224 5034
rect 6564 4758 6592 6938
rect 6656 6633 6684 7262
rect 6734 7239 6790 7248
rect 6840 6882 6868 7890
rect 6748 6854 6868 6882
rect 6642 6624 6698 6633
rect 6642 6559 6698 6568
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5920 3670 5948 4014
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6196 3670 6224 3946
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6656 3398 6684 4558
rect 6748 4282 6776 6854
rect 6932 6798 6960 8366
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 8090 7052 8298
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7010 7984 7066 7993
rect 7010 7919 7012 7928
rect 7064 7919 7066 7928
rect 7012 7890 7064 7896
rect 7116 7834 7144 8570
rect 7208 7970 7236 9143
rect 7484 9042 7512 9998
rect 7576 9654 7604 10202
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7300 8401 7328 8978
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7484 8072 7512 8774
rect 7576 8634 7604 9318
rect 7668 9178 7696 10542
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7668 8430 7696 8978
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7392 8044 7512 8072
rect 7564 8084 7616 8090
rect 7208 7942 7328 7970
rect 7012 7812 7064 7818
rect 7116 7806 7236 7834
rect 7012 7754 7064 7760
rect 7024 7546 7052 7754
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 7410 7144 7686
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7208 7290 7236 7806
rect 7300 7410 7328 7942
rect 7392 7886 7420 8044
rect 7564 8026 7616 8032
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7116 7262 7236 7290
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6840 5370 6868 6734
rect 6932 6322 6960 6734
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6918 5944 6974 5953
rect 6918 5879 6920 5888
rect 6972 5879 6974 5888
rect 6920 5850 6972 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7024 4622 7052 5714
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6748 3058 6776 4218
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 3194 6868 3674
rect 7024 3670 7052 4422
rect 7116 4078 7144 7262
rect 7196 7200 7248 7206
rect 7300 7177 7328 7346
rect 7196 7142 7248 7148
rect 7286 7168 7342 7177
rect 7208 6254 7236 7142
rect 7286 7103 7342 7112
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7300 6458 7328 6938
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5098 7236 6190
rect 7392 5914 7420 7686
rect 7484 7274 7512 7822
rect 7576 7342 7604 8026
rect 7668 8022 7696 8230
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7484 7002 7512 7210
rect 7668 7206 7696 7958
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7576 7002 7604 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7760 6882 7788 10639
rect 7852 7478 7880 10950
rect 7944 10062 7972 11154
rect 8036 10538 8064 14826
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8312 14006 8340 14350
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8404 13716 8432 14418
rect 8496 14278 8524 14418
rect 8588 14362 8616 14962
rect 8680 14618 8708 15302
rect 8772 14958 8800 16186
rect 8864 15162 8892 20266
rect 9048 20058 9076 20266
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8956 17338 8984 19790
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9048 19242 9076 19450
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9036 18760 9088 18766
rect 9140 18737 9168 21286
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9416 20398 9444 21082
rect 9692 20942 9720 21422
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9784 20874 9812 21490
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9968 20466 9996 20878
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 10152 20262 10180 21898
rect 10336 21010 10364 21898
rect 12059 21788 12367 21797
rect 12059 21786 12065 21788
rect 12121 21786 12145 21788
rect 12201 21786 12225 21788
rect 12281 21786 12305 21788
rect 12361 21786 12367 21788
rect 12121 21734 12123 21786
rect 12303 21734 12305 21786
rect 12059 21732 12065 21734
rect 12121 21732 12145 21734
rect 12201 21732 12225 21734
rect 12281 21732 12305 21734
rect 12361 21732 12367 21734
rect 12059 21723 12367 21732
rect 12544 21690 12572 21927
rect 13358 21720 13414 21729
rect 12532 21684 12584 21690
rect 13358 21655 13414 21664
rect 12532 21626 12584 21632
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10414 21040 10470 21049
rect 10324 21004 10376 21010
rect 10414 20975 10470 20984
rect 10324 20946 10376 20952
rect 10336 20777 10364 20946
rect 10322 20768 10378 20777
rect 10322 20703 10378 20712
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9508 19417 9536 19722
rect 10060 19514 10088 19858
rect 10152 19689 10180 20198
rect 10428 20058 10456 20975
rect 10520 20602 10548 21422
rect 12360 21418 12388 21558
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 11256 21010 11284 21354
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10612 20262 10640 20946
rect 10796 20806 10824 20946
rect 10888 20874 11100 20890
rect 10876 20868 11100 20874
rect 10928 20862 11100 20868
rect 10876 20810 10928 20816
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10796 19961 10824 20402
rect 10782 19952 10838 19961
rect 10980 19922 11008 20742
rect 10782 19887 10838 19896
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10138 19680 10194 19689
rect 10138 19615 10194 19624
rect 10244 19514 10272 19722
rect 11072 19718 11100 20862
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 9494 19408 9550 19417
rect 10046 19408 10102 19417
rect 9494 19343 9550 19352
rect 9956 19372 10008 19378
rect 10046 19343 10102 19352
rect 9956 19314 10008 19320
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 18970 9904 19178
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9036 18702 9088 18708
rect 9126 18728 9182 18737
rect 9048 18329 9076 18702
rect 9126 18663 9182 18672
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9034 18320 9090 18329
rect 9034 18255 9090 18264
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 15910 8984 16526
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8956 15042 8984 15846
rect 8864 15014 8984 15042
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8680 14464 8708 14554
rect 8680 14436 8800 14464
rect 8588 14334 8708 14362
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8574 13968 8630 13977
rect 8574 13903 8630 13912
rect 8588 13870 8616 13903
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8404 13688 8616 13716
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 8392 13524 8444 13530
rect 8588 13512 8616 13688
rect 8392 13466 8444 13472
rect 8496 13484 8616 13512
rect 8404 13297 8432 13466
rect 8390 13288 8446 13297
rect 8390 13223 8446 13232
rect 8496 13190 8524 13484
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8588 13190 8616 13330
rect 8680 13258 8708 14334
rect 8772 13462 8800 14436
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8300 13184 8352 13190
rect 8114 13152 8170 13161
rect 8300 13126 8352 13132
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8114 13087 8170 13096
rect 8128 12850 8156 13087
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8312 12714 8340 13126
rect 8496 13002 8524 13126
rect 8496 12974 8708 13002
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8496 11540 8524 12310
rect 8496 11512 8616 11540
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8588 11234 8616 11512
rect 8680 11506 8708 12974
rect 8864 12782 8892 15014
rect 8944 14952 8996 14958
rect 8942 14920 8944 14929
rect 8996 14920 8998 14929
rect 8942 14855 8998 14864
rect 9048 14822 9076 17818
rect 9140 17134 9168 18566
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9404 17808 9456 17814
rect 9324 17768 9404 17796
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9232 17377 9260 17682
rect 9218 17368 9274 17377
rect 9218 17303 9274 17312
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 15570 9168 16390
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12442 8800 12582
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8772 11626 8800 12378
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8680 11478 8800 11506
rect 8588 11206 8708 11234
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 10180 8064 10474
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10192 8260 10198
rect 8036 10160 8208 10180
rect 8260 10160 8262 10169
rect 8036 10152 8206 10160
rect 8206 10095 8262 10104
rect 7932 10056 7984 10062
rect 8312 10033 8340 10202
rect 7932 9998 7984 10004
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 8809 7972 9522
rect 8036 9382 8064 9658
rect 8312 9518 8340 9959
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 9217 8064 9318
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8022 9208 8078 9217
rect 8172 9211 8480 9220
rect 8022 9143 8078 9152
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8496 8945 8524 9114
rect 8588 9110 8616 11018
rect 8680 10713 8708 11206
rect 8666 10704 8722 10713
rect 8666 10639 8722 10648
rect 8680 10130 8708 10639
rect 8772 10606 8800 11478
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8772 10062 8800 10406
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8114 8936 8170 8945
rect 8024 8900 8076 8906
rect 8114 8871 8116 8880
rect 8024 8842 8076 8848
rect 8168 8871 8170 8880
rect 8482 8936 8538 8945
rect 8482 8871 8538 8880
rect 8576 8900 8628 8906
rect 8116 8842 8168 8848
rect 7930 8800 7986 8809
rect 7930 8735 7986 8744
rect 7930 8664 7986 8673
rect 8036 8634 8064 8842
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8634 8432 8774
rect 7930 8599 7986 8608
rect 8024 8628 8076 8634
rect 7944 7818 7972 8599
rect 8024 8570 8076 8576
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8036 7954 8064 8570
rect 8390 8528 8446 8537
rect 8390 8463 8392 8472
rect 8444 8463 8446 8472
rect 8392 8434 8444 8440
rect 8390 8392 8446 8401
rect 8390 8327 8392 8336
rect 8444 8327 8446 8336
rect 8392 8298 8444 8304
rect 8496 8294 8524 8871
rect 8576 8842 8628 8848
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 8300 8016 8352 8022
rect 8588 7993 8616 8842
rect 8680 8498 8708 9318
rect 8772 8906 8800 9998
rect 8864 9654 8892 11630
rect 8956 11218 8984 13874
rect 9048 13394 9076 14418
rect 9140 14278 9168 15030
rect 9232 14618 9260 17303
rect 9324 16969 9352 17768
rect 9404 17750 9456 17756
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9310 16960 9366 16969
rect 9310 16895 9366 16904
rect 9416 16833 9444 17070
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9324 16250 9352 16526
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 16250 9444 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15706 9352 15982
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9416 15706 9444 15914
rect 9508 15706 9536 17546
rect 9600 16794 9628 17682
rect 9692 17338 9720 18022
rect 9784 17796 9812 18906
rect 9968 18766 9996 19314
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18329 9996 18702
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9956 18216 10008 18222
rect 10060 18204 10088 19343
rect 10612 19310 10640 19654
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10600 19304 10652 19310
rect 10704 19281 10732 19450
rect 10980 19310 11008 19654
rect 10968 19304 11020 19310
rect 10600 19246 10652 19252
rect 10690 19272 10746 19281
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10008 18176 10088 18204
rect 9956 18158 10008 18164
rect 10152 17921 10180 18838
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 18358 10364 18770
rect 10612 18748 10640 19246
rect 10968 19246 11020 19252
rect 10690 19207 10746 19216
rect 11072 18834 11100 19654
rect 11164 19553 11192 19858
rect 11150 19544 11206 19553
rect 11150 19479 11206 19488
rect 11256 19334 11284 20946
rect 11164 19306 11284 19334
rect 11164 19009 11192 19306
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11150 19000 11206 19009
rect 11256 18970 11284 19110
rect 11150 18935 11206 18944
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10692 18760 10744 18766
rect 10612 18720 10692 18748
rect 10692 18702 10744 18708
rect 11058 18728 11114 18737
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10336 18222 10364 18294
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10138 17912 10194 17921
rect 9956 17876 10008 17882
rect 10138 17847 10194 17856
rect 9956 17818 10008 17824
rect 9864 17808 9916 17814
rect 9784 17768 9864 17796
rect 9864 17750 9916 17756
rect 9968 17626 9996 17818
rect 10138 17776 10194 17785
rect 10138 17711 10140 17720
rect 10192 17711 10194 17720
rect 10140 17682 10192 17688
rect 9784 17598 9996 17626
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9784 17202 9812 17598
rect 10152 17338 10180 17682
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10244 17270 10272 17546
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9876 17082 9904 17206
rect 10336 17134 10364 18158
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10428 17882 10456 18022
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10520 17746 10548 18362
rect 10704 18222 10732 18702
rect 10968 18692 11020 18698
rect 11058 18663 11060 18672
rect 10968 18634 11020 18640
rect 11112 18663 11114 18672
rect 11060 18634 11112 18640
rect 10980 18426 11008 18634
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17882 10640 18022
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10506 17368 10562 17377
rect 10416 17332 10468 17338
rect 10612 17354 10640 17682
rect 10704 17610 10732 18158
rect 10968 18080 11020 18086
rect 10874 18048 10930 18057
rect 10968 18022 11020 18028
rect 10874 17983 10930 17992
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10562 17326 10640 17354
rect 10506 17303 10562 17312
rect 10416 17274 10468 17280
rect 9956 17128 10008 17134
rect 9876 17076 9956 17082
rect 9876 17070 10008 17076
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9876 17054 9996 17070
rect 9784 16794 9812 17002
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9784 16590 9812 16730
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9692 16250 9720 16526
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9588 16040 9640 16046
rect 9640 16000 9720 16028
rect 9588 15982 9640 15988
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9600 15586 9628 15642
rect 9692 15609 9720 16000
rect 9324 15558 9628 15586
rect 9678 15600 9734 15609
rect 9324 15434 9352 15558
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9310 15192 9366 15201
rect 9310 15127 9366 15136
rect 9324 14958 9352 15127
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14618 9352 14758
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9232 14278 9260 14554
rect 9416 14346 9444 15370
rect 9508 15042 9536 15558
rect 9678 15535 9734 15544
rect 9784 15502 9812 16526
rect 9876 16250 9904 17054
rect 10048 16788 10100 16794
rect 10152 16776 10180 17070
rect 10100 16748 10180 16776
rect 10048 16730 10100 16736
rect 9956 16652 10008 16658
rect 10008 16612 10180 16640
rect 9956 16594 10008 16600
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9508 15026 9628 15042
rect 9508 15020 9640 15026
rect 9508 15014 9588 15020
rect 9588 14962 9640 14968
rect 9784 14958 9812 15438
rect 9876 15434 9904 16186
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15638 9996 15914
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9954 15464 10010 15473
rect 9864 15428 9916 15434
rect 9954 15399 10010 15408
rect 9864 15370 9916 15376
rect 9876 14958 9904 15370
rect 9968 15026 9996 15399
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9508 14618 9536 14894
rect 9770 14784 9826 14793
rect 9770 14719 9826 14728
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9140 13870 9168 14214
rect 9416 13870 9444 14282
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9508 13870 9536 13942
rect 9600 13870 9628 14486
rect 9784 14414 9812 14719
rect 9876 14498 9904 14894
rect 10060 14618 10088 14894
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9876 14470 9996 14498
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9864 14408 9916 14414
rect 9968 14385 9996 14470
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9864 14350 9916 14356
rect 9954 14376 10010 14385
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13938 9720 14214
rect 9876 14006 9904 14350
rect 9954 14311 10010 14320
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9128 13864 9180 13870
rect 9404 13864 9456 13870
rect 9180 13824 9260 13852
rect 9128 13806 9180 13812
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13462 9168 13670
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9232 13258 9260 13824
rect 9404 13806 9456 13812
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9048 12646 9076 13194
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9140 12374 9168 12786
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9126 12200 9182 12209
rect 9126 12135 9182 12144
rect 9140 11898 9168 12135
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11665 9076 11698
rect 9034 11656 9090 11665
rect 9034 11591 9090 11600
rect 9232 11558 9260 12922
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9416 12442 9444 13806
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9508 12986 9536 13398
rect 9588 13388 9640 13394
rect 9692 13376 9720 13874
rect 9956 13864 10008 13870
rect 9954 13832 9956 13841
rect 10008 13832 10010 13841
rect 9954 13767 10010 13776
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9772 13524 9824 13530
rect 9824 13484 9904 13512
rect 9772 13466 9824 13472
rect 9640 13348 9720 13376
rect 9588 13330 9640 13336
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9600 12918 9628 13330
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9324 11694 9352 12242
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10985 8984 11018
rect 8942 10976 8998 10985
rect 8942 10911 8998 10920
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 9722 8984 10542
rect 9048 10266 9076 11494
rect 9416 11336 9444 12242
rect 9508 11898 9536 12718
rect 9600 12374 9628 12854
rect 9876 12628 9904 13484
rect 9968 12753 9996 13631
rect 10060 13394 10088 14418
rect 10152 14346 10180 16612
rect 10244 16522 10272 17070
rect 10428 16776 10456 17274
rect 10612 16794 10640 17326
rect 10796 17218 10824 17682
rect 10888 17542 10916 17983
rect 10980 17814 11008 18022
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10876 17536 10928 17542
rect 10980 17513 11008 17750
rect 10876 17478 10928 17484
rect 10966 17504 11022 17513
rect 10966 17439 11022 17448
rect 10874 17232 10930 17241
rect 10692 17196 10744 17202
rect 10796 17190 10874 17218
rect 10980 17202 11008 17439
rect 11072 17338 11100 18362
rect 11150 17912 11206 17921
rect 11150 17847 11206 17856
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10874 17167 10930 17176
rect 10968 17196 11020 17202
rect 10692 17138 10744 17144
rect 10968 17138 11020 17144
rect 10336 16748 10456 16776
rect 10600 16788 10652 16794
rect 10336 16658 10364 16748
rect 10600 16730 10652 16736
rect 10598 16688 10654 16697
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10508 16652 10560 16658
rect 10598 16623 10600 16632
rect 10508 16594 10560 16600
rect 10652 16623 10654 16632
rect 10600 16594 10652 16600
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 15162 10272 15438
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10336 14618 10364 16594
rect 10428 16153 10456 16594
rect 10520 16538 10548 16594
rect 10704 16538 10732 17138
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10520 16510 10732 16538
rect 10690 16416 10746 16425
rect 10796 16402 10824 17002
rect 10980 16969 11008 17002
rect 11060 16992 11112 16998
rect 10966 16960 11022 16969
rect 11060 16934 11112 16940
rect 10966 16895 11022 16904
rect 11072 16658 11100 16934
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10746 16374 10916 16402
rect 10690 16351 10746 16360
rect 10888 16250 10916 16374
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10414 16144 10470 16153
rect 10414 16079 10470 16088
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10324 14612 10376 14618
rect 10376 14572 10456 14600
rect 10324 14554 10376 14560
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 13977 10180 14282
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10138 13968 10194 13977
rect 10138 13903 10194 13912
rect 10244 13394 10272 14214
rect 10336 13734 10364 14350
rect 10428 13870 10456 14572
rect 10416 13864 10468 13870
rect 10520 13841 10548 15370
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15026 10732 15302
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10796 14929 10824 15438
rect 10782 14920 10838 14929
rect 10600 14884 10652 14890
rect 10888 14890 10916 15574
rect 10980 15065 11008 16458
rect 11072 16114 11100 16594
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11164 15892 11192 17847
rect 11242 17776 11298 17785
rect 11242 17711 11298 17720
rect 11256 17610 11284 17711
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11256 16130 11284 17274
rect 11348 16250 11376 21354
rect 11428 20936 11480 20942
rect 11426 20904 11428 20913
rect 11520 20936 11572 20942
rect 11480 20904 11482 20913
rect 11520 20878 11572 20884
rect 11426 20839 11482 20848
rect 11532 19854 11560 20878
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11624 20398 11652 20742
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 19922 11652 20198
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11440 19514 11468 19790
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11428 19304 11480 19310
rect 11426 19272 11428 19281
rect 11480 19272 11482 19281
rect 11426 19207 11482 19216
rect 11532 19156 11560 19790
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11440 19128 11560 19156
rect 11624 19145 11652 19178
rect 11610 19136 11666 19145
rect 11440 18358 11468 19128
rect 11610 19071 11666 19080
rect 11518 18864 11574 18873
rect 11518 18799 11574 18808
rect 11612 18828 11664 18834
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11440 17814 11468 18158
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11532 17134 11560 18799
rect 11612 18770 11664 18776
rect 11624 18426 11652 18770
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11624 16998 11652 18158
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11440 16726 11468 16934
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11624 16153 11652 16934
rect 11610 16144 11666 16153
rect 11256 16102 11376 16130
rect 11244 15904 11296 15910
rect 11164 15864 11244 15892
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11072 15434 11100 15642
rect 11164 15570 11192 15864
rect 11244 15846 11296 15852
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11058 15192 11114 15201
rect 11164 15178 11192 15506
rect 11114 15150 11192 15178
rect 11058 15127 11114 15136
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10782 14855 10838 14864
rect 10876 14884 10928 14890
rect 10600 14826 10652 14832
rect 10876 14826 10928 14832
rect 10416 13806 10468 13812
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10428 13530 10456 13670
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10520 13462 10548 13670
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 9954 12744 10010 12753
rect 10060 12714 10088 13330
rect 10140 13320 10192 13326
rect 10138 13288 10140 13297
rect 10192 13288 10194 13297
rect 10138 13223 10194 13232
rect 10232 13184 10284 13190
rect 10508 13184 10560 13190
rect 10232 13126 10284 13132
rect 10506 13152 10508 13161
rect 10560 13152 10562 13161
rect 9954 12679 10010 12688
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9956 12640 10008 12646
rect 9876 12600 9956 12628
rect 9956 12582 10008 12588
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9600 11694 9628 12310
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 11348 9548 11354
rect 9416 11308 9496 11336
rect 9496 11290 9548 11296
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9588 11212 9640 11218
rect 9692 11200 9720 12378
rect 9968 12374 9996 12582
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9640 11172 9720 11200
rect 9588 11154 9640 11160
rect 9140 11014 9168 11154
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8850 9480 8906 9489
rect 8850 9415 8852 9424
rect 8904 9415 8906 9424
rect 8852 9386 8904 9392
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 8906 8984 9318
rect 9048 9110 9076 9522
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8850 8528 8906 8537
rect 8668 8492 8720 8498
rect 8850 8463 8906 8472
rect 8668 8434 8720 8440
rect 8864 8242 8892 8463
rect 8772 8214 8892 8242
rect 8772 8072 8800 8214
rect 8680 8044 8800 8072
rect 8852 8084 8904 8090
rect 8300 7958 8352 7964
rect 8574 7984 8630 7993
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8022 7848 8078 7857
rect 7932 7812 7984 7818
rect 8022 7783 8078 7792
rect 8206 7848 8262 7857
rect 8206 7783 8262 7792
rect 7932 7754 7984 7760
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 8036 7342 8064 7783
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7484 6854 7788 6882
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5710 7512 6854
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7576 6322 7604 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6338 7788 6598
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7668 6310 7788 6338
rect 7838 6352 7894 6361
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4758 7236 5034
rect 7484 4826 7512 5646
rect 7576 5370 7604 6258
rect 7668 5914 7696 6310
rect 7838 6287 7894 6296
rect 7852 6254 7880 6287
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7760 6089 7788 6190
rect 7746 6080 7802 6089
rect 7746 6015 7802 6024
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7944 5658 7972 7278
rect 8128 7256 8156 7686
rect 8220 7478 8248 7783
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8312 7342 8340 7958
rect 8484 7948 8536 7954
rect 8680 7954 8708 8044
rect 8956 8072 8984 8842
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9048 8129 9076 8570
rect 8904 8044 8984 8072
rect 9034 8120 9090 8129
rect 9034 8055 9090 8064
rect 8852 8026 8904 8032
rect 8942 7984 8998 7993
rect 8574 7919 8630 7928
rect 8668 7948 8720 7954
rect 8484 7890 8536 7896
rect 8668 7890 8720 7896
rect 8760 7948 8812 7954
rect 8812 7908 8892 7936
rect 8942 7919 8998 7928
rect 8760 7890 8812 7896
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8496 7290 8524 7890
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8666 7848 8722 7857
rect 8588 7528 8616 7822
rect 8864 7834 8892 7908
rect 8666 7783 8668 7792
rect 8720 7783 8722 7792
rect 8772 7806 8892 7834
rect 8668 7754 8720 7760
rect 8772 7562 8800 7806
rect 8956 7750 8984 7919
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8772 7534 8984 7562
rect 8588 7500 8708 7528
rect 8680 7460 8708 7500
rect 8852 7472 8904 7478
rect 8680 7432 8852 7460
rect 8852 7414 8904 7420
rect 8760 7336 8812 7342
rect 8496 7262 8708 7290
rect 8760 7278 8812 7284
rect 8127 7228 8156 7256
rect 8127 7188 8155 7228
rect 8072 7160 8155 7188
rect 8576 7200 8628 7206
rect 8072 7154 8100 7160
rect 8036 7126 8100 7154
rect 8576 7142 8628 7148
rect 8036 6254 8064 7126
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 8116 6928 8168 6934
rect 8168 6888 8248 6916
rect 8116 6870 8168 6876
rect 8220 6769 8248 6888
rect 8206 6760 8262 6769
rect 8206 6695 8262 6704
rect 8482 6760 8538 6769
rect 8482 6695 8538 6704
rect 8496 6458 8524 6695
rect 8588 6458 8616 7142
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7852 5630 7972 5658
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7208 4282 7236 4694
rect 7484 4282 7512 4762
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7576 4146 7604 4762
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 7116 2990 7144 4014
rect 7760 3058 7788 5510
rect 7852 5370 7880 5630
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7852 3194 7880 5034
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7944 2990 7972 5510
rect 8036 5098 8064 6054
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 3534 8064 5034
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 8588 4146 8616 5510
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8404 3194 8432 3606
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8496 3058 8524 3606
rect 8588 3194 8616 3878
rect 8680 3380 8708 7262
rect 8772 7041 8800 7278
rect 8758 7032 8814 7041
rect 8758 6967 8814 6976
rect 8772 6798 8800 6967
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8864 6390 8892 7414
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5914 8800 6054
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8772 5778 8800 5850
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4010 8800 4490
rect 8864 4282 8892 5034
rect 8956 4826 8984 7534
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 7206 9076 7278
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9140 6984 9168 10406
rect 9232 7410 9260 11018
rect 9600 10962 9628 11154
rect 9678 11112 9734 11121
rect 9678 11047 9680 11056
rect 9732 11047 9734 11056
rect 9680 11018 9732 11024
rect 9600 10934 9720 10962
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 8634 9352 10610
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9416 8378 9444 9386
rect 9508 9058 9536 10406
rect 9600 9178 9628 10474
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9508 9030 9628 9058
rect 9496 8832 9548 8838
rect 9494 8800 9496 8809
rect 9548 8800 9550 8809
rect 9494 8735 9550 8744
rect 9600 8430 9628 9030
rect 9692 8838 9720 10934
rect 9784 10742 9812 12242
rect 9968 12073 9996 12310
rect 10060 12288 10088 12650
rect 10244 12442 10272 13126
rect 10506 13087 10562 13096
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10324 12708 10376 12714
rect 10428 12696 10456 12854
rect 10612 12782 10640 14826
rect 10784 13864 10836 13870
rect 10782 13832 10784 13841
rect 10836 13832 10838 13841
rect 10704 13790 10782 13818
rect 10704 13530 10732 13790
rect 10888 13818 10916 14826
rect 11072 14414 11100 14962
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11164 14074 11192 14418
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11256 13977 11284 14418
rect 11242 13968 11298 13977
rect 11242 13903 11298 13912
rect 10888 13790 11008 13818
rect 10782 13767 10838 13776
rect 10980 13734 11008 13790
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 11244 13728 11296 13734
rect 11348 13705 11376 16102
rect 11610 16079 11666 16088
rect 11716 15706 11744 21354
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21078 12296 21286
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12346 21040 12402 21049
rect 12346 20975 12348 20984
rect 12400 20975 12402 20984
rect 12808 21004 12860 21010
rect 12348 20946 12400 20952
rect 12808 20946 12860 20952
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11794 20632 11850 20641
rect 11794 20567 11796 20576
rect 11848 20567 11850 20576
rect 11796 20538 11848 20544
rect 11992 19922 12020 20810
rect 12394 20800 12446 20806
rect 12394 20742 12446 20748
rect 12059 20700 12367 20709
rect 12059 20698 12065 20700
rect 12121 20698 12145 20700
rect 12201 20698 12225 20700
rect 12281 20698 12305 20700
rect 12361 20698 12367 20700
rect 12121 20646 12123 20698
rect 12303 20646 12305 20698
rect 12059 20644 12065 20646
rect 12121 20644 12145 20646
rect 12201 20644 12225 20646
rect 12281 20644 12305 20646
rect 12361 20644 12367 20646
rect 12059 20635 12367 20644
rect 12406 20584 12434 20742
rect 12268 20556 12434 20584
rect 12268 20330 12296 20556
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12268 20058 12296 20266
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12820 19990 12848 20946
rect 13004 20466 13032 21354
rect 13188 21146 13216 21490
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13280 21321 13308 21354
rect 13372 21350 13400 21655
rect 13648 21622 13676 22086
rect 13726 22063 13782 22072
rect 15200 22024 15252 22030
rect 13726 21992 13782 22001
rect 15200 21966 15252 21972
rect 24584 22024 24636 22030
rect 26884 22024 26936 22030
rect 24584 21966 24636 21972
rect 26054 21992 26110 22001
rect 13726 21927 13782 21936
rect 13636 21616 13688 21622
rect 13542 21584 13598 21593
rect 13636 21558 13688 21564
rect 13542 21519 13598 21528
rect 13556 21486 13584 21519
rect 13544 21480 13596 21486
rect 13464 21440 13544 21468
rect 13360 21344 13412 21350
rect 13266 21312 13322 21321
rect 13360 21286 13412 21292
rect 13266 21247 13322 21256
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13096 20942 13124 21082
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11796 19848 11848 19854
rect 11848 19808 11928 19836
rect 11796 19790 11848 19796
rect 11900 19310 11928 19808
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11808 18358 11836 18566
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11808 18057 11836 18158
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11808 17270 11836 17682
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16697 11836 17070
rect 11900 16726 11928 18770
rect 11992 18086 12020 19858
rect 12268 19802 12296 19858
rect 12532 19848 12584 19854
rect 12268 19774 12480 19802
rect 12532 19790 12584 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12059 19612 12367 19621
rect 12059 19610 12065 19612
rect 12121 19610 12145 19612
rect 12201 19610 12225 19612
rect 12281 19610 12305 19612
rect 12361 19610 12367 19612
rect 12121 19558 12123 19610
rect 12303 19558 12305 19610
rect 12059 19556 12065 19558
rect 12121 19556 12145 19558
rect 12201 19556 12225 19558
rect 12281 19556 12305 19558
rect 12361 19556 12367 19558
rect 12059 19547 12367 19556
rect 12059 18524 12367 18533
rect 12059 18522 12065 18524
rect 12121 18522 12145 18524
rect 12201 18522 12225 18524
rect 12281 18522 12305 18524
rect 12361 18522 12367 18524
rect 12121 18470 12123 18522
rect 12303 18470 12305 18522
rect 12059 18468 12065 18470
rect 12121 18468 12145 18470
rect 12201 18468 12225 18470
rect 12281 18468 12305 18470
rect 12361 18468 12367 18470
rect 12059 18459 12367 18468
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11978 17912 12034 17921
rect 12360 17882 12388 18090
rect 11978 17847 12034 17856
rect 12348 17876 12400 17882
rect 11992 17746 12020 17847
rect 12348 17818 12400 17824
rect 12452 17746 12480 19774
rect 12544 18970 12572 19790
rect 12636 19378 12664 19790
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12544 17898 12572 18906
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18358 12664 18566
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12544 17870 12756 17898
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17320 12020 17478
rect 12059 17436 12367 17445
rect 12059 17434 12065 17436
rect 12121 17434 12145 17436
rect 12201 17434 12225 17436
rect 12281 17434 12305 17436
rect 12361 17434 12367 17436
rect 12121 17382 12123 17434
rect 12303 17382 12305 17434
rect 12059 17380 12065 17382
rect 12121 17380 12145 17382
rect 12201 17380 12225 17382
rect 12281 17380 12305 17382
rect 12361 17380 12367 17382
rect 12059 17371 12367 17380
rect 11992 17292 12112 17320
rect 11978 17096 12034 17105
rect 11978 17031 11980 17040
rect 12032 17031 12034 17040
rect 11980 17002 12032 17008
rect 11978 16960 12034 16969
rect 11978 16895 12034 16904
rect 11888 16720 11940 16726
rect 11794 16688 11850 16697
rect 11888 16662 11940 16668
rect 11794 16623 11850 16632
rect 11992 16250 12020 16895
rect 12084 16658 12112 17292
rect 12532 17264 12584 17270
rect 12452 17224 12532 17252
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16726 12204 16934
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12084 16561 12112 16594
rect 12070 16552 12126 16561
rect 12070 16487 12126 16496
rect 12059 16348 12367 16357
rect 12059 16346 12065 16348
rect 12121 16346 12145 16348
rect 12201 16346 12225 16348
rect 12281 16346 12305 16348
rect 12361 16346 12367 16348
rect 12121 16294 12123 16346
rect 12303 16294 12305 16346
rect 12059 16292 12065 16294
rect 12121 16292 12145 16294
rect 12201 16292 12225 16294
rect 12281 16292 12305 16294
rect 12361 16292 12367 16294
rect 12059 16283 12367 16292
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 14793 11560 15438
rect 11624 15026 11652 15506
rect 11808 15094 11836 15574
rect 11900 15434 11928 16050
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11900 15162 11928 15370
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11886 14920 11942 14929
rect 11886 14855 11942 14864
rect 11900 14822 11928 14855
rect 11888 14816 11940 14822
rect 11518 14784 11574 14793
rect 11888 14758 11940 14764
rect 11518 14719 11574 14728
rect 11992 14550 12020 15370
rect 12059 15260 12367 15269
rect 12059 15258 12065 15260
rect 12121 15258 12145 15260
rect 12201 15258 12225 15260
rect 12281 15258 12305 15260
rect 12361 15258 12367 15260
rect 12121 15206 12123 15258
rect 12303 15206 12305 15258
rect 12059 15204 12065 15206
rect 12121 15204 12145 15206
rect 12201 15204 12225 15206
rect 12281 15204 12305 15206
rect 12361 15204 12367 15206
rect 12059 15195 12367 15204
rect 12452 15094 12480 17224
rect 12532 17206 12584 17212
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12544 15706 12572 17070
rect 12636 16590 12664 17750
rect 12728 17524 12756 17870
rect 12820 17678 12848 19450
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12728 17496 12848 17524
rect 12820 17066 12848 17496
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16590 12756 16934
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12820 16182 12848 17002
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15706 12756 15846
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12440 15088 12492 15094
rect 12728 15076 12756 15506
rect 12808 15088 12860 15094
rect 12728 15048 12808 15076
rect 12440 15030 12492 15036
rect 12808 15030 12860 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12530 14920 12586 14929
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11244 13670 11296 13676
rect 11334 13696 11390 13705
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10376 12668 10456 12696
rect 10324 12650 10376 12656
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10704 12345 10732 13330
rect 10796 12918 10824 13670
rect 11256 13394 11284 13670
rect 11334 13631 11390 13640
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10874 12880 10930 12889
rect 10874 12815 10930 12824
rect 10784 12776 10836 12782
rect 10782 12744 10784 12753
rect 10836 12744 10838 12753
rect 10782 12679 10838 12688
rect 10690 12336 10746 12345
rect 10416 12300 10468 12306
rect 10060 12260 10180 12288
rect 10152 12170 10180 12260
rect 10690 12271 10746 12280
rect 10416 12242 10468 12248
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 9954 12064 10010 12073
rect 9954 11999 10010 12008
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11150 9904 11630
rect 9968 11558 9996 11999
rect 10060 11801 10088 12106
rect 10152 11830 10180 12106
rect 10140 11824 10192 11830
rect 10046 11792 10102 11801
rect 10140 11766 10192 11772
rect 10046 11727 10102 11736
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9784 9586 9812 10678
rect 9968 9926 9996 11222
rect 10060 10810 10088 11727
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10810 10180 11154
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10152 10606 10180 10746
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10152 10130 10180 10367
rect 10244 10266 10272 11630
rect 10322 10976 10378 10985
rect 10322 10911 10378 10920
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 8974 9904 9386
rect 9864 8968 9916 8974
rect 9968 8945 9996 9862
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9864 8910 9916 8916
rect 9954 8936 10010 8945
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8424 9640 8430
rect 9416 8350 9536 8378
rect 9692 8412 9720 8774
rect 9876 8634 9904 8910
rect 9954 8871 10010 8880
rect 9968 8838 9996 8871
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8424 9824 8430
rect 9692 8384 9772 8412
rect 9588 8366 9640 8372
rect 9772 8366 9824 8372
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9324 7954 9352 8230
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7546 9352 7686
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9140 6956 9260 6984
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6322 9076 6734
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9140 5216 9168 6802
rect 9232 6254 9260 6956
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9218 6080 9274 6089
rect 9218 6015 9274 6024
rect 9232 5914 9260 6015
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9220 5228 9272 5234
rect 9140 5188 9220 5216
rect 9220 5170 9272 5176
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9232 4758 9260 5170
rect 9220 4752 9272 4758
rect 9140 4712 9220 4740
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8760 3392 8812 3398
rect 8680 3352 8760 3380
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2650 7512 2790
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 8680 2514 8708 3352
rect 8760 3334 8812 3340
rect 8864 3126 8892 3470
rect 9048 3398 9076 3946
rect 9140 3670 9168 4712
rect 9220 4694 9272 4700
rect 9324 4468 9352 7142
rect 9416 5846 9444 8230
rect 9508 6662 9536 8350
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9508 6118 9536 6394
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9404 5840 9456 5846
rect 9600 5817 9628 8055
rect 9770 7984 9826 7993
rect 9680 7948 9732 7954
rect 9770 7919 9826 7928
rect 9680 7890 9732 7896
rect 9692 6798 9720 7890
rect 9784 7721 9812 7919
rect 9876 7886 9904 8055
rect 9968 7970 9996 8366
rect 10060 8090 10088 9454
rect 10140 9376 10192 9382
rect 10138 9344 10140 9353
rect 10192 9344 10194 9353
rect 10138 9279 10194 9288
rect 10152 8412 10180 9279
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8634 10272 9046
rect 10336 9042 10364 10911
rect 10428 10266 10456 12242
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11778 10548 12174
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10600 11824 10652 11830
rect 10520 11772 10600 11778
rect 10520 11766 10652 11772
rect 10520 11750 10640 11766
rect 10520 10985 10548 11750
rect 10704 11694 10732 12106
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11898 10824 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10888 11694 10916 12815
rect 10980 11898 11008 12922
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12640 11112 12646
rect 11164 12617 11192 12786
rect 11060 12582 11112 12588
rect 11150 12608 11206 12617
rect 11072 12238 11100 12582
rect 11150 12543 11206 12552
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11058 12064 11114 12073
rect 11058 11999 11114 12008
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10506 10976 10562 10985
rect 10506 10911 10562 10920
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10441 10548 10610
rect 10506 10432 10562 10441
rect 10506 10367 10562 10376
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10520 9382 10548 10134
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10336 8634 10364 8978
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10244 8480 10272 8570
rect 10244 8452 10364 8480
rect 10152 8384 10272 8412
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10244 8242 10272 8384
rect 10336 8362 10364 8452
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9968 7942 10088 7970
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7744 9916 7750
rect 9770 7712 9826 7721
rect 9864 7686 9916 7692
rect 9770 7647 9826 7656
rect 9772 7472 9824 7478
rect 9876 7460 9904 7686
rect 9968 7585 9996 7822
rect 9954 7576 10010 7585
rect 9954 7511 10010 7520
rect 9876 7432 9996 7460
rect 9772 7414 9824 7420
rect 9784 6866 9812 7414
rect 9968 7342 9996 7432
rect 10060 7342 10088 7942
rect 10152 7410 10180 8230
rect 10244 8214 10364 8242
rect 10230 8120 10286 8129
rect 10230 8055 10286 8064
rect 10244 7546 10272 8055
rect 10336 7886 10364 8214
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9770 6760 9826 6769
rect 9692 6322 9720 6734
rect 9770 6695 9826 6704
rect 9784 6662 9812 6695
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9876 6458 9904 7278
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9770 6080 9826 6089
rect 9770 6015 9826 6024
rect 9404 5782 9456 5788
rect 9586 5808 9642 5817
rect 9586 5743 9642 5752
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9404 4480 9456 4486
rect 9324 4440 9404 4468
rect 9404 4422 9456 4428
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 3738 9260 4082
rect 9324 3738 9352 4150
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9416 3534 9444 4422
rect 9508 3942 9536 5306
rect 9600 4282 9628 5743
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9784 4010 9812 6015
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9968 3534 9996 7142
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10060 6866 10088 6938
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10152 6662 10180 7346
rect 10232 7336 10284 7342
rect 10230 7304 10232 7313
rect 10284 7304 10286 7313
rect 10230 7239 10286 7248
rect 10428 7002 10456 8871
rect 10520 8498 10548 9114
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10414 6896 10470 6905
rect 10414 6831 10470 6840
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10322 6624 10378 6633
rect 10322 6559 10378 6568
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5778 10272 6258
rect 10336 5953 10364 6559
rect 10322 5944 10378 5953
rect 10322 5879 10378 5888
rect 10336 5778 10364 5879
rect 10428 5778 10456 6831
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10336 5370 10364 5471
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10336 5001 10364 5034
rect 10322 4992 10378 5001
rect 10322 4927 10378 4936
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 9048 2990 9076 3334
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2650 9260 2790
rect 9968 2774 9996 3470
rect 10336 2854 10364 4927
rect 10428 4865 10456 5714
rect 10414 4856 10470 4865
rect 10414 4791 10470 4800
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10428 4282 10456 4626
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10520 4010 10548 8298
rect 10612 7342 10640 11018
rect 10704 9217 10732 11154
rect 10980 11150 11008 11630
rect 11072 11286 11100 11999
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11164 11268 11192 12106
rect 11256 11762 11284 13330
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11348 11694 11376 13330
rect 11532 13326 11560 13874
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11440 12986 11468 13126
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11532 12306 11560 13126
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11624 11898 11652 14214
rect 11716 12714 11744 14418
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 14074 11928 14350
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11992 14074 12020 14282
rect 12059 14172 12367 14181
rect 12059 14170 12065 14172
rect 12121 14170 12145 14172
rect 12201 14170 12225 14172
rect 12281 14170 12305 14172
rect 12361 14170 12367 14172
rect 12121 14118 12123 14170
rect 12303 14118 12305 14170
rect 12059 14116 12065 14118
rect 12121 14116 12145 14118
rect 12201 14116 12225 14118
rect 12281 14116 12305 14118
rect 12361 14116 12367 14118
rect 12059 14107 12367 14116
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11992 13920 12020 14010
rect 11900 13892 12020 13920
rect 11900 13841 11928 13892
rect 11886 13832 11942 13841
rect 11886 13767 11942 13776
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11794 13696 11850 13705
rect 11794 13631 11850 13640
rect 11808 13297 11836 13631
rect 11992 13546 12020 13738
rect 11992 13518 12296 13546
rect 12268 13462 12296 13518
rect 12348 13524 12400 13530
rect 12452 13512 12480 14894
rect 12530 14855 12586 14864
rect 12544 14550 12572 14855
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12820 14482 12848 15030
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12714 14376 12770 14385
rect 12714 14311 12770 14320
rect 12400 13484 12480 13512
rect 12348 13466 12400 13472
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12256 13456 12308 13462
rect 12308 13404 12388 13410
rect 12256 13398 12388 13404
rect 12084 13326 12112 13398
rect 12268 13382 12388 13398
rect 11980 13320 12032 13326
rect 11794 13288 11850 13297
rect 11794 13223 11850 13232
rect 11900 13280 11980 13308
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11716 12306 11744 12650
rect 11900 12442 11928 13280
rect 11980 13262 12032 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12360 13274 12388 13382
rect 12360 13246 12434 13274
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12850 12020 13126
rect 12059 13084 12367 13093
rect 12059 13082 12065 13084
rect 12121 13082 12145 13084
rect 12201 13082 12225 13084
rect 12281 13082 12305 13084
rect 12361 13082 12367 13084
rect 12121 13030 12123 13082
rect 12303 13030 12305 13082
rect 12059 13028 12065 13030
rect 12121 13028 12145 13030
rect 12201 13028 12225 13030
rect 12281 13028 12305 13030
rect 12361 13028 12367 13030
rect 12059 13019 12367 13028
rect 12406 12866 12434 13246
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12360 12838 12434 12866
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11808 11762 11836 12174
rect 11900 11898 11928 12174
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11336 11688 11388 11694
rect 11704 11688 11756 11694
rect 11336 11630 11388 11636
rect 11702 11656 11704 11665
rect 11888 11688 11940 11694
rect 11756 11656 11758 11665
rect 11888 11630 11940 11636
rect 11702 11591 11758 11600
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11244 11280 11296 11286
rect 11164 11240 11244 11268
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 9738 10824 10950
rect 10874 10840 10930 10849
rect 10874 10775 10930 10784
rect 10888 10062 10916 10775
rect 10968 10464 11020 10470
rect 10966 10432 10968 10441
rect 11020 10432 11022 10441
rect 10966 10367 11022 10376
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9897 10916 9998
rect 11072 9926 11100 10066
rect 11164 10062 11192 11240
rect 11244 11222 11296 11228
rect 11336 11280 11388 11286
rect 11532 11257 11560 11494
rect 11900 11286 11928 11630
rect 11888 11280 11940 11286
rect 11336 11222 11388 11228
rect 11518 11248 11574 11257
rect 11348 11150 11376 11222
rect 11428 11212 11480 11218
rect 11888 11222 11940 11228
rect 11518 11183 11520 11192
rect 11428 11154 11480 11160
rect 11572 11183 11574 11192
rect 11704 11212 11756 11218
rect 11520 11154 11572 11160
rect 11704 11154 11756 11160
rect 11336 11144 11388 11150
rect 11334 11112 11336 11121
rect 11388 11112 11390 11121
rect 11256 11070 11334 11098
rect 11256 10130 11284 11070
rect 11334 11047 11390 11056
rect 11334 10704 11390 10713
rect 11334 10639 11390 10648
rect 11348 10538 11376 10639
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11348 10010 11376 10474
rect 11440 10130 11468 11154
rect 11532 10130 11560 11154
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11624 10674 11652 11018
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11612 10056 11664 10062
rect 11348 9982 11468 10010
rect 11612 9998 11664 10004
rect 11060 9920 11112 9926
rect 10874 9888 10930 9897
rect 11060 9862 11112 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 10874 9823 10930 9832
rect 11164 9738 11192 9862
rect 10796 9710 11192 9738
rect 11440 9432 11468 9982
rect 11624 9874 11652 9998
rect 11532 9846 11652 9874
rect 11532 9722 11560 9846
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9586 11652 9658
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11716 9450 11744 11154
rect 11992 11150 12020 12786
rect 12360 12714 12388 12838
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12059 11996 12367 12005
rect 12059 11994 12065 11996
rect 12121 11994 12145 11996
rect 12201 11994 12225 11996
rect 12281 11994 12305 11996
rect 12361 11994 12367 11996
rect 12121 11942 12123 11994
rect 12303 11942 12305 11994
rect 12059 11940 12065 11942
rect 12121 11940 12145 11942
rect 12201 11940 12225 11942
rect 12281 11940 12305 11942
rect 12361 11940 12367 11942
rect 12059 11931 12367 11940
rect 12070 11792 12126 11801
rect 12070 11727 12126 11736
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 11008 11940 11014
rect 11794 10976 11850 10985
rect 12084 10996 12112 11727
rect 12438 11520 12494 11529
rect 12438 11455 12494 11464
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12176 11132 12204 11222
rect 12256 11144 12308 11150
rect 12176 11104 12256 11132
rect 12256 11086 12308 11092
rect 11888 10950 11940 10956
rect 11992 10968 12112 10996
rect 11794 10911 11850 10920
rect 11808 10470 11836 10911
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11900 10266 11928 10950
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11808 9722 11836 10202
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9897 11928 9930
rect 11886 9888 11942 9897
rect 11886 9823 11942 9832
rect 11992 9722 12020 10968
rect 12059 10908 12367 10917
rect 12059 10906 12065 10908
rect 12121 10906 12145 10908
rect 12201 10906 12225 10908
rect 12281 10906 12305 10908
rect 12361 10906 12367 10908
rect 12121 10854 12123 10906
rect 12303 10854 12305 10906
rect 12059 10852 12065 10854
rect 12121 10852 12145 10854
rect 12201 10852 12225 10854
rect 12281 10852 12305 10854
rect 12361 10852 12367 10854
rect 12059 10843 12367 10852
rect 12452 10674 12480 11455
rect 12544 11286 12572 12038
rect 12728 11762 12756 14311
rect 12912 13274 12940 20334
rect 13188 20058 13216 20334
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 13004 19310 13032 19926
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13004 18902 13032 19246
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 13096 18630 13124 19926
rect 13280 19417 13308 20946
rect 13266 19408 13322 19417
rect 13266 19343 13322 19352
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12990 18456 13046 18465
rect 12990 18391 13046 18400
rect 13004 18358 13032 18391
rect 12992 18352 13044 18358
rect 13372 18329 13400 18770
rect 12992 18294 13044 18300
rect 13358 18320 13414 18329
rect 13004 16114 13032 18294
rect 13358 18255 13414 18264
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13358 18184 13414 18193
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13096 16794 13124 17070
rect 13188 16998 13216 17070
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13096 15910 13124 16526
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13188 15570 13216 16390
rect 13176 15564 13228 15570
rect 13280 15552 13308 18158
rect 13464 18170 13492 21440
rect 13544 21422 13596 21428
rect 13648 19514 13676 21558
rect 13740 21146 13768 21927
rect 13818 21856 13874 21865
rect 13818 21791 13874 21800
rect 13832 21690 13860 21791
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 14738 21584 14794 21593
rect 13912 21548 13964 21554
rect 14738 21519 14794 21528
rect 13912 21490 13964 21496
rect 13924 21350 13952 21490
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 13912 21344 13964 21350
rect 14188 21344 14240 21350
rect 13912 21286 13964 21292
rect 14186 21312 14188 21321
rect 14372 21344 14424 21350
rect 14240 21312 14242 21321
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13924 21010 13952 21286
rect 14372 21286 14424 21292
rect 14186 21247 14242 21256
rect 14384 21146 14412 21286
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 20641 13768 20742
rect 13726 20632 13782 20641
rect 13726 20567 13782 20576
rect 13832 20534 13860 20878
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13636 19304 13688 19310
rect 13912 19304 13964 19310
rect 13636 19246 13688 19252
rect 13910 19272 13912 19281
rect 13964 19272 13966 19281
rect 13648 18834 13676 19246
rect 13728 19236 13780 19242
rect 13910 19207 13966 19216
rect 13728 19178 13780 19184
rect 13740 19009 13768 19178
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13726 19000 13782 19009
rect 13726 18935 13782 18944
rect 13740 18834 13768 18935
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13414 18142 13492 18170
rect 13358 18119 13414 18128
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 16658 13400 17614
rect 13464 16998 13492 18022
rect 13542 17776 13598 17785
rect 13542 17711 13544 17720
rect 13596 17711 13598 17720
rect 13636 17740 13688 17746
rect 13544 17682 13596 17688
rect 13636 17682 13688 17688
rect 13648 17202 13676 17682
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13372 16250 13400 16458
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13372 15722 13400 16186
rect 13464 15910 13492 16934
rect 13542 16688 13598 16697
rect 13542 16623 13598 16632
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13372 15694 13492 15722
rect 13360 15564 13412 15570
rect 13280 15524 13360 15552
rect 13176 15506 13228 15512
rect 13360 15506 13412 15512
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 14958 13032 15302
rect 13372 15094 13400 15506
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13004 13938 13032 14894
rect 13464 14414 13492 15694
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 14074 13492 14214
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12912 13258 13032 13274
rect 12912 13252 13044 13258
rect 12912 13246 12992 13252
rect 12992 13194 13044 13200
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13096 12617 13124 12854
rect 13082 12608 13138 12617
rect 13082 12543 13138 12552
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11898 13032 12174
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13096 11830 13124 12038
rect 13084 11824 13136 11830
rect 12990 11792 13046 11801
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12900 11756 12952 11762
rect 12952 11736 12990 11744
rect 13084 11766 13136 11772
rect 12952 11727 13046 11736
rect 12952 11716 13032 11727
rect 12900 11698 12952 11704
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12714 11384 12770 11393
rect 12714 11319 12770 11328
rect 12728 11286 12756 11319
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12440 10668 12492 10674
rect 12360 10628 12440 10656
rect 12162 10296 12218 10305
rect 12162 10231 12218 10240
rect 12176 10033 12204 10231
rect 12360 10130 12388 10628
rect 12440 10610 12492 10616
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12532 10056 12584 10062
rect 12162 10024 12218 10033
rect 12162 9959 12218 9968
rect 12346 10024 12402 10033
rect 12532 9998 12584 10004
rect 12346 9959 12348 9968
rect 12400 9959 12402 9968
rect 12348 9930 12400 9936
rect 12059 9820 12367 9829
rect 12059 9818 12065 9820
rect 12121 9818 12145 9820
rect 12201 9818 12225 9820
rect 12281 9818 12305 9820
rect 12361 9818 12367 9820
rect 12121 9766 12123 9818
rect 12303 9766 12305 9818
rect 12059 9764 12065 9766
rect 12121 9764 12145 9766
rect 12201 9764 12225 9766
rect 12281 9764 12305 9766
rect 12361 9764 12367 9766
rect 12059 9755 12367 9764
rect 11796 9716 11848 9722
rect 11980 9716 12032 9722
rect 11796 9658 11848 9664
rect 11900 9664 11980 9674
rect 11900 9658 12032 9664
rect 11900 9646 12020 9658
rect 12544 9654 12572 9998
rect 12532 9648 12584 9654
rect 11520 9444 11572 9450
rect 11440 9404 11520 9432
rect 11520 9386 11572 9392
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11058 9344 11114 9353
rect 10980 9302 11058 9330
rect 10690 9208 10746 9217
rect 10784 9172 10836 9178
rect 10746 9152 10784 9160
rect 10690 9143 10784 9152
rect 10704 9132 10784 9143
rect 10784 9114 10836 9120
rect 10692 8832 10744 8838
rect 10690 8800 10692 8809
rect 10744 8800 10746 8809
rect 10690 8735 10746 8744
rect 10692 8560 10744 8566
rect 10690 8528 10692 8537
rect 10744 8528 10746 8537
rect 10690 8463 10746 8472
rect 10784 8288 10836 8294
rect 10704 8248 10784 8276
rect 10704 8090 10732 8248
rect 10784 8230 10836 8236
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10980 7954 11008 9302
rect 11058 9279 11114 9288
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8809 11100 8910
rect 11058 8800 11114 8809
rect 11058 8735 11114 8744
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 11072 8090 11100 8599
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7528 10732 7822
rect 10796 7721 10824 7890
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10782 7712 10838 7721
rect 10782 7647 10838 7656
rect 10966 7712 11022 7721
rect 10966 7647 11022 7656
rect 10980 7546 11008 7647
rect 10968 7540 11020 7546
rect 10704 7500 10824 7528
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10704 7342 10732 7375
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10690 6216 10746 6225
rect 10690 6151 10692 6160
rect 10744 6151 10746 6160
rect 10692 6122 10744 6128
rect 10692 5840 10744 5846
rect 10796 5817 10824 7500
rect 10968 7482 11020 7488
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10888 6848 10916 7210
rect 10980 7206 11008 7278
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10968 6860 11020 6866
rect 10888 6820 10968 6848
rect 10968 6802 11020 6808
rect 10692 5782 10744 5788
rect 10782 5808 10838 5817
rect 10598 5128 10654 5137
rect 10598 5063 10654 5072
rect 10612 4146 10640 5063
rect 10704 4826 10732 5782
rect 10782 5743 10838 5752
rect 10876 5772 10928 5778
rect 11072 5760 11100 7754
rect 11164 7546 11192 8978
rect 11256 8401 11284 9114
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11426 8800 11482 8809
rect 11348 8634 11376 8774
rect 11426 8735 11482 8744
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10928 5732 11100 5760
rect 10876 5714 10928 5720
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4690 10824 5510
rect 10980 5302 11008 5578
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10980 4826 11008 5238
rect 11164 5030 11192 7142
rect 11256 7002 11284 7686
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11348 6798 11376 8298
rect 11440 7410 11468 8735
rect 11532 8634 11560 9386
rect 11900 8956 11928 9646
rect 12254 9616 12310 9625
rect 12532 9590 12584 9596
rect 12254 9551 12310 9560
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 9042 12020 9318
rect 12268 9042 12296 9551
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12360 9178 12388 9454
rect 12544 9382 12572 9454
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11716 8928 11928 8956
rect 12084 8945 12112 8978
rect 12070 8936 12126 8945
rect 11716 8650 11744 8928
rect 12070 8871 12126 8880
rect 12059 8732 12367 8741
rect 12059 8730 12065 8732
rect 12121 8730 12145 8732
rect 12201 8730 12225 8732
rect 12281 8730 12305 8732
rect 12361 8730 12367 8732
rect 12121 8678 12123 8730
rect 12303 8678 12305 8730
rect 12059 8676 12065 8678
rect 12121 8676 12145 8678
rect 12201 8676 12225 8678
rect 12281 8676 12305 8678
rect 12361 8676 12367 8678
rect 12059 8667 12367 8676
rect 12636 8650 12664 10134
rect 12716 9920 12768 9926
rect 12820 9897 12848 11630
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12716 9862 12768 9868
rect 12806 9888 12862 9897
rect 12728 9722 12756 9862
rect 12806 9823 12862 9832
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12714 9208 12770 9217
rect 12714 9143 12716 9152
rect 12768 9143 12770 9152
rect 12716 9114 12768 9120
rect 12728 8906 12756 9114
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12820 8820 12848 9318
rect 12912 8974 12940 9522
rect 13004 9382 13032 11290
rect 13188 10810 13216 13806
rect 13464 13462 13492 14010
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13556 13394 13584 16623
rect 13648 16114 13676 17138
rect 13832 17082 13860 19110
rect 13924 18834 13952 19207
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13924 17338 13952 18158
rect 14016 17610 14044 20538
rect 14108 17649 14136 20946
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14200 19718 14228 20334
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14384 19514 14412 20334
rect 14568 19786 14596 21354
rect 14752 21078 14780 21519
rect 15106 21448 15162 21457
rect 15106 21383 15108 21392
rect 15160 21383 15162 21392
rect 15108 21354 15160 21360
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 15212 21010 15240 21966
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15750 21448 15806 21457
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14464 19440 14516 19446
rect 14660 19394 14688 20946
rect 15106 20904 15162 20913
rect 15106 20839 15162 20848
rect 15120 20398 15148 20839
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14752 19514 14780 20334
rect 14844 19990 14872 20334
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14832 19984 14884 19990
rect 14832 19926 14884 19932
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14464 19382 14516 19388
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18630 14412 19246
rect 14188 18624 14240 18630
rect 14372 18624 14424 18630
rect 14188 18566 14240 18572
rect 14278 18592 14334 18601
rect 14094 17640 14150 17649
rect 14004 17604 14056 17610
rect 14094 17575 14150 17584
rect 14004 17546 14056 17552
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13912 17196 13964 17202
rect 14016 17184 14044 17546
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13964 17156 14044 17184
rect 13912 17138 13964 17144
rect 13832 17054 13952 17082
rect 13924 16726 13952 17054
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14108 16454 14136 17478
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13648 12434 13676 14554
rect 13924 14482 13952 14758
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 12714 13860 13670
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13648 12406 13768 12434
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13280 11082 13308 11290
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13464 10985 13492 12310
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 12209 13676 12242
rect 13634 12200 13690 12209
rect 13634 12135 13690 12144
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11830 13584 12038
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 11014 13584 11630
rect 13740 11529 13768 12406
rect 13832 12306 13860 12650
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13726 11520 13782 11529
rect 13726 11455 13782 11464
rect 13726 11384 13782 11393
rect 13832 11370 13860 11562
rect 13782 11342 13860 11370
rect 13924 11354 13952 14418
rect 14016 14090 14044 16118
rect 14200 15706 14228 18566
rect 14372 18566 14424 18572
rect 14278 18527 14334 18536
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14096 14272 14148 14278
rect 14094 14240 14096 14249
rect 14148 14240 14150 14249
rect 14094 14175 14150 14184
rect 14016 14062 14136 14090
rect 14200 14074 14228 15506
rect 14292 14958 14320 18527
rect 14476 18204 14504 19382
rect 14568 19366 14688 19394
rect 14568 18698 14596 19366
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14660 18465 14688 19246
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14646 18456 14702 18465
rect 14646 18391 14702 18400
rect 14648 18216 14700 18222
rect 14476 18176 14648 18204
rect 14648 18158 14700 18164
rect 14646 18048 14702 18057
rect 14646 17983 14702 17992
rect 14660 17377 14688 17983
rect 14646 17368 14702 17377
rect 14752 17338 14780 19178
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14646 17303 14702 17312
rect 14740 17332 14792 17338
rect 14660 17218 14688 17303
rect 14740 17274 14792 17280
rect 14660 17190 14780 17218
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14384 16454 14412 16594
rect 14476 16522 14504 16730
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14462 16416 14518 16425
rect 14462 16351 14518 16360
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14384 15706 14412 15914
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14384 14414 14412 15302
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13258 14044 13806
rect 14108 13734 14136 14062
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14016 12782 14044 13194
rect 14200 12782 14228 13806
rect 14384 13734 14412 14350
rect 14476 13802 14504 16351
rect 14568 16250 14596 17070
rect 14660 16658 14688 17070
rect 14752 16658 14780 17190
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14752 16153 14780 16458
rect 14738 16144 14794 16153
rect 14738 16079 14794 16088
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14844 15994 14872 18566
rect 14936 18222 14964 20198
rect 15028 18630 15056 20334
rect 15106 19816 15162 19825
rect 15106 19751 15162 19760
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18222 15056 18566
rect 15120 18358 15148 19751
rect 15212 19242 15240 20946
rect 15304 20602 15332 21422
rect 15750 21383 15806 21392
rect 15764 21146 15792 21383
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15856 21010 15884 21830
rect 19833 21788 20141 21797
rect 19833 21786 19839 21788
rect 19895 21786 19919 21788
rect 19975 21786 19999 21788
rect 20055 21786 20079 21788
rect 20135 21786 20141 21788
rect 19895 21734 19897 21786
rect 20077 21734 20079 21786
rect 19833 21732 19839 21734
rect 19895 21732 19919 21734
rect 19975 21732 19999 21734
rect 20055 21732 20079 21734
rect 20135 21732 20141 21734
rect 19833 21723 20141 21732
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 15946 21244 16254 21253
rect 15946 21242 15952 21244
rect 16008 21242 16032 21244
rect 16088 21242 16112 21244
rect 16168 21242 16192 21244
rect 16248 21242 16254 21244
rect 16008 21190 16010 21242
rect 16190 21190 16192 21242
rect 15946 21188 15952 21190
rect 16008 21188 16032 21190
rect 16088 21188 16112 21190
rect 16168 21188 16192 21190
rect 16248 21188 16254 21190
rect 15946 21179 16254 21188
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15396 20482 15424 20946
rect 15396 20454 15516 20482
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 19514 15424 20266
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15304 19310 15332 19450
rect 15488 19310 15516 20454
rect 15672 20398 15700 20946
rect 16040 20602 16068 21014
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16316 20602 16344 20946
rect 16396 20936 16448 20942
rect 16500 20913 16528 20946
rect 16396 20878 16448 20884
rect 16486 20904 16542 20913
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 15934 20496 15990 20505
rect 15752 20460 15804 20466
rect 15934 20431 15990 20440
rect 15752 20402 15804 20408
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15580 19922 15608 20334
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15212 19009 15240 19178
rect 15290 19136 15346 19145
rect 15290 19071 15346 19080
rect 15198 19000 15254 19009
rect 15198 18935 15254 18944
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15212 18358 15240 18634
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14936 17048 14964 18158
rect 15212 17542 15240 18294
rect 15304 18068 15332 19071
rect 15488 18306 15516 19246
rect 15580 18766 15608 19246
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15396 18278 15516 18306
rect 15396 18222 15424 18278
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15488 18068 15516 18158
rect 15304 18040 15516 18068
rect 15200 17536 15252 17542
rect 15488 17490 15516 18040
rect 15200 17478 15252 17484
rect 15212 17134 15240 17478
rect 15396 17462 15516 17490
rect 15290 17368 15346 17377
rect 15290 17303 15346 17312
rect 15304 17134 15332 17303
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15016 17060 15068 17066
rect 14936 17020 15016 17048
rect 14936 16658 14964 17020
rect 15016 17002 15068 17008
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14936 16250 14964 16458
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15396 16182 15424 17462
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15292 16040 15344 16046
rect 14922 16008 14978 16017
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13394 14412 13670
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14016 12238 14044 12718
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13726 11319 13782 11328
rect 13544 11008 13596 11014
rect 13450 10976 13506 10985
rect 13544 10950 13596 10956
rect 13450 10911 13506 10920
rect 13556 10810 13584 10950
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13358 10704 13414 10713
rect 13268 10668 13320 10674
rect 13358 10639 13414 10648
rect 13268 10610 13320 10616
rect 13174 10432 13230 10441
rect 13174 10367 13230 10376
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13096 9042 13124 9590
rect 13188 9450 13216 10367
rect 13280 9500 13308 10610
rect 13372 9568 13400 10639
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13556 10169 13584 10474
rect 13634 10432 13690 10441
rect 13634 10367 13690 10376
rect 13542 10160 13598 10169
rect 13542 10095 13598 10104
rect 13648 9722 13676 10367
rect 13740 10062 13768 10746
rect 13832 10198 13860 11342
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14108 11286 14136 12242
rect 14200 12102 14228 12718
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11762 14228 12038
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14292 11286 14320 12582
rect 14476 12345 14504 12650
rect 14462 12336 14518 12345
rect 14462 12271 14518 12280
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14476 10742 14504 11086
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 13820 10192 13872 10198
rect 13872 10140 14136 10146
rect 13820 10134 14136 10140
rect 13832 10130 14136 10134
rect 13832 10124 14148 10130
rect 13832 10118 14096 10124
rect 14096 10066 14148 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9722 13768 9998
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 14004 9580 14056 9586
rect 13372 9540 14004 9568
rect 14004 9522 14056 9528
rect 13280 9472 13584 9500
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12820 8792 12940 8820
rect 11520 8628 11572 8634
rect 11716 8622 11928 8650
rect 11520 8570 11572 8576
rect 11518 8256 11574 8265
rect 11518 8191 11574 8200
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 7002 11468 7142
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11532 6746 11560 8191
rect 11900 7886 11928 8622
rect 12348 8628 12400 8634
rect 12636 8622 12848 8650
rect 12348 8570 12400 8576
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11624 7313 11652 7482
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11610 7304 11666 7313
rect 11610 7239 11666 7248
rect 11624 7002 11652 7239
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11716 6798 11744 7414
rect 11808 7002 11836 7822
rect 11992 7750 12020 8434
rect 12084 8090 12112 8434
rect 12360 8344 12388 8570
rect 12716 8356 12768 8362
rect 12360 8316 12716 8344
rect 12716 8298 12768 8304
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 12059 7644 12367 7653
rect 12059 7642 12065 7644
rect 12121 7642 12145 7644
rect 12201 7642 12225 7644
rect 12281 7642 12305 7644
rect 12361 7642 12367 7644
rect 12121 7590 12123 7642
rect 12303 7590 12305 7642
rect 12059 7588 12065 7590
rect 12121 7588 12145 7590
rect 12201 7588 12225 7590
rect 12281 7588 12305 7590
rect 12361 7588 12367 7590
rect 12059 7579 12367 7588
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 7002 12480 7346
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 11794 6896 11850 6905
rect 11794 6831 11850 6840
rect 11704 6792 11756 6798
rect 11532 6718 11652 6746
rect 11704 6734 11756 6740
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11242 6488 11298 6497
rect 11242 6423 11298 6432
rect 11256 6322 11284 6423
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5710 11376 6122
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 5545 11376 5646
rect 11334 5536 11390 5545
rect 11334 5471 11390 5480
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 10980 4282 11008 4626
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3534 10456 3878
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10428 2922 10456 3470
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10324 2848 10376 2854
rect 10612 2836 10640 4082
rect 11256 3602 11284 4626
rect 11440 3738 11468 6598
rect 11532 6458 11560 6598
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11532 5234 11560 6394
rect 11624 5817 11652 6718
rect 11610 5808 11666 5817
rect 11610 5743 11666 5752
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11532 4146 11560 5170
rect 11808 5098 11836 6831
rect 11992 6458 12020 6938
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12059 6556 12367 6565
rect 12059 6554 12065 6556
rect 12121 6554 12145 6556
rect 12201 6554 12225 6556
rect 12281 6554 12305 6556
rect 12361 6554 12367 6556
rect 12121 6502 12123 6554
rect 12303 6502 12305 6554
rect 12059 6500 12065 6502
rect 12121 6500 12145 6502
rect 12201 6500 12225 6502
rect 12281 6500 12305 6502
rect 12361 6500 12367 6502
rect 12059 6491 12367 6500
rect 12452 6497 12480 6734
rect 12438 6488 12494 6497
rect 11980 6452 12032 6458
rect 12438 6423 12494 6432
rect 11980 6394 12032 6400
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11164 3194 11192 3538
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11440 3126 11468 3334
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11532 3058 11560 4082
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11624 3534 11652 3946
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11808 3126 11836 5034
rect 11900 4826 11928 6326
rect 12059 5468 12367 5477
rect 12059 5466 12065 5468
rect 12121 5466 12145 5468
rect 12201 5466 12225 5468
rect 12281 5466 12305 5468
rect 12361 5466 12367 5468
rect 12121 5414 12123 5466
rect 12303 5414 12305 5466
rect 12059 5412 12065 5414
rect 12121 5412 12145 5414
rect 12201 5412 12225 5414
rect 12281 5412 12305 5414
rect 12361 5412 12367 5414
rect 12059 5403 12367 5412
rect 12544 5234 12572 6802
rect 12636 6662 12664 7822
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12624 6180 12676 6186
rect 12728 6168 12756 8298
rect 12820 8294 12848 8622
rect 12912 8362 12940 8792
rect 13004 8498 13032 8978
rect 13556 8974 13584 9472
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8498 13124 8842
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8022 12848 8230
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12912 7392 12940 8298
rect 13004 8090 13032 8434
rect 13280 8344 13308 8570
rect 13464 8566 13492 8910
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13096 8316 13308 8344
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12820 7364 12940 7392
rect 12820 6905 12848 7364
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12806 6896 12862 6905
rect 12806 6831 12862 6840
rect 12912 6798 12940 7210
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12676 6140 12756 6168
rect 12624 6122 12676 6128
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 12636 4690 12664 6122
rect 12820 5642 12848 6734
rect 12912 5846 12940 6734
rect 13004 6633 13032 7890
rect 12990 6624 13046 6633
rect 12990 6559 13046 6568
rect 12992 6452 13044 6458
rect 13096 6440 13124 8316
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13044 6412 13124 6440
rect 12992 6394 13044 6400
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12912 5166 12940 5782
rect 13004 5778 13032 6394
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12990 5128 13046 5137
rect 12912 5001 12940 5102
rect 12990 5063 13046 5072
rect 12898 4992 12954 5001
rect 12898 4927 12954 4936
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12059 4380 12367 4389
rect 12059 4378 12065 4380
rect 12121 4378 12145 4380
rect 12201 4378 12225 4380
rect 12281 4378 12305 4380
rect 12361 4378 12367 4380
rect 12121 4326 12123 4378
rect 12303 4326 12305 4378
rect 12059 4324 12065 4326
rect 12121 4324 12145 4326
rect 12201 4324 12225 4326
rect 12281 4324 12305 4326
rect 12361 4324 12367 4326
rect 12059 4315 12367 4324
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11992 2990 12020 3674
rect 12636 3670 12664 4626
rect 13004 4554 13032 5063
rect 13096 4554 13124 6190
rect 13188 4554 13216 8026
rect 13372 7954 13400 8366
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7970 13676 8230
rect 13360 7948 13412 7954
rect 13648 7942 13768 7970
rect 13360 7890 13412 7896
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13372 7274 13400 7414
rect 13464 7410 13492 7686
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13464 7002 13492 7346
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13464 6746 13492 6938
rect 13648 6769 13676 6938
rect 13372 6718 13492 6746
rect 13634 6760 13690 6769
rect 13372 6322 13400 6718
rect 13634 6695 13690 6704
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13464 5953 13492 6598
rect 13542 6352 13598 6361
rect 13740 6338 13768 7942
rect 13832 7410 13860 9386
rect 14108 9110 14136 10066
rect 14476 10062 14504 10678
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14568 9625 14596 14486
rect 14660 14482 14688 15506
rect 14752 15473 14780 15982
rect 14844 15966 14922 15994
rect 15292 15982 15344 15988
rect 14922 15943 14978 15952
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14738 15464 14794 15473
rect 14738 15399 14794 15408
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14074 14688 14418
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14752 13954 14780 14758
rect 14844 14550 14872 15506
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14660 13926 14780 13954
rect 14660 12442 14688 13926
rect 14738 13288 14794 13297
rect 14936 13258 14964 15943
rect 15304 15026 15332 15982
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15488 14822 15516 17274
rect 15580 16794 15608 18702
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15672 17785 15700 18158
rect 15658 17776 15714 17785
rect 15658 17711 15714 17720
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15672 15586 15700 17711
rect 15764 17218 15792 20402
rect 15948 20398 15976 20431
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 16408 20210 16436 20878
rect 16486 20839 16542 20848
rect 16592 20534 16620 21626
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 19064 21480 19116 21486
rect 19156 21480 19208 21486
rect 19064 21422 19116 21428
rect 19154 21448 19156 21457
rect 19524 21480 19576 21486
rect 19208 21448 19210 21457
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 18510 21312 18566 21321
rect 16684 21078 16712 21286
rect 18510 21247 18566 21256
rect 18524 21146 18552 21247
rect 19076 21146 19104 21422
rect 19524 21422 19576 21428
rect 19154 21383 19210 21392
rect 18512 21140 18564 21146
rect 19064 21140 19116 21146
rect 18512 21082 18564 21088
rect 18984 21100 19064 21128
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 16580 20528 16632 20534
rect 16632 20476 16804 20482
rect 16580 20470 16804 20476
rect 16592 20454 16804 20470
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16316 20182 16436 20210
rect 15946 20156 16254 20165
rect 15946 20154 15952 20156
rect 16008 20154 16032 20156
rect 16088 20154 16112 20156
rect 16168 20154 16192 20156
rect 16248 20154 16254 20156
rect 16008 20102 16010 20154
rect 16190 20102 16192 20154
rect 15946 20100 15952 20102
rect 16008 20100 16032 20102
rect 16088 20100 16112 20102
rect 16168 20100 16192 20102
rect 16248 20100 16254 20102
rect 15946 20091 16254 20100
rect 15946 19068 16254 19077
rect 15946 19066 15952 19068
rect 16008 19066 16032 19068
rect 16088 19066 16112 19068
rect 16168 19066 16192 19068
rect 16248 19066 16254 19068
rect 16008 19014 16010 19066
rect 16190 19014 16192 19066
rect 15946 19012 15952 19014
rect 16008 19012 16032 19014
rect 16088 19012 16112 19014
rect 16168 19012 16192 19014
rect 16248 19012 16254 19014
rect 15946 19003 16254 19012
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15856 18306 15884 18362
rect 15856 18290 16160 18306
rect 15856 18284 16172 18290
rect 15856 18278 16120 18284
rect 15856 17338 15884 18278
rect 16120 18226 16172 18232
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 18086 16068 18158
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15946 17980 16254 17989
rect 15946 17978 15952 17980
rect 16008 17978 16032 17980
rect 16088 17978 16112 17980
rect 16168 17978 16192 17980
rect 16248 17978 16254 17980
rect 16008 17926 16010 17978
rect 16190 17926 16192 17978
rect 15946 17924 15952 17926
rect 16008 17924 16032 17926
rect 16088 17924 16112 17926
rect 16168 17924 16192 17926
rect 16248 17924 16254 17926
rect 15946 17915 16254 17924
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15764 17190 15884 17218
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16114 15792 17070
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15750 15600 15806 15609
rect 15672 15558 15750 15586
rect 15750 15535 15806 15544
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 14958 15792 15302
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15476 14612 15528 14618
rect 15672 14600 15700 14894
rect 15672 14572 15792 14600
rect 15476 14554 15528 14560
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15028 13870 15056 14418
rect 15396 13938 15424 14486
rect 15488 14482 15516 14554
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14074 15700 14418
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13394 15056 13806
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14738 13223 14794 13232
rect 14924 13252 14976 13258
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14752 12170 14780 13223
rect 14924 13194 14976 13200
rect 15120 12986 15148 13330
rect 15212 12986 15240 13738
rect 15396 13394 15424 13874
rect 15672 13870 15700 14010
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15488 13394 15516 13738
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15200 12776 15252 12782
rect 15120 12736 15200 12764
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14936 11898 14964 12650
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15028 12073 15056 12310
rect 15014 12064 15070 12073
rect 15014 11999 15070 12008
rect 15014 11928 15070 11937
rect 14924 11892 14976 11898
rect 15014 11863 15070 11872
rect 14924 11834 14976 11840
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14660 10266 14688 11018
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14752 10062 14780 10610
rect 14844 10606 14872 11154
rect 14924 11144 14976 11150
rect 14922 11112 14924 11121
rect 14976 11112 14978 11121
rect 15028 11082 15056 11863
rect 14922 11047 14978 11056
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15120 10810 15148 12736
rect 15200 12718 15252 12724
rect 15476 12708 15528 12714
rect 15304 12668 15476 12696
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12481 15240 12582
rect 15198 12472 15254 12481
rect 15198 12407 15254 12416
rect 15304 12306 15332 12668
rect 15476 12650 15528 12656
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15304 11694 15332 12242
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 10266 14872 10542
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10305 14964 10406
rect 14922 10296 14978 10305
rect 14832 10260 14884 10266
rect 15212 10266 15240 11018
rect 15396 10849 15424 11494
rect 15488 11354 15516 12378
rect 15580 11898 15608 13398
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15580 11354 15608 11562
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15672 11257 15700 13670
rect 15764 13258 15792 14572
rect 15856 13394 15884 17190
rect 16224 17082 16252 17614
rect 16316 17202 16344 20182
rect 16500 20058 16528 20334
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16488 20052 16540 20058
rect 16408 20012 16488 20040
rect 16408 19718 16436 20012
rect 16488 19994 16540 20000
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16500 19514 16528 19790
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16592 19417 16620 20198
rect 16578 19408 16634 19417
rect 16396 19372 16448 19378
rect 16448 19332 16528 19360
rect 16578 19343 16634 19352
rect 16396 19314 16448 19320
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16408 18329 16436 19178
rect 16394 18320 16450 18329
rect 16500 18306 16528 19332
rect 16580 19304 16632 19310
rect 16632 19264 16712 19292
rect 16580 19246 16632 19252
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16592 18766 16620 19110
rect 16684 19009 16712 19264
rect 16776 19145 16804 20454
rect 17328 20398 17356 20742
rect 17972 20602 18000 21014
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18248 20602 18276 20946
rect 17960 20596 18012 20602
rect 18236 20596 18288 20602
rect 18012 20556 18092 20584
rect 17960 20538 18012 20544
rect 16948 20392 17000 20398
rect 16946 20360 16948 20369
rect 17040 20392 17092 20398
rect 17000 20360 17002 20369
rect 17040 20334 17092 20340
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 16946 20295 17002 20304
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16960 19310 16988 20198
rect 17052 19922 17080 20334
rect 17328 19990 17356 20334
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16762 19136 16818 19145
rect 16762 19071 16818 19080
rect 16670 19000 16726 19009
rect 16670 18935 16726 18944
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16684 18465 16712 18838
rect 16776 18578 16804 19071
rect 16868 18698 16896 19246
rect 17052 18850 17080 19858
rect 17222 19544 17278 19553
rect 17222 19479 17278 19488
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17144 18970 17172 19314
rect 17236 19310 17264 19479
rect 17224 19304 17276 19310
rect 17222 19272 17224 19281
rect 17276 19272 17278 19281
rect 17222 19207 17278 19216
rect 17222 19000 17278 19009
rect 17132 18964 17184 18970
rect 17222 18935 17224 18944
rect 17132 18906 17184 18912
rect 17276 18935 17278 18944
rect 17224 18906 17276 18912
rect 16948 18828 17000 18834
rect 17052 18822 17172 18850
rect 16948 18770 17000 18776
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16854 18592 16910 18601
rect 16776 18550 16854 18578
rect 16960 18578 16988 18770
rect 16910 18550 16988 18578
rect 16854 18527 16910 18536
rect 16670 18456 16726 18465
rect 16670 18391 16726 18400
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16500 18278 16712 18306
rect 16394 18255 16450 18264
rect 16408 17660 16436 18255
rect 16488 18080 16540 18086
rect 16580 18080 16632 18086
rect 16488 18022 16540 18028
rect 16578 18048 16580 18057
rect 16632 18048 16634 18057
rect 16500 17762 16528 18022
rect 16578 17983 16634 17992
rect 16578 17912 16634 17921
rect 16578 17847 16580 17856
rect 16632 17847 16634 17856
rect 16580 17818 16632 17824
rect 16500 17734 16620 17762
rect 16684 17746 16712 18278
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16776 17785 16804 18090
rect 16762 17776 16818 17785
rect 16408 17632 16528 17660
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16396 17128 16448 17134
rect 16224 17054 16344 17082
rect 16396 17070 16448 17076
rect 15946 16892 16254 16901
rect 15946 16890 15952 16892
rect 16008 16890 16032 16892
rect 16088 16890 16112 16892
rect 16168 16890 16192 16892
rect 16248 16890 16254 16892
rect 16008 16838 16010 16890
rect 16190 16838 16192 16890
rect 15946 16836 15952 16838
rect 16008 16836 16032 16838
rect 16088 16836 16112 16838
rect 16168 16836 16192 16838
rect 16248 16836 16254 16838
rect 15946 16827 16254 16836
rect 16316 16522 16344 17054
rect 16408 16658 16436 17070
rect 16500 17066 16528 17632
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16500 16538 16528 16759
rect 16592 16726 16620 17734
rect 16672 17740 16724 17746
rect 16762 17711 16818 17720
rect 16672 17682 16724 17688
rect 16868 17660 16896 18158
rect 16960 17882 16988 18158
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16868 17632 16988 17660
rect 16960 17338 16988 17632
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17052 17184 17080 18362
rect 17144 18204 17172 18822
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17236 18426 17264 18770
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17224 18216 17276 18222
rect 17144 18176 17224 18204
rect 17224 18158 17276 18164
rect 17224 18080 17276 18086
rect 17144 18040 17224 18068
rect 17144 17377 17172 18040
rect 17224 18022 17276 18028
rect 17328 17746 17356 19926
rect 17512 19922 17540 20198
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17130 17368 17186 17377
rect 17130 17303 17186 17312
rect 16960 17156 17080 17184
rect 17222 17232 17278 17241
rect 17222 17167 17278 17176
rect 16960 16810 16988 17156
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16960 16782 17080 16810
rect 16580 16720 16632 16726
rect 16578 16688 16580 16697
rect 16632 16688 16634 16697
rect 16578 16623 16634 16632
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16408 16510 16528 16538
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16946 16552 17002 16561
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 15946 15804 16254 15813
rect 15946 15802 15952 15804
rect 16008 15802 16032 15804
rect 16088 15802 16112 15804
rect 16168 15802 16192 15804
rect 16248 15802 16254 15804
rect 16008 15750 16010 15802
rect 16190 15750 16192 15802
rect 15946 15748 15952 15750
rect 16008 15748 16032 15750
rect 16088 15748 16112 15750
rect 16168 15748 16192 15750
rect 16248 15748 16254 15750
rect 15946 15739 16254 15748
rect 16316 15706 16344 16186
rect 16408 16182 16436 16510
rect 16684 16425 16712 16526
rect 16764 16448 16816 16454
rect 16670 16416 16726 16425
rect 16764 16390 16816 16396
rect 16670 16351 16726 16360
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16040 14958 16068 15506
rect 16224 15162 16252 15574
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 15946 14716 16254 14725
rect 15946 14714 15952 14716
rect 16008 14714 16032 14716
rect 16088 14714 16112 14716
rect 16168 14714 16192 14716
rect 16248 14714 16254 14716
rect 16008 14662 16010 14714
rect 16190 14662 16192 14714
rect 15946 14660 15952 14662
rect 16008 14660 16032 14662
rect 16088 14660 16112 14662
rect 16168 14660 16192 14662
rect 16248 14660 16254 14662
rect 15946 14651 16254 14660
rect 16316 14618 16344 14894
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16408 14278 16436 16118
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16500 15570 16528 15642
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 14618 16620 15506
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16684 14414 16712 16351
rect 16776 16182 16804 16390
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16776 15162 16804 15370
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 14414 16804 14894
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16500 13841 16528 14282
rect 16486 13832 16542 13841
rect 16486 13767 16542 13776
rect 15946 13628 16254 13637
rect 15946 13626 15952 13628
rect 16008 13626 16032 13628
rect 16088 13626 16112 13628
rect 16168 13626 16192 13628
rect 16248 13626 16254 13628
rect 16008 13574 16010 13626
rect 16190 13574 16192 13626
rect 15946 13572 15952 13574
rect 16008 13572 16032 13574
rect 16088 13572 16112 13574
rect 16168 13572 16192 13574
rect 16248 13572 16254 13574
rect 15946 13563 16254 13572
rect 16592 13394 16620 14350
rect 16684 14074 16712 14350
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16868 13716 16896 16526
rect 16946 16487 17002 16496
rect 16960 16454 16988 16487
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16960 15337 16988 15574
rect 16946 15328 17002 15337
rect 16946 15263 17002 15272
rect 17052 15094 17080 16782
rect 17144 16454 17172 17070
rect 17236 16998 17264 17167
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17130 15736 17186 15745
rect 17130 15671 17186 15680
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16946 14920 17002 14929
rect 16946 14855 17002 14864
rect 16960 13870 16988 14855
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 17052 14260 17080 14486
rect 17144 14414 17172 15671
rect 17236 14958 17264 16594
rect 17328 16250 17356 17682
rect 17420 17202 17448 19654
rect 17512 19446 17540 19722
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17512 18426 17540 19246
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17512 17746 17540 18362
rect 17604 18086 17632 20334
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17880 20233 17908 20266
rect 17866 20224 17922 20233
rect 17866 20159 17922 20168
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17696 19310 17724 19994
rect 17880 19854 17908 20159
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17868 19848 17920 19854
rect 17788 19808 17868 19836
rect 17788 19689 17816 19808
rect 17868 19790 17920 19796
rect 17868 19712 17920 19718
rect 17774 19680 17830 19689
rect 17868 19654 17920 19660
rect 17774 19615 17830 19624
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17696 18970 17724 19110
rect 17788 18970 17816 19178
rect 17880 19174 17908 19654
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17696 18154 17724 18634
rect 17776 18624 17828 18630
rect 17880 18612 17908 19110
rect 17972 18834 18000 19858
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17828 18584 17908 18612
rect 17776 18566 17828 18572
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17420 16538 17448 17002
rect 17512 16833 17540 17546
rect 17696 17490 17724 18090
rect 17788 17882 17816 18566
rect 17868 18216 17920 18222
rect 17866 18184 17868 18193
rect 17920 18184 17922 18193
rect 17866 18119 17922 18128
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17774 17776 17830 17785
rect 17880 17746 17908 18119
rect 17774 17711 17830 17720
rect 17868 17740 17920 17746
rect 17788 17592 17816 17711
rect 17868 17682 17920 17688
rect 17788 17564 17908 17592
rect 17696 17462 17816 17490
rect 17684 17332 17736 17338
rect 17604 17292 17684 17320
rect 17498 16824 17554 16833
rect 17498 16759 17554 16768
rect 17512 16658 17540 16759
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17420 16510 17540 16538
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17420 16182 17448 16390
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17512 16130 17540 16510
rect 17604 16504 17632 17292
rect 17684 17274 17736 17280
rect 17604 16476 17724 16504
rect 17512 16102 17632 16130
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17328 14822 17356 15982
rect 17420 15881 17448 15982
rect 17406 15872 17462 15881
rect 17406 15807 17462 15816
rect 17406 15736 17462 15745
rect 17512 15706 17540 15982
rect 17604 15910 17632 16102
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15706 17632 15846
rect 17406 15671 17462 15680
rect 17500 15700 17552 15706
rect 17420 15638 17448 15671
rect 17500 15642 17552 15648
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17604 15162 17632 15302
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17236 14618 17264 14758
rect 17420 14618 17448 14826
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17236 14521 17264 14554
rect 17222 14512 17278 14521
rect 17222 14447 17278 14456
rect 17132 14408 17184 14414
rect 17316 14408 17368 14414
rect 17184 14368 17316 14396
rect 17132 14350 17184 14356
rect 17316 14350 17368 14356
rect 17132 14272 17184 14278
rect 17052 14232 17132 14260
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16868 13688 16988 13716
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16212 13320 16264 13326
rect 16764 13320 16816 13326
rect 16264 13268 16620 13274
rect 16212 13262 16620 13268
rect 16764 13262 16816 13268
rect 15752 13252 15804 13258
rect 16224 13246 16620 13262
rect 15752 13194 15804 13200
rect 15764 12918 15792 13194
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15844 12640 15896 12646
rect 16408 12594 16436 12922
rect 16486 12608 16542 12617
rect 15844 12582 15896 12588
rect 15750 12472 15806 12481
rect 15750 12407 15806 12416
rect 15856 12424 15884 12582
rect 16316 12566 16486 12594
rect 15946 12540 16254 12549
rect 15946 12538 15952 12540
rect 16008 12538 16032 12540
rect 16088 12538 16112 12540
rect 16168 12538 16192 12540
rect 16248 12538 16254 12540
rect 16008 12486 16010 12538
rect 16190 12486 16192 12538
rect 15946 12484 15952 12486
rect 16008 12484 16032 12486
rect 16088 12484 16112 12486
rect 16168 12484 16192 12486
rect 16248 12484 16254 12486
rect 15946 12475 16254 12484
rect 16212 12436 16264 12442
rect 15764 12374 15792 12407
rect 15856 12396 16212 12424
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15750 12200 15806 12209
rect 15750 12135 15806 12144
rect 15764 12102 15792 12135
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15856 11558 15884 12396
rect 16212 12378 16264 12384
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15948 11558 15976 12242
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 11694 16160 12106
rect 16224 11830 16252 12242
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15844 11552 15896 11558
rect 15750 11520 15806 11529
rect 15844 11494 15896 11500
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15750 11455 15806 11464
rect 15474 11248 15530 11257
rect 15658 11248 15714 11257
rect 15530 11218 15608 11234
rect 15530 11212 15620 11218
rect 15530 11206 15568 11212
rect 15474 11183 15530 11192
rect 15658 11183 15714 11192
rect 15568 11154 15620 11160
rect 15382 10840 15438 10849
rect 15382 10775 15438 10784
rect 15672 10538 15700 11183
rect 15764 10690 15792 11455
rect 15856 11014 15884 11494
rect 15946 11452 16254 11461
rect 15946 11450 15952 11452
rect 16008 11450 16032 11452
rect 16088 11450 16112 11452
rect 16168 11450 16192 11452
rect 16248 11450 16254 11452
rect 16008 11398 16010 11450
rect 16190 11398 16192 11450
rect 15946 11396 15952 11398
rect 16008 11396 16032 11398
rect 16088 11396 16112 11398
rect 16168 11396 16192 11398
rect 16248 11396 16254 11398
rect 15946 11387 16254 11396
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 16132 10713 16160 11018
rect 16118 10704 16174 10713
rect 15764 10662 15884 10690
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 14922 10231 14978 10240
rect 15200 10260 15252 10266
rect 14832 10202 14884 10208
rect 15200 10202 15252 10208
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 14740 10056 14792 10062
rect 14738 10024 14740 10033
rect 14792 10024 14794 10033
rect 14738 9959 14794 9968
rect 15580 9926 15608 10066
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15568 9648 15620 9654
rect 14554 9616 14610 9625
rect 15568 9590 15620 9596
rect 14554 9551 14610 9560
rect 15384 9580 15436 9586
rect 14186 9344 14242 9353
rect 14186 9279 14242 9288
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8294 13952 8910
rect 14200 8362 14228 9279
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 7834 14044 8230
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 13924 7806 14044 7834
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13598 6310 13768 6338
rect 13542 6287 13598 6296
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13450 5944 13506 5953
rect 13450 5879 13506 5888
rect 13464 5710 13492 5879
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 5296 13412 5302
rect 13358 5264 13360 5273
rect 13412 5264 13414 5273
rect 13358 5199 13414 5208
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13004 4146 13032 4490
rect 13556 4146 13584 6190
rect 13636 6112 13688 6118
rect 13924 6066 13952 7806
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 6254 14044 7686
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6458 14136 7210
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14200 6662 14228 6870
rect 14188 6656 14240 6662
rect 14280 6656 14332 6662
rect 14188 6598 14240 6604
rect 14278 6624 14280 6633
rect 14332 6624 14334 6633
rect 14278 6559 14334 6568
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13636 6054 13688 6060
rect 13648 5914 13676 6054
rect 13832 6038 13952 6066
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3942 13584 4082
rect 13832 4010 13860 6038
rect 14200 5302 14228 6258
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14292 5574 14320 6190
rect 14384 5778 14412 6394
rect 14476 6089 14504 7346
rect 14568 6798 14596 9551
rect 15384 9522 15436 9528
rect 15396 9382 15424 9522
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9217 15424 9318
rect 15382 9208 15438 9217
rect 15382 9143 15438 9152
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15120 8514 15148 8570
rect 14844 8486 15148 8514
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 14844 8430 14872 8486
rect 14832 8424 14884 8430
rect 15212 8378 15240 8502
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14832 8366 14884 8372
rect 15120 8350 15240 8378
rect 15120 7206 15148 8350
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7342 15240 8230
rect 15304 7886 15332 8434
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 14556 6792 14608 6798
rect 14924 6792 14976 6798
rect 14556 6734 14608 6740
rect 14738 6760 14794 6769
rect 14738 6695 14794 6704
rect 14844 6752 14924 6780
rect 14752 6458 14780 6695
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14462 6080 14518 6089
rect 14462 6015 14518 6024
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4752 13964 4758
rect 13910 4720 13912 4729
rect 13964 4720 13966 4729
rect 13910 4655 13966 4664
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13832 3670 13860 3946
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 12059 3292 12367 3301
rect 12059 3290 12065 3292
rect 12121 3290 12145 3292
rect 12201 3290 12225 3292
rect 12281 3290 12305 3292
rect 12361 3290 12367 3292
rect 12121 3238 12123 3290
rect 12303 3238 12305 3290
rect 12059 3236 12065 3238
rect 12121 3236 12145 3238
rect 12201 3236 12225 3238
rect 12281 3236 12305 3238
rect 12361 3236 12367 3238
rect 12059 3227 12367 3236
rect 13924 3058 13952 4655
rect 14016 4622 14044 4966
rect 14108 4826 14136 5102
rect 14200 5001 14228 5238
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14186 4992 14242 5001
rect 14186 4927 14242 4936
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 4214 14044 4558
rect 14292 4282 14320 5102
rect 14476 4690 14504 5714
rect 14568 5574 14596 6258
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14660 4690 14688 5238
rect 14752 4826 14780 5714
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14016 3670 14044 4150
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14016 2990 14044 3606
rect 14476 3602 14504 3878
rect 14844 3738 14872 6752
rect 14924 6734 14976 6740
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15028 6322 15056 6666
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15120 6254 15148 6870
rect 15212 6662 15240 7278
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15396 6186 15424 8910
rect 15488 8362 15516 9454
rect 15580 9110 15608 9590
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 8090 15608 8230
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15580 7478 15608 8026
rect 15672 8022 15700 10474
rect 15764 10198 15792 10474
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15856 9704 15884 10662
rect 16118 10639 16174 10648
rect 15946 10364 16254 10373
rect 15946 10362 15952 10364
rect 16008 10362 16032 10364
rect 16088 10362 16112 10364
rect 16168 10362 16192 10364
rect 16248 10362 16254 10364
rect 16008 10310 16010 10362
rect 16190 10310 16192 10362
rect 15946 10308 15952 10310
rect 16008 10308 16032 10310
rect 16088 10308 16112 10310
rect 16168 10308 16192 10310
rect 16248 10308 16254 10310
rect 15946 10299 16254 10308
rect 16316 10198 16344 12566
rect 16486 12543 16542 12552
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16408 12170 16436 12242
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16408 11218 16436 11319
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10198 16436 10406
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 15764 9676 15884 9704
rect 15764 8786 15792 9676
rect 16408 9654 16436 9998
rect 16396 9648 16448 9654
rect 15842 9616 15898 9625
rect 16396 9590 16448 9596
rect 15842 9551 15844 9560
rect 15896 9551 15898 9560
rect 15844 9522 15896 9528
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 15946 9276 16254 9285
rect 15946 9274 15952 9276
rect 16008 9274 16032 9276
rect 16088 9274 16112 9276
rect 16168 9274 16192 9276
rect 16248 9274 16254 9276
rect 16008 9222 16010 9274
rect 16190 9222 16192 9274
rect 15946 9220 15952 9222
rect 16008 9220 16032 9222
rect 16088 9220 16112 9222
rect 16168 9220 16192 9222
rect 16248 9220 16254 9222
rect 15946 9211 16254 9220
rect 16316 9042 16344 9386
rect 16408 9178 16436 9386
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 15764 8758 15884 8786
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15764 6458 15792 8570
rect 15856 7970 15884 8758
rect 15946 8188 16254 8197
rect 15946 8186 15952 8188
rect 16008 8186 16032 8188
rect 16088 8186 16112 8188
rect 16168 8186 16192 8188
rect 16248 8186 16254 8188
rect 16008 8134 16010 8186
rect 16190 8134 16192 8186
rect 15946 8132 15952 8134
rect 16008 8132 16032 8134
rect 16088 8132 16112 8134
rect 16168 8132 16192 8134
rect 16248 8132 16254 8134
rect 15946 8123 16254 8132
rect 15856 7942 15976 7970
rect 15948 7410 15976 7942
rect 16316 7410 16344 8978
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 8673 16436 8774
rect 16394 8664 16450 8673
rect 16500 8634 16528 11494
rect 16592 11286 16620 13246
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12866 16712 13194
rect 16776 12986 16804 13262
rect 16868 13025 16896 13398
rect 16960 13297 16988 13688
rect 17052 13462 17080 14232
rect 17132 14214 17184 14220
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16946 13288 17002 13297
rect 16946 13223 17002 13232
rect 16854 13016 16910 13025
rect 16764 12980 16816 12986
rect 16854 12951 16910 12960
rect 16764 12922 16816 12928
rect 16684 12838 16804 12866
rect 16776 12646 16804 12838
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12442 16804 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16856 12300 16908 12306
rect 16960 12288 16988 12378
rect 17052 12374 17080 13398
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16908 12260 16988 12288
rect 16856 12242 16908 12248
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16670 12064 16726 12073
rect 16670 11999 16726 12008
rect 16684 11762 16712 11999
rect 16868 11762 16896 12106
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16580 11144 16632 11150
rect 16684 11132 16712 11698
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16632 11121 16712 11132
rect 16632 11112 16726 11121
rect 16632 11104 16670 11112
rect 16580 11086 16632 11092
rect 16670 11047 16726 11056
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 9518 16620 10406
rect 16776 9654 16804 11630
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 10266 16896 11562
rect 16960 11558 16988 12260
rect 17144 11801 17172 13874
rect 17420 13394 17448 14554
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 13161 17448 13330
rect 17604 13326 17632 14010
rect 17696 13870 17724 16476
rect 17788 16046 17816 17462
rect 17880 17338 17908 17564
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17972 17134 18000 18770
rect 18064 17218 18092 20556
rect 18236 20538 18288 20544
rect 18340 20262 18368 20946
rect 18880 20936 18932 20942
rect 18984 20924 19012 21100
rect 19064 21082 19116 21088
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19260 21049 19288 21082
rect 19432 21072 19484 21078
rect 19246 21040 19302 21049
rect 19432 21014 19484 21020
rect 19246 20975 19302 20984
rect 18932 20896 19012 20924
rect 19064 20936 19116 20942
rect 18880 20878 18932 20884
rect 19064 20878 19116 20884
rect 18788 20800 18840 20806
rect 18418 20768 18474 20777
rect 18788 20742 18840 20748
rect 18418 20703 18474 20712
rect 18432 20534 18460 20703
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18524 20058 18552 20402
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18420 19984 18472 19990
rect 18616 19938 18644 20470
rect 18420 19926 18472 19932
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 18902 18184 19790
rect 18432 19378 18460 19926
rect 18524 19910 18644 19938
rect 18694 19952 18750 19961
rect 18524 19718 18552 19910
rect 18694 19887 18750 19896
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18602 19680 18658 19689
rect 18602 19615 18658 19624
rect 18616 19446 18644 19615
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18156 17377 18184 18838
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18142 17368 18198 17377
rect 18142 17303 18198 17312
rect 18064 17190 18184 17218
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17880 16425 17908 16662
rect 17972 16454 18000 16934
rect 18064 16522 18092 17070
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17960 16448 18012 16454
rect 17866 16416 17922 16425
rect 17960 16390 18012 16396
rect 17866 16351 17922 16360
rect 18156 16182 18184 17190
rect 17960 16176 18012 16182
rect 17880 16136 17960 16164
rect 17880 16130 17908 16136
rect 17864 16102 17908 16130
rect 17960 16118 18012 16124
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17864 15960 17892 16102
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17864 15932 17908 15960
rect 17774 15736 17830 15745
rect 17774 15671 17830 15680
rect 17788 15434 17816 15671
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17880 15366 17908 15932
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17972 15194 18000 15982
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17788 15166 18000 15194
rect 17788 14249 17816 15166
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17774 14240 17830 14249
rect 17774 14175 17830 14184
rect 17774 14104 17830 14113
rect 17774 14039 17776 14048
rect 17828 14039 17830 14048
rect 17776 14010 17828 14016
rect 17880 14006 17908 15030
rect 18064 14822 18092 15438
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14618 18092 14758
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17774 13696 17830 13705
rect 17830 13654 17908 13682
rect 17774 13631 17830 13640
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17880 13190 17908 13654
rect 17972 13394 18000 14282
rect 18064 13462 18092 14418
rect 18248 14414 18276 17546
rect 18340 17338 18368 18906
rect 18432 18766 18460 18906
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18432 17218 18460 18702
rect 18524 18086 18552 18799
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18524 17649 18552 17818
rect 18510 17640 18566 17649
rect 18510 17575 18566 17584
rect 18340 17190 18460 17218
rect 18340 15978 18368 17190
rect 18512 16992 18564 16998
rect 18418 16960 18474 16969
rect 18512 16934 18564 16940
rect 18418 16895 18474 16904
rect 18432 16794 18460 16895
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18340 15366 18368 15642
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18432 15162 18460 16730
rect 18524 15706 18552 16934
rect 18616 16590 18644 19178
rect 18708 18222 18736 19887
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18708 17882 18736 18158
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18800 17066 18828 20742
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18892 19922 18920 19994
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18892 19689 18920 19858
rect 18878 19680 18934 19689
rect 18878 19615 18934 19624
rect 19076 19514 19104 20878
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19168 19990 19196 20402
rect 19352 20262 19380 20810
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19246 20088 19302 20097
rect 19246 20023 19302 20032
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19260 19836 19288 20023
rect 19352 19922 19380 20198
rect 19444 19922 19472 21014
rect 19536 20777 19564 21422
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19522 20768 19578 20777
rect 19522 20703 19578 20712
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19168 19808 19288 19836
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18892 17746 18920 19450
rect 19076 19310 19104 19450
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 18984 18816 19012 19246
rect 19168 18834 19196 19808
rect 19352 19530 19380 19858
rect 19260 19502 19380 19530
rect 19064 18828 19116 18834
rect 18984 18788 19064 18816
rect 19064 18770 19116 18776
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19076 18306 19104 18770
rect 19154 18320 19210 18329
rect 18972 18284 19024 18290
rect 19076 18278 19154 18306
rect 19154 18255 19210 18264
rect 18972 18226 19024 18232
rect 18984 18057 19012 18226
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18970 18048 19026 18057
rect 18970 17983 19026 17992
rect 18970 17912 19026 17921
rect 18970 17847 19026 17856
rect 18984 17814 19012 17847
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16046 18644 16390
rect 18708 16182 18736 17002
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18524 15484 18552 15642
rect 18604 15496 18656 15502
rect 18524 15456 18604 15484
rect 18604 15438 18656 15444
rect 18708 15194 18736 16118
rect 18800 15484 18828 17002
rect 18892 16969 18920 17682
rect 18878 16960 18934 16969
rect 18878 16895 18934 16904
rect 18984 16250 19012 17750
rect 19076 17134 19104 18158
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19168 17746 19196 18022
rect 19260 17898 19288 19502
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19444 19174 19472 19382
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19536 18970 19564 19858
rect 19628 19446 19656 21286
rect 20272 21010 20300 21558
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 19833 20700 20141 20709
rect 19833 20698 19839 20700
rect 19895 20698 19919 20700
rect 19975 20698 19999 20700
rect 20055 20698 20079 20700
rect 20135 20698 20141 20700
rect 19895 20646 19897 20698
rect 20077 20646 20079 20698
rect 19833 20644 19839 20646
rect 19895 20644 19919 20646
rect 19975 20644 19999 20646
rect 20055 20644 20079 20646
rect 20135 20644 20141 20646
rect 19833 20635 20141 20644
rect 20272 20534 20300 20946
rect 19800 20528 19852 20534
rect 19800 20470 19852 20476
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19720 19961 19748 20334
rect 19706 19952 19762 19961
rect 19706 19887 19762 19896
rect 19812 19786 19840 20470
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20272 20262 20300 20334
rect 19984 20256 20036 20262
rect 20260 20256 20312 20262
rect 20036 20216 20116 20244
rect 19984 20198 20036 20204
rect 20088 19922 20116 20216
rect 20260 20198 20312 20204
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19833 19612 20141 19621
rect 19833 19610 19839 19612
rect 19895 19610 19919 19612
rect 19975 19610 19999 19612
rect 20055 19610 20079 19612
rect 20135 19610 20141 19612
rect 19895 19558 19897 19610
rect 20077 19558 20079 19610
rect 19833 19556 19839 19558
rect 19895 19556 19919 19558
rect 19975 19556 19999 19558
rect 20055 19556 20079 19558
rect 20135 19556 20141 19558
rect 19833 19547 20141 19556
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19430 18864 19486 18873
rect 19340 18828 19392 18834
rect 19430 18799 19432 18808
rect 19340 18770 19392 18776
rect 19484 18799 19486 18808
rect 19432 18770 19484 18776
rect 19352 18714 19380 18770
rect 19352 18686 19564 18714
rect 19340 18624 19392 18630
rect 19392 18584 19472 18612
rect 19340 18566 19392 18572
rect 19338 18456 19394 18465
rect 19338 18391 19394 18400
rect 19352 18154 19380 18391
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19444 18057 19472 18584
rect 19536 18426 19564 18686
rect 19628 18426 19656 19382
rect 20456 19310 20484 21626
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20548 21146 20576 21422
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20352 19304 20404 19310
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 20088 19230 20300 19258
rect 20352 19246 20404 19252
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19720 18306 19748 19178
rect 20088 19174 20116 19230
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 19812 18952 19840 19110
rect 19812 18924 20116 18952
rect 19812 18834 19840 18924
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18630 20024 18770
rect 19984 18624 20036 18630
rect 20088 18612 20116 18924
rect 20180 18816 20208 19110
rect 20272 19009 20300 19230
rect 20364 19174 20392 19246
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20258 19000 20314 19009
rect 20548 18986 20576 20198
rect 20640 19310 20668 21286
rect 20732 21010 20760 21626
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 21486 21496 21558
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20718 20904 20774 20913
rect 20718 20839 20774 20848
rect 20732 20602 20760 20839
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20732 20398 20760 20538
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20904 20324 20956 20330
rect 20904 20266 20956 20272
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20732 19378 20760 19858
rect 20916 19854 20944 20266
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20824 19310 20852 19654
rect 20916 19514 20944 19654
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 21008 19310 21036 21354
rect 21456 21072 21508 21078
rect 21508 21032 21680 21060
rect 21456 21014 21508 21020
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21546 20768 21602 20777
rect 21284 20398 21312 20742
rect 21546 20703 21602 20712
rect 21560 20398 21588 20703
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21456 20256 21508 20262
rect 21362 20224 21418 20233
rect 21418 20204 21456 20210
rect 21418 20198 21508 20204
rect 21546 20224 21602 20233
rect 21418 20182 21496 20198
rect 21362 20159 21418 20168
rect 21086 20088 21142 20097
rect 21142 20046 21312 20074
rect 21086 20023 21142 20032
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20732 19122 20760 19178
rect 20810 19136 20866 19145
rect 20732 19094 20810 19122
rect 20810 19071 20866 19080
rect 20626 19000 20682 19009
rect 20548 18958 20626 18986
rect 20258 18935 20314 18944
rect 21008 18970 21036 19246
rect 20626 18935 20682 18944
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20536 18828 20588 18834
rect 20180 18788 20484 18816
rect 20260 18624 20312 18630
rect 20088 18584 20208 18612
rect 19984 18566 20036 18572
rect 19833 18524 20141 18533
rect 19833 18522 19839 18524
rect 19895 18522 19919 18524
rect 19975 18522 19999 18524
rect 20055 18522 20079 18524
rect 20135 18522 20141 18524
rect 19895 18470 19897 18522
rect 20077 18470 20079 18522
rect 19833 18468 19839 18470
rect 19895 18468 19919 18470
rect 19975 18468 19999 18470
rect 20055 18468 20079 18470
rect 20135 18468 20141 18470
rect 19833 18459 20141 18468
rect 20180 18408 20208 18584
rect 20312 18584 20392 18612
rect 20260 18566 20312 18572
rect 19536 18278 19748 18306
rect 20088 18380 20208 18408
rect 20258 18456 20314 18465
rect 20258 18391 20314 18400
rect 19430 18048 19486 18057
rect 19430 17983 19486 17992
rect 19430 17912 19486 17921
rect 19260 17870 19430 17898
rect 19430 17847 19486 17856
rect 19444 17814 19472 17847
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19156 17740 19208 17746
rect 19208 17700 19288 17728
rect 19156 17682 19208 17688
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19168 16522 19196 17478
rect 19260 17338 19288 17700
rect 19432 17672 19484 17678
rect 19338 17640 19394 17649
rect 19432 17614 19484 17620
rect 19338 17575 19340 17584
rect 19392 17575 19394 17584
rect 19340 17546 19392 17552
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 15638 18920 15846
rect 18984 15706 19012 15982
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18880 15632 18932 15638
rect 19076 15586 19104 15982
rect 18880 15574 18932 15580
rect 18984 15558 19104 15586
rect 18984 15502 19012 15558
rect 18972 15496 19024 15502
rect 18800 15456 18920 15484
rect 18892 15348 18920 15456
rect 18972 15438 19024 15444
rect 18616 15166 18736 15194
rect 18800 15320 18920 15348
rect 18970 15328 19026 15337
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18616 14482 18644 15166
rect 18694 15056 18750 15065
rect 18694 14991 18750 15000
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18236 14408 18288 14414
rect 18420 14408 18472 14414
rect 18236 14350 18288 14356
rect 18418 14376 18420 14385
rect 18472 14376 18474 14385
rect 18418 14311 18474 14320
rect 18234 13968 18290 13977
rect 18708 13938 18736 14991
rect 18800 14414 18828 15320
rect 18970 15263 19026 15272
rect 18984 15194 19012 15263
rect 18892 15166 19012 15194
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18234 13903 18290 13912
rect 18696 13932 18748 13938
rect 18248 13870 18276 13903
rect 18696 13874 18748 13880
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17868 13184 17920 13190
rect 17406 13152 17462 13161
rect 17972 13161 18000 13194
rect 17868 13126 17920 13132
rect 17958 13152 18014 13161
rect 17406 13087 17462 13096
rect 17958 13087 18014 13096
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17328 12617 17356 12650
rect 17592 12640 17644 12646
rect 17314 12608 17370 12617
rect 17592 12582 17644 12588
rect 17314 12543 17370 12552
rect 17604 12434 17632 12582
rect 17420 12406 17632 12434
rect 17420 12306 17448 12406
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11801 17632 12038
rect 17130 11792 17186 11801
rect 17130 11727 17186 11736
rect 17590 11792 17646 11801
rect 17590 11727 17646 11736
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 10810 16988 11154
rect 17144 11082 17172 11727
rect 17696 11286 17724 12174
rect 17788 11898 17816 12922
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17880 12306 17908 12650
rect 17972 12646 18000 13087
rect 18064 12782 18092 13398
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18248 12442 18276 13806
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 13258 18552 13670
rect 18892 13274 18920 15166
rect 19168 14890 19196 16458
rect 19260 16250 19288 17002
rect 19444 16522 19472 17614
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19536 16402 19564 18278
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19628 17241 19656 17682
rect 19614 17232 19670 17241
rect 19720 17202 19748 18158
rect 20088 18154 20116 18380
rect 20272 18358 20300 18391
rect 20260 18352 20312 18358
rect 20166 18320 20222 18329
rect 20260 18294 20312 18300
rect 20166 18255 20222 18264
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19812 17746 19840 17818
rect 20180 17814 20208 18255
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19833 17436 20141 17445
rect 19833 17434 19839 17436
rect 19895 17434 19919 17436
rect 19975 17434 19999 17436
rect 20055 17434 20079 17436
rect 20135 17434 20141 17436
rect 19895 17382 19897 17434
rect 20077 17382 20079 17434
rect 19833 17380 19839 17382
rect 19895 17380 19919 17382
rect 19975 17380 19999 17382
rect 20055 17380 20079 17382
rect 20135 17380 20141 17382
rect 19833 17371 20141 17380
rect 20258 17368 20314 17377
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 20180 17326 20258 17354
rect 19904 17241 19932 17274
rect 19890 17232 19946 17241
rect 19614 17167 19670 17176
rect 19708 17196 19760 17202
rect 19890 17167 19946 17176
rect 19708 17138 19760 17144
rect 19904 16658 19932 17167
rect 20180 16658 20208 17326
rect 20364 17354 20392 18584
rect 20456 18426 20484 18788
rect 20536 18770 20588 18776
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20314 17326 20392 17354
rect 20258 17303 20314 17312
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 19708 16652 19760 16658
rect 19892 16652 19944 16658
rect 19760 16612 19840 16640
rect 19708 16594 19760 16600
rect 19812 16538 19840 16612
rect 19892 16594 19944 16600
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 19984 16584 20036 16590
rect 19812 16532 19984 16538
rect 19812 16526 20036 16532
rect 19708 16516 19760 16522
rect 19812 16510 20024 16526
rect 20168 16516 20220 16522
rect 19708 16458 19760 16464
rect 20168 16458 20220 16464
rect 19352 16374 19564 16402
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15366 19288 16050
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19062 14648 19118 14657
rect 19062 14583 19118 14592
rect 19076 14414 19104 14583
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 18984 13938 19012 14350
rect 19168 14278 19196 14826
rect 19352 14618 19380 16374
rect 19628 16289 19656 16390
rect 19614 16280 19670 16289
rect 19614 16215 19670 16224
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19444 15706 19472 15914
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19522 15600 19578 15609
rect 19522 15535 19524 15544
rect 19576 15535 19578 15544
rect 19524 15506 19576 15512
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19444 14482 19472 14758
rect 19536 14657 19564 15098
rect 19628 14890 19656 15914
rect 19720 15638 19748 16458
rect 19833 16348 20141 16357
rect 19833 16346 19839 16348
rect 19895 16346 19919 16348
rect 19975 16346 19999 16348
rect 20055 16346 20079 16348
rect 20135 16346 20141 16348
rect 19895 16294 19897 16346
rect 20077 16294 20079 16346
rect 19833 16292 19839 16294
rect 19895 16292 19919 16294
rect 19975 16292 19999 16294
rect 20055 16292 20079 16294
rect 20135 16292 20141 16294
rect 19833 16283 20141 16292
rect 20076 16108 20128 16114
rect 19812 16068 20076 16096
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19812 15484 19840 16068
rect 20076 16050 20128 16056
rect 20180 15978 20208 16458
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20074 15736 20130 15745
rect 20074 15671 20130 15680
rect 19720 15456 19840 15484
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19522 14648 19578 14657
rect 19522 14583 19524 14592
rect 19576 14583 19578 14592
rect 19720 14600 19748 15456
rect 20088 15366 20116 15671
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19833 15260 20141 15269
rect 19833 15258 19839 15260
rect 19895 15258 19919 15260
rect 19975 15258 19999 15260
rect 20055 15258 20079 15260
rect 20135 15258 20141 15260
rect 19895 15206 19897 15258
rect 20077 15206 20079 15258
rect 19833 15204 19839 15206
rect 19895 15204 19919 15206
rect 19975 15204 19999 15206
rect 20055 15204 20079 15206
rect 20135 15204 20141 15206
rect 19833 15195 20141 15204
rect 20180 15162 20208 15914
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 19984 15088 20036 15094
rect 20036 15036 20116 15042
rect 19984 15030 20116 15036
rect 19996 15014 20116 15030
rect 19892 14816 19944 14822
rect 19890 14784 19892 14793
rect 19984 14816 20036 14822
rect 19944 14784 19946 14793
rect 19984 14758 20036 14764
rect 19890 14719 19946 14728
rect 19720 14572 19840 14600
rect 19524 14554 19576 14560
rect 19522 14512 19578 14521
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19432 14476 19484 14482
rect 19522 14447 19578 14456
rect 19706 14512 19762 14521
rect 19812 14482 19840 14572
rect 19996 14550 20024 14758
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19706 14447 19762 14456
rect 19800 14476 19852 14482
rect 19432 14418 19484 14424
rect 19260 14278 19288 14418
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19352 14074 19380 14350
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18984 13530 19012 13874
rect 19444 13870 19472 14418
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19248 13320 19300 13326
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18512 13252 18564 13258
rect 18892 13246 19196 13274
rect 19248 13262 19300 13268
rect 18512 13194 18564 13200
rect 18340 12986 18368 13194
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18418 13016 18474 13025
rect 18328 12980 18380 12986
rect 18418 12951 18420 12960
rect 18328 12922 18380 12928
rect 18472 12951 18474 12960
rect 18420 12922 18472 12928
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17880 11898 17908 12242
rect 17972 12209 18000 12242
rect 17958 12200 18014 12209
rect 17958 12135 18014 12144
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17788 11218 17816 11290
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 17236 10130 17264 11086
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10130 17356 10406
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 17328 9382 17356 10066
rect 17420 9722 17448 10542
rect 17880 10266 17908 11834
rect 18064 11762 18092 12106
rect 18156 11898 18184 12378
rect 18432 12306 18460 12650
rect 19076 12646 19104 13126
rect 19168 12918 19196 13246
rect 19260 12986 19288 13262
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19246 12880 19302 12889
rect 19246 12815 19302 12824
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19076 12442 19104 12582
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18248 11218 18276 12242
rect 18524 11778 18552 12378
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18432 11750 18552 11778
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18052 11144 18104 11150
rect 17972 11104 18052 11132
rect 17972 10674 18000 11104
rect 18052 11086 18104 11092
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17972 10112 18000 10610
rect 18064 10606 18092 10950
rect 18248 10810 18276 11154
rect 18340 11121 18368 11630
rect 18432 11558 18460 11750
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18524 11354 18552 11630
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18616 11218 18644 12174
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18708 11626 18736 12106
rect 18800 11762 18828 12242
rect 18892 11937 18920 12242
rect 19168 12238 19196 12378
rect 18972 12232 19024 12238
rect 19156 12232 19208 12238
rect 18972 12174 19024 12180
rect 19076 12192 19156 12220
rect 18878 11928 18934 11937
rect 18878 11863 18934 11872
rect 18984 11812 19012 12174
rect 18892 11784 19012 11812
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18892 11694 18920 11784
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18970 11656 19026 11665
rect 18696 11620 18748 11626
rect 18970 11591 19026 11600
rect 18696 11562 18748 11568
rect 18984 11218 19012 11591
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18420 11144 18472 11150
rect 18326 11112 18382 11121
rect 18420 11086 18472 11092
rect 18326 11047 18328 11056
rect 18380 11047 18382 11056
rect 18328 11018 18380 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18340 10146 18368 10542
rect 18432 10266 18460 11086
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18524 10266 18552 10911
rect 18616 10266 18644 11154
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10810 18736 11086
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 19076 10606 19104 12192
rect 19156 12174 19208 12180
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19168 10810 19196 10950
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 10464 19024 10470
rect 18970 10432 18972 10441
rect 19024 10432 19026 10441
rect 18970 10367 19026 10376
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 18616 10146 18644 10202
rect 18052 10124 18104 10130
rect 17972 10084 18052 10112
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17696 9722 17724 9930
rect 17408 9716 17460 9722
rect 17684 9716 17736 9722
rect 17408 9658 17460 9664
rect 17604 9676 17684 9704
rect 17604 9586 17632 9676
rect 17972 9674 18000 10084
rect 18052 10066 18104 10072
rect 18236 10124 18288 10130
rect 18340 10118 18644 10146
rect 18878 10160 18934 10169
rect 18878 10095 18880 10104
rect 18236 10066 18288 10072
rect 18932 10095 18934 10104
rect 18880 10066 18932 10072
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17684 9658 17736 9664
rect 17880 9646 18000 9674
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 16592 8634 16620 9318
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16946 8936 17002 8945
rect 16946 8871 17002 8880
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16394 8599 16450 8608
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 15946 7100 16254 7109
rect 15946 7098 15952 7100
rect 16008 7098 16032 7100
rect 16088 7098 16112 7100
rect 16168 7098 16192 7100
rect 16248 7098 16254 7100
rect 16008 7046 16010 7098
rect 16190 7046 16192 7098
rect 15946 7044 15952 7046
rect 16008 7044 16032 7046
rect 16088 7044 16112 7046
rect 16168 7044 16192 7046
rect 16248 7044 16254 7046
rect 15946 7035 16254 7044
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5914 14964 6054
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 14004 2984 14056 2990
rect 14188 2984 14240 2990
rect 14004 2926 14056 2932
rect 14186 2952 14188 2961
rect 14240 2952 14242 2961
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 10784 2848 10836 2854
rect 10612 2808 10784 2836
rect 10324 2790 10376 2796
rect 10784 2790 10836 2796
rect 9692 2746 9996 2774
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9692 2514 9720 2746
rect 13556 2582 13584 2858
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 14016 2514 14044 2926
rect 14186 2887 14242 2896
rect 14200 2774 14228 2887
rect 14200 2746 14320 2774
rect 14292 2514 14320 2746
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14200 2394 14228 2450
rect 14568 2394 14596 3470
rect 14936 3194 14964 5102
rect 15028 4214 15056 5510
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15304 4826 15332 5170
rect 15580 5137 15608 6122
rect 15856 5846 15884 6598
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 15946 6012 16254 6021
rect 15946 6010 15952 6012
rect 16008 6010 16032 6012
rect 16088 6010 16112 6012
rect 16168 6010 16192 6012
rect 16248 6010 16254 6012
rect 16008 5958 16010 6010
rect 16190 5958 16192 6010
rect 15946 5956 15952 5958
rect 16008 5956 16032 5958
rect 16088 5956 16112 5958
rect 16168 5956 16192 5958
rect 16248 5956 16254 5958
rect 15946 5947 16254 5956
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 16316 5710 16344 6054
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16132 5302 16160 5646
rect 16210 5400 16266 5409
rect 16210 5335 16266 5344
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16224 5166 16252 5335
rect 15752 5160 15804 5166
rect 15566 5128 15622 5137
rect 15566 5063 15622 5072
rect 15750 5128 15752 5137
rect 16212 5160 16264 5166
rect 15804 5128 15806 5137
rect 15750 5063 15806 5072
rect 15856 5120 16212 5148
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15474 4992 15530 5001
rect 15396 4826 15424 4966
rect 15474 4927 15530 4936
rect 15488 4826 15516 4927
rect 15750 4856 15806 4865
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15476 4820 15528 4826
rect 15750 4791 15752 4800
rect 15476 4762 15528 4768
rect 15804 4791 15806 4800
rect 15752 4762 15804 4768
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15028 4078 15056 4150
rect 15120 4078 15148 4558
rect 15212 4162 15240 4762
rect 15856 4706 15884 5120
rect 16212 5102 16264 5108
rect 15946 4924 16254 4933
rect 15946 4922 15952 4924
rect 16008 4922 16032 4924
rect 16088 4922 16112 4924
rect 16168 4922 16192 4924
rect 16248 4922 16254 4924
rect 16008 4870 16010 4922
rect 16190 4870 16192 4922
rect 15946 4868 15952 4870
rect 16008 4868 16032 4870
rect 16088 4868 16112 4870
rect 16168 4868 16192 4870
rect 16248 4868 16254 4870
rect 15946 4859 16254 4868
rect 15396 4690 15884 4706
rect 15384 4684 15884 4690
rect 15436 4678 15884 4684
rect 15384 4626 15436 4632
rect 15212 4134 15332 4162
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3618 15148 3878
rect 15212 3738 15240 3946
rect 15304 3738 15332 4134
rect 15396 4078 15424 4626
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15120 3590 15240 3618
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15212 2514 15240 3590
rect 15304 3058 15332 3674
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15396 3194 15424 3538
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15488 3194 15516 3334
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15396 2514 15424 3130
rect 15580 3058 15608 4490
rect 15672 4282 15700 4490
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16040 4078 16068 4218
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16224 4010 16252 4558
rect 16316 4146 16344 5646
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 15946 3836 16254 3845
rect 15946 3834 15952 3836
rect 16008 3834 16032 3836
rect 16088 3834 16112 3836
rect 16168 3834 16192 3836
rect 16248 3834 16254 3836
rect 16008 3782 16010 3834
rect 16190 3782 16192 3834
rect 15946 3780 15952 3782
rect 16008 3780 16032 3782
rect 16088 3780 16112 3782
rect 16168 3780 16192 3782
rect 16248 3780 16254 3782
rect 15946 3771 16254 3780
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15672 2650 15700 2926
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15856 2582 15884 2926
rect 16408 2922 16436 8230
rect 16592 8090 16620 8298
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16684 8022 16712 8502
rect 16776 8430 16804 8774
rect 16868 8498 16896 8774
rect 16960 8498 16988 8871
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7478 16528 7686
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16500 6798 16528 7414
rect 16776 7206 16804 8026
rect 16868 7410 16896 8434
rect 17052 8022 17080 9046
rect 17420 8634 17448 9454
rect 17696 8634 17724 9454
rect 17880 9382 17908 9646
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 18156 8514 18184 9862
rect 18248 9722 18276 10066
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8906 18460 8978
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 17972 8486 18184 8514
rect 17972 8430 18000 8486
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17052 7886 17080 7958
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16592 6633 16620 6831
rect 16856 6656 16908 6662
rect 16578 6624 16634 6633
rect 16856 6598 16908 6604
rect 16578 6559 16634 6568
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 5030 16528 6054
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16578 4856 16634 4865
rect 16578 4791 16634 4800
rect 16592 4486 16620 4791
rect 16684 4570 16712 6258
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16776 4826 16804 5306
rect 16868 5302 16896 6598
rect 16960 6497 16988 7142
rect 17500 6928 17552 6934
rect 17604 6916 17632 7822
rect 17696 7342 17724 7822
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17552 6888 17632 6916
rect 17500 6870 17552 6876
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 16946 6488 17002 6497
rect 17696 6458 17724 6802
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17880 6458 17908 7346
rect 17972 6984 18000 8230
rect 18064 7546 18092 8366
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7342 18184 8486
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 7585 18276 7890
rect 18234 7576 18290 7585
rect 18234 7511 18290 7520
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 17972 6956 18276 6984
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 16946 6423 17002 6432
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17052 5778 17080 6122
rect 17972 5778 18000 6666
rect 18064 6458 18092 6802
rect 18248 6798 18276 6956
rect 18340 6934 18368 7278
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18432 6798 18460 8298
rect 18524 7342 18552 9318
rect 18616 8974 18644 9454
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18616 7954 18644 8910
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18708 7410 18736 8842
rect 18984 8022 19012 9862
rect 19168 9518 19196 10202
rect 19260 9926 19288 12815
rect 19352 12434 19380 13806
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12714 19472 13126
rect 19536 12918 19564 14447
rect 19720 14249 19748 14447
rect 19800 14418 19852 14424
rect 20088 14260 20116 15014
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14414 20208 14894
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19706 14240 19762 14249
rect 20088 14232 20208 14260
rect 19706 14175 19762 14184
rect 19833 14172 20141 14181
rect 19833 14170 19839 14172
rect 19895 14170 19919 14172
rect 19975 14170 19999 14172
rect 20055 14170 20079 14172
rect 20135 14170 20141 14172
rect 19895 14118 19897 14170
rect 20077 14118 20079 14170
rect 19833 14116 19839 14118
rect 19895 14116 19919 14118
rect 19975 14116 19999 14118
rect 20055 14116 20079 14118
rect 20135 14116 20141 14118
rect 19833 14107 20141 14116
rect 20180 13802 20208 14232
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 19706 13424 19762 13433
rect 19616 13388 19668 13394
rect 20272 13394 20300 17138
rect 20456 16289 20484 18362
rect 20548 17678 20576 18770
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20640 18358 20668 18702
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20534 17504 20590 17513
rect 20534 17439 20590 17448
rect 20548 17134 20576 17439
rect 20640 17270 20668 18294
rect 20732 17746 20760 18362
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20824 17814 20852 18294
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20626 17096 20682 17105
rect 20548 16658 20576 17070
rect 20626 17031 20682 17040
rect 20640 16794 20668 17031
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20732 16522 20760 17682
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 17134 20852 17614
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20442 16280 20498 16289
rect 20442 16215 20498 16224
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15745 20392 15914
rect 20350 15736 20406 15745
rect 20350 15671 20406 15680
rect 20456 15502 20484 16215
rect 20824 16114 20852 17070
rect 20916 16658 20944 18906
rect 21192 18834 21220 19858
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 18086 21036 18566
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17338 21036 17614
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20994 16960 21050 16969
rect 20994 16895 21050 16904
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20628 16040 20680 16046
rect 20548 16000 20628 16028
rect 20548 15502 20576 16000
rect 20628 15982 20680 15988
rect 20718 16008 20774 16017
rect 20916 15994 20944 16186
rect 21008 16114 21036 16895
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20718 15943 20774 15952
rect 20824 15966 20944 15994
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20640 15337 20668 15506
rect 20626 15328 20682 15337
rect 20626 15263 20682 15272
rect 20534 15192 20590 15201
rect 20534 15127 20590 15136
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 14414 20392 14758
rect 20456 14482 20484 15030
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 14074 20392 14350
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20456 14074 20484 14282
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 13954 20576 15127
rect 20640 14890 20668 15263
rect 20732 14929 20760 15943
rect 20824 15434 20852 15966
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15570 21036 15846
rect 20996 15564 21048 15570
rect 20916 15524 20996 15552
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20916 15026 20944 15524
rect 20996 15506 21048 15512
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20996 14952 21048 14958
rect 20718 14920 20774 14929
rect 20628 14884 20680 14890
rect 20996 14894 21048 14900
rect 20718 14855 20774 14864
rect 20628 14826 20680 14832
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 14074 20668 14214
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20456 13926 20576 13954
rect 20456 13394 20484 13926
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 19706 13359 19762 13368
rect 20260 13388 20312 13394
rect 19616 13330 19668 13336
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19628 12646 19656 13330
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19720 12434 19748 13359
rect 20260 13330 20312 13336
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 19833 13084 20141 13093
rect 19833 13082 19839 13084
rect 19895 13082 19919 13084
rect 19975 13082 19999 13084
rect 20055 13082 20079 13084
rect 20135 13082 20141 13084
rect 19895 13030 19897 13082
rect 20077 13030 20079 13082
rect 19833 13028 19839 13030
rect 19895 13028 19919 13030
rect 19975 13028 19999 13030
rect 20055 13028 20079 13030
rect 20135 13028 20141 13030
rect 19833 13019 20141 13028
rect 20180 12986 20208 13194
rect 20272 13161 20300 13330
rect 20352 13184 20404 13190
rect 20258 13152 20314 13161
rect 20352 13126 20404 13132
rect 20258 13087 20314 13096
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20076 12912 20128 12918
rect 20074 12880 20076 12889
rect 20128 12880 20130 12889
rect 20364 12850 20392 13126
rect 20548 12986 20576 13466
rect 20732 13394 20760 14010
rect 20916 13734 20944 14758
rect 21008 14618 21036 14894
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20074 12815 20130 12824
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20628 12776 20680 12782
rect 20442 12744 20498 12753
rect 20628 12718 20680 12724
rect 20442 12679 20498 12688
rect 19352 12406 19472 12434
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19352 11014 19380 11562
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10742 19380 10950
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19338 10432 19394 10441
rect 19444 10418 19472 12406
rect 19628 12406 19748 12434
rect 20168 12436 20220 12442
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19536 10470 19564 11698
rect 19394 10390 19472 10418
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19338 10367 19394 10376
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19154 9072 19210 9081
rect 19154 9007 19210 9016
rect 19168 8634 19196 9007
rect 19260 8974 19288 9454
rect 19352 9382 19380 9998
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19260 8566 19288 8910
rect 19248 8560 19300 8566
rect 19154 8528 19210 8537
rect 19248 8502 19300 8508
rect 19154 8463 19210 8472
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 19168 7886 19196 8463
rect 19338 7984 19394 7993
rect 19338 7919 19340 7928
rect 19392 7919 19394 7928
rect 19340 7890 19392 7896
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18156 6390 18184 6734
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18432 6338 18460 6734
rect 18984 6730 19012 7346
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18616 6458 18644 6598
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17960 5772 18012 5778
rect 18156 5760 18184 6326
rect 18432 6310 18552 6338
rect 18524 6254 18552 6310
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18248 5914 18276 6122
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18236 5772 18288 5778
rect 18156 5732 18236 5760
rect 17960 5714 18012 5720
rect 18236 5714 18288 5720
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 16868 4826 16896 5238
rect 17052 5166 17080 5714
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16684 4542 16804 4570
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4146 16712 4422
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16684 3398 16712 3878
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3194 16712 3334
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16776 2990 16804 4542
rect 17052 4486 17080 5102
rect 17144 4826 17172 5170
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17236 4758 17264 4966
rect 17788 4826 17816 5714
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18064 5234 18092 5646
rect 18340 5409 18368 6122
rect 18326 5400 18382 5409
rect 18326 5335 18382 5344
rect 18432 5234 18460 6190
rect 18892 5846 18920 6666
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18064 4826 18092 5170
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18326 5128 18382 5137
rect 18156 4826 18184 5102
rect 18326 5063 18382 5072
rect 18340 4826 18368 5063
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4078 17816 4422
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3534 17172 3878
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3194 16896 3334
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 15946 2748 16254 2757
rect 15946 2746 15952 2748
rect 16008 2746 16032 2748
rect 16088 2746 16112 2748
rect 16168 2746 16192 2748
rect 16248 2746 16254 2748
rect 16008 2694 16010 2746
rect 16190 2694 16192 2746
rect 15946 2692 15952 2694
rect 16008 2692 16032 2694
rect 16088 2692 16112 2694
rect 16168 2692 16192 2694
rect 16248 2692 16254 2694
rect 15946 2683 16254 2692
rect 15844 2576 15896 2582
rect 15844 2518 15896 2524
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 14200 2366 14596 2394
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 4285 2204 4593 2213
rect 4285 2202 4291 2204
rect 4347 2202 4371 2204
rect 4427 2202 4451 2204
rect 4507 2202 4531 2204
rect 4587 2202 4593 2204
rect 4347 2150 4349 2202
rect 4529 2150 4531 2202
rect 4285 2148 4291 2150
rect 4347 2148 4371 2150
rect 4427 2148 4451 2150
rect 4507 2148 4531 2150
rect 4587 2148 4593 2150
rect 4285 2139 4593 2148
rect 12059 2204 12367 2213
rect 12059 2202 12065 2204
rect 12121 2202 12145 2204
rect 12201 2202 12225 2204
rect 12281 2202 12305 2204
rect 12361 2202 12367 2204
rect 12121 2150 12123 2202
rect 12303 2150 12305 2202
rect 12059 2148 12065 2150
rect 12121 2148 12145 2150
rect 12201 2148 12225 2150
rect 12281 2148 12305 2150
rect 12361 2148 12367 2150
rect 12059 2139 12367 2148
rect 8172 1660 8480 1669
rect 8172 1658 8178 1660
rect 8234 1658 8258 1660
rect 8314 1658 8338 1660
rect 8394 1658 8418 1660
rect 8474 1658 8480 1660
rect 8234 1606 8236 1658
rect 8416 1606 8418 1658
rect 8172 1604 8178 1606
rect 8234 1604 8258 1606
rect 8314 1604 8338 1606
rect 8394 1604 8418 1606
rect 8474 1604 8480 1606
rect 8172 1595 8480 1604
rect 14200 1494 14228 2366
rect 15304 2106 15332 2382
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15764 1766 15792 2382
rect 15856 2106 15884 2518
rect 16592 2446 16620 2790
rect 16776 2774 16804 2926
rect 16684 2746 16804 2774
rect 16684 2514 16712 2746
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 15844 2100 15896 2106
rect 15844 2042 15896 2048
rect 16592 1902 16620 2382
rect 17144 2106 17172 2926
rect 17328 2650 17356 4014
rect 18156 3890 18184 4490
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 17880 3862 18184 3890
rect 17880 3602 17908 3862
rect 18156 3738 18184 3862
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17420 2990 17448 3538
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17512 3194 17540 3402
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17132 2100 17184 2106
rect 17132 2042 17184 2048
rect 17512 2038 17540 3130
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17604 2650 17632 2858
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17696 2650 17724 2790
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17696 2514 17724 2586
rect 17972 2514 18000 3674
rect 18248 2650 18276 4150
rect 18432 2922 18460 5170
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 4078 18828 4422
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18524 2514 18552 2586
rect 18616 2514 18644 3130
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18708 2774 18736 2858
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18708 2746 18828 2774
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18800 2446 18828 2746
rect 18892 2650 18920 2790
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18156 2106 18184 2314
rect 18892 2106 18920 2586
rect 18984 2446 19012 5578
rect 19076 3738 19104 7822
rect 19444 7002 19472 10202
rect 19628 9602 19656 12406
rect 19812 12396 20168 12424
rect 19812 12102 19840 12396
rect 20168 12378 20220 12384
rect 20166 12336 20222 12345
rect 20166 12271 20168 12280
rect 20220 12271 20222 12280
rect 20168 12242 20220 12248
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19833 11996 20141 12005
rect 19833 11994 19839 11996
rect 19895 11994 19919 11996
rect 19975 11994 19999 11996
rect 20055 11994 20079 11996
rect 20135 11994 20141 11996
rect 19895 11942 19897 11994
rect 20077 11942 20079 11994
rect 19833 11940 19839 11942
rect 19895 11940 19919 11942
rect 19975 11940 19999 11942
rect 20055 11940 20079 11942
rect 20135 11940 20141 11942
rect 19833 11931 20141 11940
rect 20180 11830 20208 12106
rect 20272 11898 20300 12106
rect 20350 11928 20406 11937
rect 20260 11892 20312 11898
rect 20350 11863 20406 11872
rect 20260 11834 20312 11840
rect 20168 11824 20220 11830
rect 20364 11778 20392 11863
rect 20456 11830 20484 12679
rect 20640 12374 20668 12718
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20220 11772 20392 11778
rect 20168 11766 20392 11772
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20180 11750 20392 11766
rect 20364 11694 20392 11750
rect 20352 11688 20404 11694
rect 19798 11656 19854 11665
rect 20352 11630 20404 11636
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 19798 11591 19854 11600
rect 19812 11286 19840 11591
rect 20456 11393 20484 11630
rect 20442 11384 20498 11393
rect 20548 11354 20576 12174
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20442 11319 20498 11328
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 20640 11218 20668 12106
rect 20732 11830 20760 13330
rect 20824 12986 20852 13398
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20824 12782 20852 12922
rect 20916 12918 20944 13670
rect 21008 13190 21036 13738
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20824 11830 20852 12271
rect 20916 12238 20944 12650
rect 20996 12436 21048 12442
rect 21100 12434 21128 17002
rect 21192 16114 21220 18634
rect 21284 18630 21312 20046
rect 21362 19952 21418 19961
rect 21468 19922 21496 20182
rect 21546 20159 21602 20168
rect 21560 19990 21588 20159
rect 21652 20058 21680 21032
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21362 19887 21418 19896
rect 21456 19916 21508 19922
rect 21376 19768 21404 19887
rect 21456 19858 21508 19864
rect 21456 19780 21508 19786
rect 21376 19740 21456 19768
rect 21456 19722 21508 19728
rect 21362 19680 21418 19689
rect 21362 19615 21418 19624
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21270 18456 21326 18465
rect 21270 18391 21326 18400
rect 21284 18358 21312 18391
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21376 17649 21404 19615
rect 21468 19553 21496 19722
rect 21454 19544 21510 19553
rect 21454 19479 21510 19488
rect 21652 19378 21680 19994
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21836 19310 21864 20946
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21928 20602 21956 20810
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21928 19553 21956 19858
rect 21914 19544 21970 19553
rect 21914 19479 21970 19488
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21454 19000 21510 19009
rect 21454 18935 21510 18944
rect 21640 18964 21692 18970
rect 21468 18834 21496 18935
rect 21640 18906 21692 18912
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21362 17640 21418 17649
rect 21362 17575 21418 17584
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17184 21312 17478
rect 21284 17156 21404 17184
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21284 16794 21312 17002
rect 21376 16998 21404 17156
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21364 16584 21416 16590
rect 21270 16552 21326 16561
rect 21364 16526 21416 16532
rect 21270 16487 21326 16496
rect 21284 16454 21312 16487
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 16114 21312 16390
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 21192 15881 21220 15914
rect 21284 15910 21312 16050
rect 21272 15904 21324 15910
rect 21178 15872 21234 15881
rect 21272 15846 21324 15852
rect 21178 15807 21234 15816
rect 21376 15570 21404 16526
rect 21468 15570 21496 18770
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21560 17882 21588 18702
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21652 17814 21680 18906
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 21638 17640 21694 17649
rect 21638 17575 21694 17584
rect 21652 16998 21680 17575
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21640 16788 21692 16794
rect 21744 16776 21772 19246
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 21692 16748 21772 16776
rect 21640 16730 21692 16736
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21560 16425 21588 16594
rect 21546 16416 21602 16425
rect 21546 16351 21602 16360
rect 21560 15978 21588 16351
rect 21548 15972 21600 15978
rect 21548 15914 21600 15920
rect 21546 15872 21602 15881
rect 21546 15807 21602 15816
rect 21560 15638 21588 15807
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21192 14278 21220 14894
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21284 14618 21312 14826
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21376 14414 21404 15506
rect 21652 14958 21680 16730
rect 21836 16250 21864 17682
rect 21928 16561 21956 18022
rect 22020 17134 22048 21626
rect 23940 21480 23992 21486
rect 23992 21428 24256 21434
rect 23940 21422 24256 21428
rect 23952 21406 24256 21422
rect 24228 21350 24256 21406
rect 24124 21344 24176 21350
rect 23386 21312 23442 21321
rect 24124 21286 24176 21292
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 23386 21247 23442 21256
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22388 20942 22416 21082
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22834 21040 22890 21049
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 19854 22232 20402
rect 22282 20224 22338 20233
rect 22282 20159 22338 20168
rect 22296 19990 22324 20159
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22388 19922 22416 20878
rect 22480 20262 22508 21014
rect 23400 21010 23428 21247
rect 23720 21244 24028 21253
rect 23720 21242 23726 21244
rect 23782 21242 23806 21244
rect 23862 21242 23886 21244
rect 23942 21242 23966 21244
rect 24022 21242 24028 21244
rect 23782 21190 23784 21242
rect 23964 21190 23966 21242
rect 23720 21188 23726 21190
rect 23782 21188 23806 21190
rect 23862 21188 23886 21190
rect 23942 21188 23966 21190
rect 24022 21188 24028 21190
rect 23720 21179 24028 21188
rect 24136 21146 24164 21286
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 22834 20975 22836 20984
rect 22888 20975 22890 20984
rect 22928 21004 22980 21010
rect 22836 20946 22888 20952
rect 22928 20946 22980 20952
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22572 20074 22600 20538
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22480 20046 22600 20074
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22112 19446 22140 19790
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22204 19242 22232 19314
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22112 16574 22140 18566
rect 22296 17542 22324 19450
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22388 18970 22416 19110
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22480 18850 22508 20046
rect 22664 19378 22692 20198
rect 22742 19816 22798 19825
rect 22742 19751 22798 19760
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22572 18970 22600 19246
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22664 18850 22692 19178
rect 22388 18822 22508 18850
rect 22572 18822 22692 18850
rect 22388 18426 22416 18822
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22284 17264 22336 17270
rect 21914 16552 21970 16561
rect 21914 16487 21970 16496
rect 22020 16546 22140 16574
rect 22204 17224 22284 17252
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21916 16244 21968 16250
rect 22020 16232 22048 16546
rect 22204 16454 22232 17224
rect 22284 17206 22336 17212
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22284 17128 22336 17134
rect 22282 17096 22284 17105
rect 22388 17116 22416 17206
rect 22336 17096 22416 17116
rect 22338 17088 22416 17096
rect 22480 17048 22508 18294
rect 22572 17105 22600 18822
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22664 18057 22692 18634
rect 22756 18290 22784 19751
rect 22940 19224 22968 20946
rect 23308 20602 23336 20946
rect 23584 20602 23612 20946
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23294 20496 23350 20505
rect 23350 20454 23520 20482
rect 23676 20466 23704 20878
rect 23860 20874 23888 21014
rect 24492 21004 24544 21010
rect 24492 20946 24544 20952
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23754 20496 23810 20505
rect 23294 20431 23350 20440
rect 23110 20360 23166 20369
rect 23110 20295 23166 20304
rect 23388 20324 23440 20330
rect 23020 19848 23072 19854
rect 23018 19816 23020 19825
rect 23072 19816 23074 19825
rect 23018 19751 23074 19760
rect 23124 19378 23152 20295
rect 23388 20266 23440 20272
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23112 19236 23164 19242
rect 22940 19196 23112 19224
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22848 18222 22876 19110
rect 22940 18970 22968 19196
rect 23112 19178 23164 19184
rect 23216 19145 23244 19246
rect 23308 19174 23336 19994
rect 23400 19922 23428 20266
rect 23492 19922 23520 20454
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23664 20460 23716 20466
rect 23754 20431 23810 20440
rect 23664 20402 23716 20408
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23492 19553 23520 19858
rect 23584 19718 23612 20402
rect 23768 20330 23796 20431
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 23756 20324 23808 20330
rect 23756 20266 23808 20272
rect 23720 20156 24028 20165
rect 23720 20154 23726 20156
rect 23782 20154 23806 20156
rect 23862 20154 23886 20156
rect 23942 20154 23966 20156
rect 24022 20154 24028 20156
rect 23782 20102 23784 20154
rect 23964 20102 23966 20154
rect 23720 20100 23726 20102
rect 23782 20100 23806 20102
rect 23862 20100 23886 20102
rect 23942 20100 23966 20102
rect 24022 20100 24028 20102
rect 23720 20091 24028 20100
rect 24320 19922 24348 20334
rect 24400 19984 24452 19990
rect 24400 19926 24452 19932
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23478 19544 23534 19553
rect 23388 19508 23440 19514
rect 23478 19479 23534 19488
rect 23388 19450 23440 19456
rect 23296 19168 23348 19174
rect 23202 19136 23258 19145
rect 23296 19110 23348 19116
rect 23202 19071 23258 19080
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22940 18329 22968 18702
rect 23032 18358 23060 18906
rect 23216 18834 23244 19071
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23020 18352 23072 18358
rect 22926 18320 22982 18329
rect 23020 18294 23072 18300
rect 22926 18255 22982 18264
rect 23112 18284 23164 18290
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22650 18048 22706 18057
rect 22650 17983 22706 17992
rect 22282 17031 22338 17040
rect 22388 17020 22508 17048
rect 22558 17096 22614 17105
rect 22558 17031 22614 17040
rect 22282 16824 22338 16833
rect 22282 16759 22338 16768
rect 22296 16726 22324 16759
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 21968 16204 22048 16232
rect 21916 16186 21968 16192
rect 21928 16046 21956 16186
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21744 14414 21772 14962
rect 21928 14618 21956 15982
rect 22204 15570 22232 16390
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22006 15056 22062 15065
rect 22204 15026 22232 15506
rect 22006 14991 22062 15000
rect 22192 15020 22244 15026
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21822 14376 21878 14385
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21560 14006 21588 14350
rect 21744 14074 21772 14350
rect 21822 14311 21878 14320
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21192 13394 21220 13466
rect 21560 13394 21588 13738
rect 21652 13530 21680 13806
rect 21836 13530 21864 14311
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21284 12782 21312 12922
rect 21272 12776 21324 12782
rect 21324 12736 21404 12764
rect 21272 12718 21324 12724
rect 21100 12406 21312 12434
rect 20996 12378 21048 12384
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 21008 11694 21036 12378
rect 21088 12300 21140 12306
rect 21140 12260 21220 12288
rect 21088 12242 21140 12248
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21100 11694 21128 12106
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 19708 11144 19760 11150
rect 19706 11112 19708 11121
rect 19760 11112 19762 11121
rect 19706 11047 19762 11056
rect 19720 10266 19748 11047
rect 19833 10908 20141 10917
rect 19833 10906 19839 10908
rect 19895 10906 19919 10908
rect 19975 10906 19999 10908
rect 20055 10906 20079 10908
rect 20135 10906 20141 10908
rect 19895 10854 19897 10906
rect 20077 10854 20079 10906
rect 19833 10852 19839 10854
rect 19895 10852 19919 10854
rect 19975 10852 19999 10854
rect 20055 10852 20079 10854
rect 20135 10852 20141 10854
rect 19833 10843 20141 10852
rect 20364 10810 20392 11154
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20456 10577 20484 10950
rect 20442 10568 20498 10577
rect 20168 10532 20220 10538
rect 20442 10503 20498 10512
rect 20168 10474 20220 10480
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19833 9820 20141 9829
rect 19833 9818 19839 9820
rect 19895 9818 19919 9820
rect 19975 9818 19999 9820
rect 20055 9818 20079 9820
rect 20135 9818 20141 9820
rect 19895 9766 19897 9818
rect 20077 9766 20079 9818
rect 19833 9764 19839 9766
rect 19895 9764 19919 9766
rect 19975 9764 19999 9766
rect 20055 9764 20079 9766
rect 20135 9764 20141 9766
rect 19833 9755 20141 9764
rect 19536 9574 19656 9602
rect 19536 8294 19564 9574
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19628 7546 19656 9386
rect 19996 9178 20024 9386
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8514 19748 8910
rect 19833 8732 20141 8741
rect 19833 8730 19839 8732
rect 19895 8730 19919 8732
rect 19975 8730 19999 8732
rect 20055 8730 20079 8732
rect 20135 8730 20141 8732
rect 19895 8678 19897 8730
rect 20077 8678 20079 8730
rect 19833 8676 19839 8678
rect 19895 8676 19919 8678
rect 19975 8676 19999 8678
rect 20055 8676 20079 8678
rect 20135 8676 20141 8678
rect 19833 8667 20141 8676
rect 19798 8528 19854 8537
rect 19720 8486 19798 8514
rect 19798 8463 19800 8472
rect 19852 8463 19854 8472
rect 19800 8434 19852 8440
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19260 6089 19288 6122
rect 19246 6080 19302 6089
rect 19246 6015 19302 6024
rect 19352 5817 19380 6598
rect 19720 6390 19748 7958
rect 20180 7818 20208 10474
rect 20548 10198 20576 11086
rect 20720 11008 20772 11014
rect 20824 10996 20852 11290
rect 20916 11286 20944 11494
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20772 10968 20852 10996
rect 20720 10950 20772 10956
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20548 10062 20576 10134
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20640 9704 20668 10406
rect 20916 10033 20944 10406
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 20640 9676 20760 9704
rect 20626 9616 20682 9625
rect 20626 9551 20682 9560
rect 20640 9382 20668 9551
rect 20732 9432 20760 9676
rect 21008 9654 21036 10134
rect 21192 9897 21220 12260
rect 21178 9888 21234 9897
rect 21100 9846 21178 9874
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 20996 9444 21048 9450
rect 20732 9404 20996 9432
rect 20996 9386 21048 9392
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20272 8362 20300 9114
rect 20548 9081 20576 9318
rect 20534 9072 20590 9081
rect 20534 9007 20590 9016
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20258 7848 20314 7857
rect 20168 7812 20220 7818
rect 20258 7783 20314 7792
rect 20168 7754 20220 7760
rect 19833 7644 20141 7653
rect 19833 7642 19839 7644
rect 19895 7642 19919 7644
rect 19975 7642 19999 7644
rect 20055 7642 20079 7644
rect 20135 7642 20141 7644
rect 19895 7590 19897 7642
rect 20077 7590 20079 7642
rect 19833 7588 19839 7590
rect 19895 7588 19919 7590
rect 19975 7588 19999 7590
rect 20055 7588 20079 7590
rect 20135 7588 20141 7590
rect 19833 7579 20141 7588
rect 20076 7336 20128 7342
rect 20180 7324 20208 7754
rect 20128 7296 20208 7324
rect 20076 7278 20128 7284
rect 20166 7168 20222 7177
rect 20166 7103 20222 7112
rect 20180 6866 20208 7103
rect 20272 7002 20300 7783
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20272 6866 20300 6938
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 19812 6662 19840 6802
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 19833 6556 20141 6565
rect 19833 6554 19839 6556
rect 19895 6554 19919 6556
rect 19975 6554 19999 6556
rect 20055 6554 20079 6556
rect 20135 6554 20141 6556
rect 19895 6502 19897 6554
rect 20077 6502 20079 6554
rect 19833 6500 19839 6502
rect 19895 6500 19919 6502
rect 19975 6500 19999 6502
rect 20055 6500 20079 6502
rect 20135 6500 20141 6502
rect 19833 6491 20141 6500
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19338 5808 19394 5817
rect 19338 5743 19394 5752
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19444 5234 19472 5510
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19260 4690 19288 4966
rect 19352 4690 19380 5034
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19536 4604 19564 5714
rect 19628 5370 19656 6054
rect 19812 5914 19840 6190
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19996 5846 20024 6190
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 20088 5778 20116 6122
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19720 5302 19748 5646
rect 19833 5468 20141 5477
rect 19833 5466 19839 5468
rect 19895 5466 19919 5468
rect 19975 5466 19999 5468
rect 20055 5466 20079 5468
rect 20135 5466 20141 5468
rect 19895 5414 19897 5466
rect 20077 5414 20079 5466
rect 19833 5412 19839 5414
rect 19895 5412 19919 5414
rect 19975 5412 19999 5414
rect 20055 5412 20079 5414
rect 20135 5412 20141 5414
rect 19833 5403 20141 5412
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19616 4616 19668 4622
rect 19536 4576 19616 4604
rect 19616 4558 19668 4564
rect 19156 4548 19208 4554
rect 19156 4490 19208 4496
rect 19168 4078 19196 4490
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4078 19472 4422
rect 19628 4146 19656 4558
rect 19720 4282 19748 5102
rect 19833 4380 20141 4389
rect 19833 4378 19839 4380
rect 19895 4378 19919 4380
rect 19975 4378 19999 4380
rect 20055 4378 20079 4380
rect 20135 4378 20141 4380
rect 19895 4326 19897 4378
rect 20077 4326 20079 4378
rect 19833 4324 19839 4326
rect 19895 4324 19919 4326
rect 19975 4324 19999 4326
rect 20055 4324 20079 4326
rect 20135 4324 20141 4326
rect 19833 4315 20141 4324
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19720 4078 19748 4218
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19076 3602 19104 3674
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19076 2514 19104 2790
rect 19352 2514 19380 2790
rect 19444 2514 19472 3878
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19628 3058 19656 3402
rect 19720 3058 19748 3878
rect 20088 3466 20116 4014
rect 20180 3602 20208 6598
rect 20260 6316 20312 6322
rect 20364 6304 20392 8570
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20456 8106 20484 8434
rect 20534 8120 20590 8129
rect 20456 8078 20534 8106
rect 20456 8022 20484 8078
rect 20534 8055 20590 8064
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20456 7177 20484 7958
rect 20442 7168 20498 7177
rect 20442 7103 20498 7112
rect 20548 7041 20576 7958
rect 20640 7886 20668 9318
rect 21100 9194 21128 9846
rect 21178 9823 21234 9832
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 20732 9166 21128 9194
rect 20732 8838 20760 9166
rect 21192 9110 21220 9658
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20720 7744 20772 7750
rect 20718 7712 20720 7721
rect 20812 7744 20864 7750
rect 20772 7712 20774 7721
rect 20812 7686 20864 7692
rect 20718 7647 20774 7656
rect 20824 7478 20852 7686
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20534 7032 20590 7041
rect 20534 6967 20590 6976
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20444 6724 20496 6730
rect 20548 6712 20576 6802
rect 20496 6684 20576 6712
rect 20444 6666 20496 6672
rect 20364 6276 20484 6304
rect 20260 6258 20312 6264
rect 20272 5778 20300 6258
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5098 20300 5510
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20456 5030 20484 6276
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 5846 20576 6122
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20628 5772 20680 5778
rect 20904 5772 20956 5778
rect 20680 5732 20852 5760
rect 20628 5714 20680 5720
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20548 5030 20576 5510
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20456 4690 20484 4966
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20548 4214 20576 4966
rect 20824 4690 20852 5732
rect 20904 5714 20956 5720
rect 20916 4690 20944 5714
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20536 4208 20588 4214
rect 20442 4176 20498 4185
rect 20272 4134 20442 4162
rect 20272 4078 20300 4134
rect 20536 4150 20588 4156
rect 20442 4111 20498 4120
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3738 20300 3878
rect 20364 3738 20392 4014
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19833 3292 20141 3301
rect 19833 3290 19839 3292
rect 19895 3290 19919 3292
rect 19975 3290 19999 3292
rect 20055 3290 20079 3292
rect 20135 3290 20141 3292
rect 19895 3238 19897 3290
rect 20077 3238 20079 3290
rect 19833 3236 19839 3238
rect 19895 3236 19919 3238
rect 19975 3236 19999 3238
rect 20055 3236 20079 3238
rect 20135 3236 20141 3238
rect 19833 3227 20141 3236
rect 20272 3074 20300 3538
rect 20456 3194 20484 4014
rect 20916 3618 20944 4626
rect 21008 3738 21036 7822
rect 21192 6730 21220 7890
rect 21284 7342 21312 12406
rect 21376 11898 21404 12736
rect 21468 11898 21496 13126
rect 21560 12646 21588 13126
rect 21652 12646 21680 13466
rect 21928 13190 21956 14554
rect 22020 14396 22048 14991
rect 22192 14962 22244 14968
rect 22100 14408 22152 14414
rect 22020 14368 22100 14396
rect 22020 14113 22048 14368
rect 22100 14350 22152 14356
rect 22006 14104 22062 14113
rect 22006 14039 22062 14048
rect 22006 13968 22062 13977
rect 22006 13903 22008 13912
rect 22060 13903 22062 13912
rect 22008 13874 22060 13880
rect 22204 13530 22232 14962
rect 22296 13841 22324 16662
rect 22388 14958 22416 17020
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22572 15706 22600 16594
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 15586 22692 17983
rect 22940 17610 22968 18255
rect 23112 18226 23164 18232
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22928 17604 22980 17610
rect 22928 17546 22980 17552
rect 22940 17134 22968 17546
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 22756 16454 22784 16662
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22848 16114 22876 16390
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22940 16046 22968 16458
rect 23032 16250 23060 18158
rect 23124 17082 23152 18226
rect 23216 17814 23244 18770
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23308 17649 23336 17818
rect 23294 17640 23350 17649
rect 23294 17575 23350 17584
rect 23124 17054 23244 17082
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23124 16658 23152 16934
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 23020 15632 23072 15638
rect 22480 15558 22692 15586
rect 22940 15592 23020 15620
rect 22744 15564 22796 15570
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22388 14618 22416 14894
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22480 14346 22508 15558
rect 22744 15506 22796 15512
rect 22560 15360 22612 15366
rect 22756 15314 22784 15506
rect 22834 15464 22890 15473
rect 22834 15399 22890 15408
rect 22560 15302 22612 15308
rect 22572 15162 22600 15302
rect 22664 15286 22784 15314
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22664 14498 22692 15286
rect 22848 15162 22876 15399
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22756 15042 22784 15098
rect 22834 15056 22890 15065
rect 22756 15014 22834 15042
rect 22834 14991 22890 15000
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22756 14521 22784 14826
rect 22572 14470 22692 14498
rect 22742 14512 22798 14521
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22282 13832 22338 13841
rect 22282 13767 22338 13776
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22572 13433 22600 14470
rect 22742 14447 22798 14456
rect 22848 14278 22876 14894
rect 22940 14890 22968 15592
rect 23020 15574 23072 15580
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23032 14958 23060 15098
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22928 14884 22980 14890
rect 22928 14826 22980 14832
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22664 13462 22692 13806
rect 22756 13802 22784 14010
rect 22940 13870 22968 14418
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22652 13456 22704 13462
rect 22558 13424 22614 13433
rect 22100 13388 22152 13394
rect 22652 13398 22704 13404
rect 22756 13394 22784 13738
rect 22558 13359 22614 13368
rect 22744 13388 22796 13394
rect 22100 13330 22152 13336
rect 22744 13330 22796 13336
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 22006 13152 22062 13161
rect 22006 13087 22062 13096
rect 22020 12850 22048 13087
rect 22112 12986 22140 13330
rect 22756 12986 22784 13330
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22468 12776 22520 12782
rect 22756 12753 22784 12922
rect 22928 12844 22980 12850
rect 23032 12832 23060 14350
rect 22980 12804 23060 12832
rect 22928 12786 22980 12792
rect 22468 12718 22520 12724
rect 22742 12744 22798 12753
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 22296 12442 22324 12718
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 21730 12336 21786 12345
rect 21928 12306 21956 12378
rect 22192 12368 22244 12374
rect 22192 12310 22244 12316
rect 21730 12271 21786 12280
rect 21916 12300 21968 12306
rect 21744 12238 21772 12271
rect 21916 12242 21968 12248
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21732 12096 21784 12102
rect 21730 12064 21732 12073
rect 22100 12096 22152 12102
rect 21784 12064 21786 12073
rect 22100 12038 22152 12044
rect 21730 11999 21786 12008
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21362 11520 21418 11529
rect 21362 11455 21418 11464
rect 21376 11286 21404 11455
rect 21468 11354 21496 11630
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21914 11248 21970 11257
rect 21914 11183 21916 11192
rect 21968 11183 21970 11192
rect 21916 11154 21968 11160
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21468 10588 21496 10746
rect 21640 10600 21692 10606
rect 21468 10560 21640 10588
rect 21640 10542 21692 10548
rect 21652 10266 21680 10542
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21362 9616 21418 9625
rect 21362 9551 21418 9560
rect 21376 9178 21404 9551
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8634 21404 9114
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21100 5710 21128 6190
rect 21192 5914 21220 6394
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21100 5302 21128 5646
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 21192 4758 21220 5850
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21192 4078 21220 4694
rect 21284 4078 21312 6326
rect 21376 5273 21404 6326
rect 21362 5264 21418 5273
rect 21362 5199 21418 5208
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21180 4072 21232 4078
rect 21272 4072 21324 4078
rect 21180 4014 21232 4020
rect 21270 4040 21272 4049
rect 21324 4040 21326 4049
rect 21270 3975 21326 3984
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20732 3590 20944 3618
rect 20994 3632 21050 3641
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20548 3194 20576 3334
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20732 3126 20760 3590
rect 20994 3567 20996 3576
rect 21048 3567 21050 3576
rect 21376 3584 21404 4490
rect 21560 4026 21588 7346
rect 21652 7274 21680 9998
rect 21744 9722 21772 11018
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21744 9178 21772 9318
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21836 8974 21864 9590
rect 21928 9518 21956 11154
rect 22112 11150 22140 12038
rect 22204 11762 22232 12310
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11830 22324 12038
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22204 11014 22232 11698
rect 22296 11694 22324 11766
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22480 10062 22508 12718
rect 22742 12679 22798 12688
rect 23124 12594 23152 16186
rect 23216 15706 23244 17054
rect 23308 16658 23336 17575
rect 23296 16652 23348 16658
rect 23296 16594 23348 16600
rect 23400 16250 23428 19450
rect 23584 19224 23612 19654
rect 23768 19334 23796 19654
rect 23952 19378 23980 19858
rect 23676 19310 23796 19334
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 23664 19306 23796 19310
rect 23664 19304 23716 19306
rect 23664 19246 23716 19252
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23492 19196 23612 19224
rect 23492 18630 23520 19196
rect 23860 19156 23888 19246
rect 23584 19128 23888 19156
rect 24124 19168 24176 19174
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23492 17882 23520 18158
rect 23584 17921 23612 19128
rect 24124 19110 24176 19116
rect 23720 19068 24028 19077
rect 23720 19066 23726 19068
rect 23782 19066 23806 19068
rect 23862 19066 23886 19068
rect 23942 19066 23966 19068
rect 24022 19066 24028 19068
rect 23782 19014 23784 19066
rect 23964 19014 23966 19066
rect 23720 19012 23726 19014
rect 23782 19012 23806 19014
rect 23862 19012 23886 19014
rect 23942 19012 23966 19014
rect 24022 19012 24028 19014
rect 23720 19003 24028 19012
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23768 18222 23796 18838
rect 24136 18766 24164 19110
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 24044 18222 24072 18566
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23720 17980 24028 17989
rect 23720 17978 23726 17980
rect 23782 17978 23806 17980
rect 23862 17978 23886 17980
rect 23942 17978 23966 17980
rect 24022 17978 24028 17980
rect 23782 17926 23784 17978
rect 23964 17926 23966 17978
rect 23720 17924 23726 17926
rect 23782 17924 23806 17926
rect 23862 17924 23886 17926
rect 23942 17924 23966 17926
rect 24022 17924 24028 17926
rect 23570 17912 23626 17921
rect 23720 17915 24028 17924
rect 23480 17876 23532 17882
rect 23570 17847 23626 17856
rect 23480 17818 23532 17824
rect 23584 17814 23612 17847
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23216 14278 23244 15506
rect 23308 14958 23336 15846
rect 23386 15736 23442 15745
rect 23386 15671 23388 15680
rect 23440 15671 23442 15680
rect 23388 15642 23440 15648
rect 23386 15600 23442 15609
rect 23386 15535 23442 15544
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23294 14512 23350 14521
rect 23400 14482 23428 15535
rect 23492 15502 23520 17206
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23584 16522 23612 17138
rect 23768 17066 23796 17206
rect 23952 17202 23980 17478
rect 24136 17338 24164 18362
rect 24228 17513 24256 19314
rect 24320 18290 24348 19858
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24320 17921 24348 18226
rect 24306 17912 24362 17921
rect 24306 17847 24362 17856
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 24214 17504 24270 17513
rect 24214 17439 24270 17448
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24216 17264 24268 17270
rect 24030 17232 24086 17241
rect 23940 17196 23992 17202
rect 24086 17212 24216 17218
rect 24086 17206 24268 17212
rect 24086 17190 24256 17206
rect 24030 17167 24086 17176
rect 23940 17138 23992 17144
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23720 16892 24028 16901
rect 23720 16890 23726 16892
rect 23782 16890 23806 16892
rect 23862 16890 23886 16892
rect 23942 16890 23966 16892
rect 24022 16890 24028 16892
rect 23782 16838 23784 16890
rect 23964 16838 23966 16890
rect 23720 16836 23726 16838
rect 23782 16836 23806 16838
rect 23862 16836 23886 16838
rect 23942 16836 23966 16838
rect 24022 16836 24028 16838
rect 23720 16827 24028 16836
rect 24122 16824 24178 16833
rect 24122 16759 24178 16768
rect 23938 16552 23994 16561
rect 23572 16516 23624 16522
rect 23938 16487 23994 16496
rect 23572 16458 23624 16464
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23584 15881 23612 15982
rect 23952 15978 23980 16487
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23570 15872 23626 15881
rect 23570 15807 23626 15816
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23584 15366 23612 15807
rect 23720 15804 24028 15813
rect 23720 15802 23726 15804
rect 23782 15802 23806 15804
rect 23862 15802 23886 15804
rect 23942 15802 23966 15804
rect 24022 15802 24028 15804
rect 23782 15750 23784 15802
rect 23964 15750 23966 15802
rect 23720 15748 23726 15750
rect 23782 15748 23806 15750
rect 23862 15748 23886 15750
rect 23942 15748 23966 15750
rect 24022 15748 24028 15750
rect 23720 15739 24028 15748
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23492 14550 23520 15098
rect 23768 15026 23796 15574
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 15026 23980 15506
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 24044 14958 24072 15642
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23720 14716 24028 14725
rect 23720 14714 23726 14716
rect 23782 14714 23806 14716
rect 23862 14714 23886 14716
rect 23942 14714 23966 14716
rect 24022 14714 24028 14716
rect 23782 14662 23784 14714
rect 23964 14662 23966 14714
rect 23720 14660 23726 14662
rect 23782 14660 23806 14662
rect 23862 14660 23886 14662
rect 23942 14660 23966 14662
rect 24022 14660 24028 14662
rect 23720 14651 24028 14660
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23294 14447 23350 14456
rect 23388 14476 23440 14482
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 23216 13326 23244 13738
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12714 23244 13262
rect 23308 13258 23336 14447
rect 23388 14418 23440 14424
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23860 14074 23888 14418
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 23952 14113 23980 14282
rect 23938 14104 23994 14113
rect 23848 14068 23900 14074
rect 23938 14039 23994 14048
rect 23848 14010 23900 14016
rect 23860 13870 23888 14010
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 24044 13734 24072 14282
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 23584 13394 23612 13670
rect 23720 13628 24028 13637
rect 23720 13626 23726 13628
rect 23782 13626 23806 13628
rect 23862 13626 23886 13628
rect 23942 13626 23966 13628
rect 24022 13626 24028 13628
rect 23782 13574 23784 13626
rect 23964 13574 23966 13626
rect 23720 13572 23726 13574
rect 23782 13572 23806 13574
rect 23862 13572 23886 13574
rect 23942 13572 23966 13574
rect 24022 13572 24028 13574
rect 23720 13563 24028 13572
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23204 12708 23256 12714
rect 23204 12650 23256 12656
rect 23584 12646 23612 13330
rect 23676 12986 23704 13330
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23572 12640 23624 12646
rect 23124 12566 23244 12594
rect 24044 12628 24072 13330
rect 24136 12850 24164 16759
rect 24228 16726 24256 17190
rect 24320 16726 24348 17614
rect 24412 16726 24440 19926
rect 24504 18426 24532 20946
rect 24596 20466 24624 21966
rect 30380 22024 30432 22030
rect 26884 21966 26936 21972
rect 29734 21992 29790 22001
rect 26054 21927 26110 21936
rect 25320 21888 25372 21894
rect 24674 21856 24730 21865
rect 25320 21830 25372 21836
rect 24674 21791 24730 21800
rect 24688 21486 24716 21791
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 21350 24900 21422
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24674 20768 24730 20777
rect 24674 20703 24730 20712
rect 24688 20602 24716 20703
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24504 17746 24532 18226
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24216 16720 24268 16726
rect 24216 16662 24268 16668
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 24400 16720 24452 16726
rect 24400 16662 24452 16668
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24228 15638 24256 16186
rect 24320 15706 24348 16662
rect 24412 16250 24440 16662
rect 24596 16454 24624 20402
rect 24688 19990 24716 20538
rect 24872 20330 24900 21286
rect 25332 21010 25360 21830
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25884 21434 25912 21490
rect 26068 21486 26096 21927
rect 26606 21856 26662 21865
rect 26606 21791 26662 21800
rect 26620 21486 26648 21791
rect 26056 21480 26108 21486
rect 25884 21406 26004 21434
rect 26056 21422 26108 21428
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25410 21040 25466 21049
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25320 21004 25372 21010
rect 25410 20975 25412 20984
rect 25320 20946 25372 20952
rect 25464 20975 25466 20984
rect 25504 21004 25556 21010
rect 25412 20946 25464 20952
rect 25504 20946 25556 20952
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25148 20602 25176 20946
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25516 20534 25544 20946
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25608 20466 25636 20810
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24676 19984 24728 19990
rect 24676 19926 24728 19932
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24780 19553 24808 19858
rect 24766 19544 24822 19553
rect 24872 19514 24900 20266
rect 24964 20058 24992 20334
rect 25700 20262 25728 20946
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25332 19922 25360 20198
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25596 19916 25648 19922
rect 25596 19858 25648 19864
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 24766 19479 24822 19488
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18970 24716 19246
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24780 18408 24808 19382
rect 24872 18630 24900 19450
rect 25148 19446 25176 19790
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 24952 18760 25004 18766
rect 24950 18728 24952 18737
rect 25044 18760 25096 18766
rect 25004 18728 25006 18737
rect 25044 18702 25096 18708
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 24950 18663 25006 18672
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24860 18420 24912 18426
rect 24780 18380 24860 18408
rect 24860 18362 24912 18368
rect 24860 18216 24912 18222
rect 24674 18184 24730 18193
rect 24860 18158 24912 18164
rect 24674 18119 24676 18128
rect 24728 18119 24730 18128
rect 24676 18090 24728 18096
rect 24872 17785 24900 18158
rect 25056 17882 25084 18702
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 24858 17776 24914 17785
rect 24858 17711 24860 17720
rect 24912 17711 24914 17720
rect 24860 17682 24912 17688
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17377 24900 17478
rect 24858 17368 24914 17377
rect 24676 17332 24728 17338
rect 24858 17303 24914 17312
rect 24676 17274 24728 17280
rect 24688 16794 24716 17274
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24228 15337 24256 15370
rect 24214 15328 24270 15337
rect 24214 15263 24270 15272
rect 24320 15026 24348 15642
rect 24412 15570 24440 15846
rect 24872 15706 24900 17303
rect 25044 16720 25096 16726
rect 24964 16680 25044 16708
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24216 14884 24268 14890
rect 24216 14826 24268 14832
rect 24228 14793 24256 14826
rect 24214 14784 24270 14793
rect 24214 14719 24270 14728
rect 24320 13462 24348 14962
rect 24412 14074 24440 15506
rect 24688 15434 24716 15642
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24490 15328 24546 15337
rect 24490 15263 24546 15272
rect 24504 14822 24532 15263
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24504 14006 24532 14758
rect 24596 14006 24624 15370
rect 24858 14920 24914 14929
rect 24858 14855 24914 14864
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24398 13832 24454 13841
rect 24398 13767 24400 13776
rect 24452 13767 24454 13776
rect 24400 13738 24452 13744
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24044 12600 24164 12628
rect 23572 12582 23624 12588
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22664 12209 22692 12242
rect 22650 12200 22706 12209
rect 22560 12164 22612 12170
rect 22650 12135 22706 12144
rect 22560 12106 22612 12112
rect 22572 11898 22600 12106
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22848 11665 22876 12038
rect 22834 11656 22890 11665
rect 22834 11591 22890 11600
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22940 10538 22968 10950
rect 23032 10674 23060 11086
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22928 10532 22980 10538
rect 22928 10474 22980 10480
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22664 10062 22692 10202
rect 22940 10198 22968 10474
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 22020 8430 22048 9386
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22572 9110 22600 9318
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22376 9036 22428 9042
rect 22428 8996 22508 9024
rect 22376 8978 22428 8984
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21744 7857 21772 8230
rect 21916 7880 21968 7886
rect 21730 7848 21786 7857
rect 21916 7822 21968 7828
rect 21730 7783 21786 7792
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21652 6866 21680 7210
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21744 6322 21772 7783
rect 21928 7342 21956 7822
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21928 6934 21956 7278
rect 21916 6928 21968 6934
rect 21916 6870 21968 6876
rect 22204 6730 22232 8910
rect 22480 8430 22508 8996
rect 22572 8498 22600 9046
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22374 7984 22430 7993
rect 22374 7919 22376 7928
rect 22428 7919 22430 7928
rect 22376 7890 22428 7896
rect 22480 7342 22508 8366
rect 22284 7336 22336 7342
rect 22468 7336 22520 7342
rect 22336 7296 22416 7324
rect 22284 7278 22336 7284
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 21822 6624 21878 6633
rect 21822 6559 21878 6568
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21652 5778 21680 6122
rect 21744 5778 21772 6258
rect 21836 6254 21864 6559
rect 22006 6488 22062 6497
rect 22006 6423 22062 6432
rect 22020 6254 22048 6423
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 21836 5778 21864 6190
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21652 5302 21680 5714
rect 21744 5370 21772 5714
rect 21916 5636 21968 5642
rect 21916 5578 21968 5584
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21744 4758 21772 4966
rect 21836 4826 21864 4966
rect 21928 4826 21956 5578
rect 22112 5234 22140 6190
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22098 5128 22154 5137
rect 22020 5086 22098 5114
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21824 4548 21876 4554
rect 21824 4490 21876 4496
rect 21836 4298 21864 4490
rect 22020 4298 22048 5086
rect 22098 5063 22154 5072
rect 21836 4270 22048 4298
rect 21836 4078 21864 4270
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21824 4072 21876 4078
rect 21560 3998 21680 4026
rect 21824 4014 21876 4020
rect 21914 4040 21970 4049
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21468 3738 21496 3878
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 21456 3596 21508 3602
rect 21376 3556 21456 3584
rect 20996 3538 21048 3544
rect 21456 3538 21508 3544
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19812 3046 20300 3074
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 19628 2514 19656 2994
rect 19812 2990 19840 3046
rect 20272 2990 20300 3046
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19984 2984 20036 2990
rect 20260 2984 20312 2990
rect 19984 2926 20036 2932
rect 20074 2952 20130 2961
rect 19996 2854 20024 2926
rect 20260 2926 20312 2932
rect 20074 2887 20130 2896
rect 20088 2854 20116 2887
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 19996 2514 20024 2790
rect 20824 2514 20852 3334
rect 20916 2774 20944 3470
rect 21468 3369 21496 3538
rect 21454 3360 21510 3369
rect 21454 3295 21510 3304
rect 21468 2938 21496 3295
rect 21560 2990 21588 3878
rect 21284 2922 21496 2938
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 21652 2938 21680 3998
rect 22020 4026 22048 4082
rect 22204 4026 22232 6054
rect 22296 5642 22324 7142
rect 22388 5914 22416 7296
rect 22468 7278 22520 7284
rect 22480 6934 22508 7278
rect 22664 7274 22692 9998
rect 23124 9625 23152 10406
rect 22834 9616 22890 9625
rect 22834 9551 22890 9560
rect 23110 9616 23166 9625
rect 23110 9551 23166 9560
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8129 22784 8978
rect 22742 8120 22798 8129
rect 22742 8055 22798 8064
rect 22756 8022 22784 8055
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22480 6322 22508 6870
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22468 6112 22520 6118
rect 22466 6080 22468 6089
rect 22520 6080 22522 6089
rect 22466 6015 22522 6024
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 22296 5370 22324 5578
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22296 4690 22324 5306
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22480 5114 22508 6015
rect 22572 5778 22600 7142
rect 22650 6896 22706 6905
rect 22650 6831 22706 6840
rect 22664 6798 22692 6831
rect 22652 6792 22704 6798
rect 22848 6769 22876 9551
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23124 8634 23152 9046
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23216 8537 23244 12566
rect 23720 12540 24028 12549
rect 23720 12538 23726 12540
rect 23782 12538 23806 12540
rect 23862 12538 23886 12540
rect 23942 12538 23966 12540
rect 24022 12538 24028 12540
rect 23782 12486 23784 12538
rect 23964 12486 23966 12538
rect 23720 12484 23726 12486
rect 23782 12484 23806 12486
rect 23862 12484 23886 12486
rect 23942 12484 23966 12486
rect 24022 12484 24028 12486
rect 23720 12475 24028 12484
rect 24136 12442 24164 12600
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 23754 12336 23810 12345
rect 23754 12271 23756 12280
rect 23808 12271 23810 12280
rect 24032 12300 24084 12306
rect 23756 12242 23808 12248
rect 24032 12242 24084 12248
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23308 9994 23336 11562
rect 23400 11558 23428 12174
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23572 12096 23624 12102
rect 23768 12073 23796 12106
rect 23572 12038 23624 12044
rect 23754 12064 23810 12073
rect 23584 11898 23612 12038
rect 23754 11999 23810 12008
rect 24044 11898 24072 12242
rect 24136 12238 24164 12378
rect 24228 12238 24256 13330
rect 24400 13320 24452 13326
rect 24306 13288 24362 13297
rect 24400 13262 24452 13268
rect 24306 13223 24362 13232
rect 24320 13190 24348 13223
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24412 12646 24440 13262
rect 24596 12986 24624 13942
rect 24688 13394 24716 14554
rect 24872 14550 24900 14855
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24780 13870 24808 14418
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 14006 24900 14214
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24490 12744 24546 12753
rect 24780 12714 24808 13806
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24872 12986 24900 13670
rect 24964 13530 24992 16680
rect 25044 16662 25096 16668
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25056 13530 25084 15506
rect 25148 14958 25176 18702
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 16833 25268 18022
rect 25332 17746 25360 19858
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 25332 17270 25360 17682
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25320 16992 25372 16998
rect 25318 16960 25320 16969
rect 25372 16960 25374 16969
rect 25318 16895 25374 16904
rect 25226 16824 25282 16833
rect 25226 16759 25282 16768
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25240 16454 25268 16662
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25424 15586 25452 18090
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25516 16522 25544 17206
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 16153 25544 16458
rect 25502 16144 25558 16153
rect 25502 16079 25558 16088
rect 25332 15558 25452 15586
rect 25228 15496 25280 15502
rect 25332 15473 25360 15558
rect 25412 15496 25464 15502
rect 25228 15438 25280 15444
rect 25318 15464 25374 15473
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25240 14482 25268 15438
rect 25412 15438 25464 15444
rect 25318 15399 25374 15408
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25332 14958 25360 15302
rect 25424 15094 25452 15438
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25228 14476 25280 14482
rect 25148 14436 25228 14464
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24490 12679 24546 12688
rect 24768 12708 24820 12714
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 12442 24440 12582
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23400 10130 23428 10610
rect 23492 10538 23520 11834
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 23720 11452 24028 11461
rect 23720 11450 23726 11452
rect 23782 11450 23806 11452
rect 23862 11450 23886 11452
rect 23942 11450 23966 11452
rect 24022 11450 24028 11452
rect 23782 11398 23784 11450
rect 23964 11398 23966 11450
rect 23720 11396 23726 11398
rect 23782 11396 23806 11398
rect 23862 11396 23886 11398
rect 23942 11396 23966 11398
rect 24022 11396 24028 11398
rect 23720 11387 24028 11396
rect 24124 11144 24176 11150
rect 24320 11098 24348 11562
rect 24176 11092 24348 11098
rect 24124 11086 24348 11092
rect 24136 11070 24348 11086
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23720 10364 24028 10373
rect 23720 10362 23726 10364
rect 23782 10362 23806 10364
rect 23862 10362 23886 10364
rect 23942 10362 23966 10364
rect 24022 10362 24028 10364
rect 23782 10310 23784 10362
rect 23964 10310 23966 10362
rect 23720 10308 23726 10310
rect 23782 10308 23806 10310
rect 23862 10308 23886 10310
rect 23942 10308 23966 10310
rect 24022 10308 24028 10310
rect 23720 10299 24028 10308
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23940 10124 23992 10130
rect 24320 10112 24348 11070
rect 24412 10810 24440 12378
rect 24504 12306 24532 12679
rect 24768 12650 24820 12656
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12458 24716 12582
rect 24766 12472 24822 12481
rect 24688 12430 24766 12458
rect 24766 12407 24822 12416
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24872 12186 24900 12718
rect 25056 12714 25084 12922
rect 25148 12850 25176 14436
rect 25228 14418 25280 14424
rect 25226 14376 25282 14385
rect 25226 14311 25282 14320
rect 25240 13802 25268 14311
rect 25332 13841 25360 14894
rect 25412 13864 25464 13870
rect 25318 13832 25374 13841
rect 25228 13796 25280 13802
rect 25412 13806 25464 13812
rect 25318 13767 25374 13776
rect 25228 13738 25280 13744
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 25148 12356 25176 12786
rect 25424 12782 25452 13806
rect 25608 13394 25636 19858
rect 25700 18154 25728 20198
rect 25688 18148 25740 18154
rect 25688 18090 25740 18096
rect 25792 17898 25820 20946
rect 25884 19310 25912 21286
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 25884 18154 25912 18294
rect 25872 18148 25924 18154
rect 25872 18090 25924 18096
rect 25792 17870 25912 17898
rect 25780 17740 25832 17746
rect 25700 17700 25780 17728
rect 25700 16114 25728 17700
rect 25780 17682 25832 17688
rect 25780 17604 25832 17610
rect 25780 17546 25832 17552
rect 25792 16794 25820 17546
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 25792 16250 25820 16458
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25700 15502 25728 16050
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25688 15088 25740 15094
rect 25686 15056 25688 15065
rect 25740 15056 25742 15065
rect 25686 14991 25742 15000
rect 25792 14550 25820 16050
rect 25884 15201 25912 17870
rect 25870 15192 25926 15201
rect 25870 15127 25926 15136
rect 25780 14544 25832 14550
rect 25780 14486 25832 14492
rect 25884 14482 25912 15127
rect 25872 14476 25924 14482
rect 25872 14418 25924 14424
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25884 13530 25912 14282
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25792 13410 25820 13466
rect 25596 13388 25648 13394
rect 25792 13382 25912 13410
rect 25596 13330 25648 13336
rect 25608 12986 25636 13330
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12986 25820 13126
rect 25884 12986 25912 13382
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25686 12472 25742 12481
rect 25686 12407 25742 12416
rect 25700 12374 25728 12407
rect 25228 12368 25280 12374
rect 25148 12328 25228 12356
rect 25228 12310 25280 12316
rect 25688 12368 25740 12374
rect 25688 12310 25740 12316
rect 24872 12170 25084 12186
rect 24872 12164 25096 12170
rect 24872 12158 25044 12164
rect 25044 12106 25096 12112
rect 24858 11792 24914 11801
rect 24858 11727 24914 11736
rect 24872 11694 24900 11727
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24582 11112 24638 11121
rect 24582 11047 24638 11056
rect 24596 10810 24624 11047
rect 24688 11014 24716 11222
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24584 10804 24636 10810
rect 24584 10746 24636 10752
rect 24596 10266 24624 10746
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24584 10124 24636 10130
rect 24320 10084 24584 10112
rect 23940 10066 23992 10072
rect 24584 10066 24636 10072
rect 23664 10056 23716 10062
rect 23662 10024 23664 10033
rect 23716 10024 23718 10033
rect 23296 9988 23348 9994
rect 23348 9948 23520 9976
rect 23662 9959 23718 9968
rect 23756 9988 23808 9994
rect 23296 9930 23348 9936
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23400 9518 23428 9658
rect 23492 9654 23520 9948
rect 23860 9976 23888 10066
rect 23808 9948 23888 9976
rect 23756 9930 23808 9936
rect 23952 9926 23980 10066
rect 24214 10024 24270 10033
rect 24214 9959 24270 9968
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23202 8528 23258 8537
rect 23112 8492 23164 8498
rect 23308 8498 23336 9318
rect 23202 8463 23204 8472
rect 23112 8434 23164 8440
rect 23256 8463 23258 8472
rect 23296 8492 23348 8498
rect 23204 8434 23256 8440
rect 23296 8434 23348 8440
rect 23124 8378 23152 8434
rect 23492 8378 23520 9590
rect 23584 8634 23612 9590
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 23720 9276 24028 9285
rect 23720 9274 23726 9276
rect 23782 9274 23806 9276
rect 23862 9274 23886 9276
rect 23942 9274 23966 9276
rect 24022 9274 24028 9276
rect 23782 9222 23784 9274
rect 23964 9222 23966 9274
rect 23720 9220 23726 9222
rect 23782 9220 23806 9222
rect 23862 9220 23886 9222
rect 23942 9220 23966 9222
rect 24022 9220 24028 9222
rect 23720 9211 24028 9220
rect 24136 9178 24164 9454
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 23756 8968 23808 8974
rect 24228 8945 24256 9959
rect 24398 9888 24454 9897
rect 24398 9823 24454 9832
rect 24412 9586 24440 9823
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24308 9512 24360 9518
rect 24688 9466 24716 10950
rect 24780 10130 24808 11494
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24964 10713 24992 10950
rect 24950 10704 25006 10713
rect 24950 10639 25006 10648
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25700 10266 25728 10406
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 24308 9454 24360 9460
rect 23756 8910 23808 8916
rect 24214 8936 24270 8945
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23768 8498 23796 8910
rect 24214 8871 24270 8880
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23124 8350 23520 8378
rect 23952 8362 23980 8570
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23400 7886 23428 8230
rect 23584 8022 23612 8230
rect 23720 8188 24028 8197
rect 23720 8186 23726 8188
rect 23782 8186 23806 8188
rect 23862 8186 23886 8188
rect 23942 8186 23966 8188
rect 24022 8186 24028 8188
rect 23782 8134 23784 8186
rect 23964 8134 23966 8186
rect 23720 8132 23726 8134
rect 23782 8132 23806 8134
rect 23862 8132 23886 8134
rect 23942 8132 23966 8134
rect 24022 8132 24028 8134
rect 23720 8123 24028 8132
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 23572 8016 23624 8022
rect 23624 7976 23704 8004
rect 23572 7958 23624 7964
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 22940 6934 22968 7822
rect 23112 7744 23164 7750
rect 23032 7692 23112 7698
rect 23400 7721 23428 7822
rect 23572 7744 23624 7750
rect 23032 7686 23164 7692
rect 23386 7712 23442 7721
rect 23032 7670 23152 7686
rect 23032 7478 23060 7670
rect 23572 7686 23624 7692
rect 23386 7647 23442 7656
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23020 7472 23072 7478
rect 23020 7414 23072 7420
rect 23216 7342 23244 7482
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 22928 6928 22980 6934
rect 22928 6870 22980 6876
rect 22652 6734 22704 6740
rect 22834 6760 22890 6769
rect 22834 6695 22890 6704
rect 22848 6186 22876 6695
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 23216 5914 23244 7278
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 23204 5908 23256 5914
rect 23308 5896 23336 6870
rect 23492 6730 23520 7142
rect 23584 6866 23612 7686
rect 23676 7546 23704 7976
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23768 7342 23796 7482
rect 23860 7342 23888 7822
rect 24136 7460 24164 8026
rect 24228 7970 24256 8871
rect 24320 8634 24348 9454
rect 24504 9438 24716 9466
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24228 7942 24348 7970
rect 24216 7472 24268 7478
rect 24136 7432 24216 7460
rect 24216 7414 24268 7420
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23720 7100 24028 7109
rect 23720 7098 23726 7100
rect 23782 7098 23806 7100
rect 23862 7098 23886 7100
rect 23942 7098 23966 7100
rect 24022 7098 24028 7100
rect 23782 7046 23784 7098
rect 23964 7046 23966 7098
rect 23720 7044 23726 7046
rect 23782 7044 23806 7046
rect 23862 7044 23886 7046
rect 23942 7044 23966 7046
rect 24022 7044 24028 7046
rect 23720 7035 24028 7044
rect 24136 6866 24164 7142
rect 24320 6866 24348 7942
rect 24412 7886 24440 9318
rect 24504 9110 24532 9438
rect 24492 9104 24544 9110
rect 24492 9046 24544 9052
rect 24504 8090 24532 9046
rect 24780 8838 24808 10066
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 24964 9926 24992 9998
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24860 9104 24912 9110
rect 24858 9072 24860 9081
rect 24912 9072 24914 9081
rect 24858 9007 24914 9016
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24688 8090 24716 8434
rect 24780 8362 24808 8774
rect 24872 8634 24900 8774
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24964 8022 24992 9590
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 24952 8016 25004 8022
rect 24952 7958 25004 7964
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 25148 7818 25176 9386
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 23308 5868 23520 5896
rect 23204 5850 23256 5856
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22848 5574 22876 5714
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22848 5166 22876 5510
rect 22940 5166 22968 5850
rect 23216 5794 23244 5850
rect 23216 5766 23428 5794
rect 23492 5778 23520 5868
rect 23584 5778 23612 6802
rect 24122 6760 24178 6769
rect 24122 6695 24178 6704
rect 24030 6352 24086 6361
rect 24030 6287 24086 6296
rect 24044 6254 24072 6287
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 24136 6186 24164 6695
rect 24124 6180 24176 6186
rect 24124 6122 24176 6128
rect 23720 6012 24028 6021
rect 23720 6010 23726 6012
rect 23782 6010 23806 6012
rect 23862 6010 23886 6012
rect 23942 6010 23966 6012
rect 24022 6010 24028 6012
rect 23782 5958 23784 6010
rect 23964 5958 23966 6010
rect 23720 5956 23726 5958
rect 23782 5956 23806 5958
rect 23862 5956 23886 5958
rect 23942 5956 23966 5958
rect 24022 5956 24028 5958
rect 23720 5947 24028 5956
rect 24136 5846 24164 6122
rect 24228 5953 24256 6802
rect 24412 6254 24440 7482
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24952 7336 25004 7342
rect 25148 7324 25176 7754
rect 25240 7750 25268 9998
rect 25424 9994 25452 10066
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25594 9888 25650 9897
rect 25516 9846 25594 9874
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25332 8294 25360 9386
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25424 7954 25452 9386
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 25424 7426 25452 7890
rect 25516 7886 25544 9846
rect 25594 9823 25650 9832
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 8090 25728 9454
rect 25792 8430 25820 10474
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 25884 9450 25912 9862
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 25884 9042 25912 9386
rect 25976 9178 26004 21406
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 26344 19922 26372 21354
rect 26896 21146 26924 21966
rect 30380 21966 30432 21972
rect 29734 21927 29790 21936
rect 28078 21856 28134 21865
rect 27607 21788 27915 21797
rect 28078 21791 28134 21800
rect 27607 21786 27613 21788
rect 27669 21786 27693 21788
rect 27749 21786 27773 21788
rect 27829 21786 27853 21788
rect 27909 21786 27915 21788
rect 27669 21734 27671 21786
rect 27851 21734 27853 21786
rect 27607 21732 27613 21734
rect 27669 21732 27693 21734
rect 27749 21732 27773 21734
rect 27829 21732 27853 21734
rect 27909 21732 27915 21734
rect 27434 21720 27490 21729
rect 27607 21723 27915 21732
rect 27434 21655 27490 21664
rect 27448 21486 27476 21655
rect 27710 21584 27766 21593
rect 27710 21519 27766 21528
rect 27724 21486 27752 21519
rect 28092 21486 28120 21791
rect 28448 21684 28500 21690
rect 28448 21626 28500 21632
rect 27436 21480 27488 21486
rect 27436 21422 27488 21428
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 27068 21072 27120 21078
rect 27068 21014 27120 21020
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26712 19990 26740 20946
rect 27080 20398 27108 21014
rect 27068 20392 27120 20398
rect 27068 20334 27120 20340
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 26804 20058 26832 20198
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26700 19984 26752 19990
rect 26700 19926 26752 19932
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26056 19712 26108 19718
rect 26344 19689 26372 19858
rect 26056 19654 26108 19660
rect 26330 19680 26386 19689
rect 26068 19310 26096 19654
rect 26330 19615 26386 19624
rect 26528 19394 26556 19858
rect 26620 19514 26648 19858
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26698 19408 26754 19417
rect 26528 19366 26648 19394
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 26424 19304 26476 19310
rect 26424 19246 26476 19252
rect 26148 19236 26200 19242
rect 26200 19196 26372 19224
rect 26148 19178 26200 19184
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26160 18426 26188 18702
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 26056 17808 26108 17814
rect 26056 17750 26108 17756
rect 26068 16250 26096 17750
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 26068 15586 26096 16186
rect 26160 15706 26188 18362
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26252 17202 26280 18294
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26238 17096 26294 17105
rect 26238 17031 26294 17040
rect 26252 16658 26280 17031
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26068 15570 26188 15586
rect 26068 15564 26200 15570
rect 26068 15558 26148 15564
rect 26148 15506 26200 15512
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26068 15337 26096 15370
rect 26054 15328 26110 15337
rect 26054 15263 26110 15272
rect 26252 14618 26280 16594
rect 26344 16425 26372 19196
rect 26436 17954 26464 19246
rect 26620 18834 26648 19366
rect 26698 19343 26754 19352
rect 26712 19174 26740 19343
rect 26700 19168 26752 19174
rect 26700 19110 26752 19116
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 18306 26648 18770
rect 26712 18426 26740 19110
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 26620 18278 26740 18306
rect 26436 17926 26556 17954
rect 26528 17746 26556 17926
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26436 16998 26464 17682
rect 26620 17649 26648 17682
rect 26606 17640 26662 17649
rect 26606 17575 26662 17584
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26330 16416 26386 16425
rect 26330 16351 26386 16360
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26344 13326 26372 16351
rect 26422 15736 26478 15745
rect 26422 15671 26478 15680
rect 26436 15638 26464 15671
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26422 14240 26478 14249
rect 26528 14226 26556 17478
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26620 16794 26648 17138
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26620 14958 26648 16730
rect 26712 15978 26740 18278
rect 26700 15972 26752 15978
rect 26700 15914 26752 15920
rect 26804 15722 26832 19790
rect 26988 19417 27016 20198
rect 27172 20058 27200 20198
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 27066 19544 27122 19553
rect 27066 19479 27122 19488
rect 26974 19408 27030 19417
rect 26974 19343 27030 19352
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26896 18970 26924 19246
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26976 18624 27028 18630
rect 26976 18566 27028 18572
rect 26988 18154 27016 18566
rect 26976 18148 27028 18154
rect 26976 18090 27028 18096
rect 27080 17882 27108 19479
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 26988 17202 27016 17478
rect 27172 17338 27200 19246
rect 27264 18290 27292 21286
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27356 20806 27384 21014
rect 27344 20800 27396 20806
rect 27344 20742 27396 20748
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27342 19816 27398 19825
rect 27342 19751 27398 19760
rect 27356 19378 27384 19751
rect 27448 19446 27476 19858
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26884 17128 26936 17134
rect 26884 17070 26936 17076
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 26896 16658 26924 17070
rect 26976 17060 27028 17066
rect 26976 17002 27028 17008
rect 26988 16969 27016 17002
rect 27080 16998 27108 17070
rect 27160 17060 27212 17066
rect 27160 17002 27212 17008
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27068 16992 27120 16998
rect 26974 16960 27030 16969
rect 27068 16934 27120 16940
rect 26974 16895 27030 16904
rect 27172 16794 27200 17002
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 26988 16658 27016 16730
rect 27264 16658 27292 17002
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26976 16652 27028 16658
rect 27252 16652 27304 16658
rect 26976 16594 27028 16600
rect 27080 16612 27252 16640
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 26712 15694 26832 15722
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26620 14482 26648 14894
rect 26712 14618 26740 15694
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26804 14940 26832 15506
rect 26988 14958 27016 16458
rect 27080 16289 27108 16612
rect 27252 16594 27304 16600
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 27066 16280 27122 16289
rect 27066 16215 27122 16224
rect 27068 16176 27120 16182
rect 27068 16118 27120 16124
rect 26884 14952 26936 14958
rect 26804 14912 26884 14940
rect 26884 14894 26936 14900
rect 26976 14952 27028 14958
rect 26976 14894 27028 14900
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26804 14482 26832 14758
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26896 14278 26924 14758
rect 26478 14198 26556 14226
rect 26884 14272 26936 14278
rect 26988 14260 27016 14894
rect 27080 14362 27108 16118
rect 27172 15026 27200 16458
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27158 14784 27214 14793
rect 27158 14719 27214 14728
rect 27172 14618 27200 14719
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27080 14334 27200 14362
rect 26988 14232 27108 14260
rect 26884 14214 26936 14220
rect 26422 14175 26478 14184
rect 26974 14104 27030 14113
rect 26974 14039 27030 14048
rect 26514 13968 26570 13977
rect 26514 13903 26570 13912
rect 26528 13802 26556 13903
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26700 13796 26752 13802
rect 26700 13738 26752 13744
rect 26712 13394 26740 13738
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26344 12345 26372 12650
rect 26330 12336 26386 12345
rect 26330 12271 26386 12280
rect 26436 12238 26464 13330
rect 26988 13326 27016 14039
rect 27080 13734 27108 14232
rect 27068 13728 27120 13734
rect 27068 13670 27120 13676
rect 26976 13320 27028 13326
rect 27068 13320 27120 13326
rect 26976 13262 27028 13268
rect 27066 13288 27068 13297
rect 27120 13288 27122 13297
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26896 12238 26924 12650
rect 26988 12646 27016 13262
rect 27066 13223 27122 13232
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26606 11928 26662 11937
rect 26896 11898 26924 12174
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26988 11898 27016 12038
rect 26606 11863 26662 11872
rect 26884 11892 26936 11898
rect 26332 11620 26384 11626
rect 26332 11562 26384 11568
rect 26344 11286 26372 11562
rect 26620 11286 26648 11863
rect 26884 11834 26936 11840
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26332 11280 26384 11286
rect 26332 11222 26384 11228
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26528 10577 26556 10678
rect 26514 10568 26570 10577
rect 26056 10532 26108 10538
rect 26514 10503 26570 10512
rect 26056 10474 26108 10480
rect 26068 10266 26096 10474
rect 26528 10266 26556 10503
rect 26056 10260 26108 10266
rect 26056 10202 26108 10208
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26620 10062 26648 11086
rect 26804 11082 26832 11630
rect 26896 11218 26924 11834
rect 27080 11218 27108 12718
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 26792 11076 26844 11082
rect 26792 11018 26844 11024
rect 26804 10674 26832 11018
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26068 9897 26096 9998
rect 26054 9888 26110 9897
rect 26054 9823 26110 9832
rect 26712 9518 26740 9998
rect 26700 9512 26752 9518
rect 26238 9480 26294 9489
rect 26700 9454 26752 9460
rect 26238 9415 26294 9424
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25792 8090 25820 8366
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25976 7993 26004 9114
rect 25962 7984 26018 7993
rect 25872 7948 25924 7954
rect 25962 7919 26018 7928
rect 25872 7890 25924 7896
rect 25504 7880 25556 7886
rect 25884 7857 25912 7890
rect 25504 7822 25556 7828
rect 25870 7848 25926 7857
rect 25004 7296 25176 7324
rect 25240 7398 25452 7426
rect 25516 7410 25544 7822
rect 25870 7783 25926 7792
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 25504 7404 25556 7410
rect 25240 7313 25268 7398
rect 25504 7346 25556 7352
rect 25226 7304 25282 7313
rect 24952 7278 25004 7284
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24412 6089 24440 6190
rect 24398 6080 24454 6089
rect 24398 6015 24454 6024
rect 24214 5944 24270 5953
rect 24504 5914 24532 6802
rect 24688 6662 24716 7278
rect 24964 6934 24992 7278
rect 25226 7239 25282 7248
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24780 6322 24808 6666
rect 25148 6390 25176 6734
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 25148 6254 25176 6326
rect 24676 6248 24728 6254
rect 24952 6248 25004 6254
rect 24676 6190 24728 6196
rect 24950 6216 24952 6225
rect 25136 6248 25188 6254
rect 25004 6216 25006 6225
rect 24214 5879 24270 5888
rect 24492 5908 24544 5914
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22836 5160 22888 5166
rect 22388 4865 22416 5102
rect 22480 5086 22600 5114
rect 22836 5102 22888 5108
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22374 4856 22430 4865
rect 22374 4791 22430 4800
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22480 4214 22508 4966
rect 22572 4758 22600 5086
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22848 4690 22876 5102
rect 23032 4826 23060 5238
rect 23124 4826 23152 5510
rect 23216 5098 23244 5646
rect 23308 5234 23336 5646
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23400 5098 23428 5766
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23204 5092 23256 5098
rect 23204 5034 23256 5040
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23584 4826 23612 5510
rect 24228 5370 24256 5879
rect 24492 5850 24544 5856
rect 24308 5704 24360 5710
rect 24306 5672 24308 5681
rect 24584 5704 24636 5710
rect 24360 5672 24362 5681
rect 24584 5646 24636 5652
rect 24306 5607 24362 5616
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 23938 5128 23994 5137
rect 23860 5098 23938 5114
rect 23848 5092 23938 5098
rect 23900 5086 23938 5092
rect 24412 5098 24440 5238
rect 23938 5063 23994 5072
rect 24400 5092 24452 5098
rect 23848 5034 23900 5040
rect 24400 5034 24452 5040
rect 23940 5024 23992 5030
rect 23992 4984 24256 5012
rect 23940 4966 23992 4972
rect 23720 4924 24028 4933
rect 23720 4922 23726 4924
rect 23782 4922 23806 4924
rect 23862 4922 23886 4924
rect 23942 4922 23966 4924
rect 24022 4922 24028 4924
rect 23782 4870 23784 4922
rect 23964 4870 23966 4922
rect 23720 4868 23726 4870
rect 23782 4868 23806 4870
rect 23862 4868 23886 4870
rect 23942 4868 23966 4870
rect 24022 4868 24028 4870
rect 23720 4859 24028 4868
rect 24228 4826 24256 4984
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 23478 4720 23534 4729
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22928 4684 22980 4690
rect 23478 4655 23534 4664
rect 22928 4626 22980 4632
rect 22940 4282 22968 4626
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 21970 3998 22048 4026
rect 21914 3975 21970 3984
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3738 21864 3878
rect 22020 3738 22048 3998
rect 22112 3998 22232 4026
rect 21732 3732 21784 3738
rect 21732 3674 21784 3680
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 21744 3097 21772 3674
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21928 3482 21956 3538
rect 21836 3126 21864 3470
rect 21928 3466 22048 3482
rect 21928 3460 22060 3466
rect 21928 3454 22008 3460
rect 22008 3402 22060 3408
rect 22112 3194 22140 3998
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21824 3120 21876 3126
rect 21730 3088 21786 3097
rect 21824 3062 21876 3068
rect 21730 3023 21732 3032
rect 21784 3023 21786 3032
rect 21732 2994 21784 3000
rect 21272 2916 21496 2922
rect 21324 2910 21496 2916
rect 21652 2910 21772 2938
rect 21272 2858 21324 2864
rect 21456 2848 21508 2854
rect 21508 2796 21680 2802
rect 21456 2790 21680 2796
rect 21468 2774 21680 2790
rect 20916 2746 21036 2774
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18144 2100 18196 2106
rect 18144 2042 18196 2048
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 18984 1766 19012 2246
rect 19064 1964 19116 1970
rect 19064 1906 19116 1912
rect 15752 1760 15804 1766
rect 15752 1702 15804 1708
rect 18972 1760 19024 1766
rect 18972 1702 19024 1708
rect 15946 1660 16254 1669
rect 15946 1658 15952 1660
rect 16008 1658 16032 1660
rect 16088 1658 16112 1660
rect 16168 1658 16192 1660
rect 16248 1658 16254 1660
rect 16008 1606 16010 1658
rect 16190 1606 16192 1658
rect 15946 1604 15952 1606
rect 16008 1604 16032 1606
rect 16088 1604 16112 1606
rect 16168 1604 16192 1606
rect 16248 1604 16254 1606
rect 15946 1595 16254 1604
rect 14188 1488 14240 1494
rect 14188 1430 14240 1436
rect 19076 1358 19104 1906
rect 19156 1760 19208 1766
rect 19156 1702 19208 1708
rect 19168 1426 19196 1702
rect 19260 1562 19288 2450
rect 20352 2440 20404 2446
rect 19628 2378 19840 2394
rect 20352 2382 20404 2388
rect 19628 2372 19852 2378
rect 19628 2366 19800 2372
rect 19340 2100 19392 2106
rect 19340 2042 19392 2048
rect 19352 1562 19380 2042
rect 19628 2038 19656 2366
rect 19800 2314 19852 2320
rect 19833 2204 20141 2213
rect 19833 2202 19839 2204
rect 19895 2202 19919 2204
rect 19975 2202 19999 2204
rect 20055 2202 20079 2204
rect 20135 2202 20141 2204
rect 19895 2150 19897 2202
rect 20077 2150 20079 2202
rect 19833 2148 19839 2150
rect 19895 2148 19919 2150
rect 19975 2148 19999 2150
rect 20055 2148 20079 2150
rect 20135 2148 20141 2150
rect 19833 2139 20141 2148
rect 19616 2032 19668 2038
rect 19616 1974 19668 1980
rect 20364 1902 20392 2382
rect 20916 2106 20944 2518
rect 21008 2514 21036 2746
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 21284 2106 21312 2450
rect 20904 2100 20956 2106
rect 20904 2042 20956 2048
rect 21272 2100 21324 2106
rect 21272 2042 21324 2048
rect 19708 1896 19760 1902
rect 19708 1838 19760 1844
rect 20352 1896 20404 1902
rect 20352 1838 20404 1844
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 19248 1556 19300 1562
rect 19248 1498 19300 1504
rect 19340 1556 19392 1562
rect 19340 1498 19392 1504
rect 19720 1426 19748 1838
rect 20444 1828 20496 1834
rect 20444 1770 20496 1776
rect 20456 1562 20484 1770
rect 20824 1766 20852 1838
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 21376 1562 21404 2586
rect 21548 2576 21600 2582
rect 21652 2564 21680 2774
rect 21600 2536 21680 2564
rect 21548 2518 21600 2524
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21468 1986 21496 2382
rect 21468 1958 21588 1986
rect 21560 1902 21588 1958
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 21744 1834 21772 2910
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 21732 1828 21784 1834
rect 21732 1770 21784 1776
rect 20444 1556 20496 1562
rect 20444 1498 20496 1504
rect 21364 1556 21416 1562
rect 21364 1498 21416 1504
rect 21836 1494 21864 2246
rect 21928 1970 21956 2586
rect 22020 2514 22048 2790
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22112 2378 22140 2858
rect 22296 2774 22324 3878
rect 22940 3602 22968 4218
rect 23216 4214 23244 4490
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23204 4208 23256 4214
rect 23204 4150 23256 4156
rect 23018 4040 23074 4049
rect 23018 3975 23074 3984
rect 23032 3942 23060 3975
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23216 3738 23244 4150
rect 23296 4072 23348 4078
rect 23294 4040 23296 4049
rect 23348 4040 23350 4049
rect 23294 3975 23350 3984
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22204 2746 22324 2774
rect 22204 2514 22232 2746
rect 22388 2650 22416 2858
rect 22940 2774 22968 3538
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 3194 23152 3334
rect 23308 3194 23336 3470
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23032 2938 23060 3130
rect 23400 2990 23428 4422
rect 23492 4214 23520 4655
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23860 4128 23888 4422
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 23768 4100 23888 4128
rect 23768 3942 23796 4100
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23584 3618 23612 3878
rect 23720 3836 24028 3845
rect 23720 3834 23726 3836
rect 23782 3834 23806 3836
rect 23862 3834 23886 3836
rect 23942 3834 23966 3836
rect 24022 3834 24028 3836
rect 23782 3782 23784 3834
rect 23964 3782 23966 3834
rect 23720 3780 23726 3782
rect 23782 3780 23806 3782
rect 23862 3780 23886 3782
rect 23942 3780 23966 3782
rect 24022 3780 24028 3782
rect 23720 3771 24028 3780
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23584 3590 23796 3618
rect 23664 3528 23716 3534
rect 23492 3488 23664 3516
rect 23204 2984 23256 2990
rect 23032 2932 23204 2938
rect 23032 2926 23256 2932
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23032 2910 23244 2926
rect 22940 2746 23428 2774
rect 23400 2650 23428 2746
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 23492 2378 23520 3488
rect 23664 3470 23716 3476
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23584 2514 23612 3334
rect 23768 3126 23796 3590
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 23860 2990 23888 3674
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 24044 3505 24072 3538
rect 24030 3496 24086 3505
rect 24030 3431 24086 3440
rect 24136 3194 24164 4218
rect 24412 4185 24440 4762
rect 24504 4690 24532 5510
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24398 4176 24454 4185
rect 24398 4111 24454 4120
rect 24412 3670 24440 4111
rect 24400 3664 24452 3670
rect 24596 3652 24624 5646
rect 24688 4214 24716 6190
rect 25136 6190 25188 6196
rect 24950 6151 25006 6160
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25148 5914 25176 6054
rect 25240 5914 25268 7142
rect 25332 6254 25360 7210
rect 25412 6928 25464 6934
rect 25412 6870 25464 6876
rect 25424 6633 25452 6870
rect 25516 6798 25544 7346
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25608 7002 25636 7142
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25594 6760 25650 6769
rect 25594 6695 25650 6704
rect 25410 6624 25466 6633
rect 25410 6559 25466 6568
rect 25502 6352 25558 6361
rect 25502 6287 25558 6296
rect 25320 6248 25372 6254
rect 25372 6208 25452 6236
rect 25320 6190 25372 6196
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 24858 5808 24914 5817
rect 24858 5743 24860 5752
rect 24912 5743 24914 5752
rect 24860 5714 24912 5720
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24964 5370 24992 5646
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24780 4593 24808 5238
rect 24766 4584 24822 4593
rect 24822 4542 24992 4570
rect 24766 4519 24822 4528
rect 24676 4208 24728 4214
rect 24676 4150 24728 4156
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24400 3606 24452 3612
rect 24504 3624 24624 3652
rect 24504 3398 24532 3624
rect 24676 3596 24728 3602
rect 24596 3556 24676 3584
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24216 3052 24268 3058
rect 23952 3012 24216 3040
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23952 2922 23980 3012
rect 24268 3012 24440 3040
rect 24216 2994 24268 3000
rect 23940 2916 23992 2922
rect 23940 2858 23992 2864
rect 24216 2916 24268 2922
rect 24216 2858 24268 2864
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 23720 2748 24028 2757
rect 23720 2746 23726 2748
rect 23782 2746 23806 2748
rect 23862 2746 23886 2748
rect 23942 2746 23966 2748
rect 24022 2746 24028 2748
rect 23782 2694 23784 2746
rect 23964 2694 23966 2746
rect 23720 2692 23726 2694
rect 23782 2692 23806 2694
rect 23862 2692 23886 2694
rect 23942 2692 23966 2694
rect 24022 2692 24028 2694
rect 23720 2683 24028 2692
rect 24136 2632 24164 2790
rect 24044 2604 24164 2632
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 24044 2446 24072 2604
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24228 2378 24256 2858
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 24216 2372 24268 2378
rect 24216 2314 24268 2320
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 22296 2106 22324 2246
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 23492 2038 23520 2314
rect 24320 2310 24348 2450
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 23768 2106 23796 2246
rect 24412 2106 24440 3012
rect 24596 2514 24624 3556
rect 24676 3538 24728 3544
rect 24674 3088 24730 3097
rect 24674 3023 24676 3032
rect 24728 3023 24730 3032
rect 24676 2994 24728 3000
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24596 2106 24624 2450
rect 24688 2428 24716 2858
rect 24780 2582 24808 3878
rect 24872 3670 24900 4014
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24964 3482 24992 4542
rect 25056 4049 25084 5510
rect 25148 5250 25176 5850
rect 25240 5778 25268 5850
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25226 5264 25282 5273
rect 25148 5222 25226 5250
rect 25148 4826 25176 5222
rect 25226 5199 25282 5208
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 4078 25176 4626
rect 25136 4072 25188 4078
rect 25042 4040 25098 4049
rect 25136 4014 25188 4020
rect 25042 3975 25098 3984
rect 24872 3454 24992 3482
rect 24872 3369 24900 3454
rect 24952 3392 25004 3398
rect 24858 3360 24914 3369
rect 24952 3334 25004 3340
rect 24858 3295 24914 3304
rect 24872 3194 24900 3295
rect 24964 3194 24992 3334
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 24964 2582 24992 2926
rect 25056 2922 25084 3975
rect 25134 3768 25190 3777
rect 25134 3703 25190 3712
rect 25148 3602 25176 3703
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25240 3505 25268 4694
rect 25332 4622 25360 6054
rect 25424 5166 25452 6208
rect 25516 5760 25544 6287
rect 25608 6254 25636 6695
rect 25700 6497 25728 7142
rect 25686 6488 25742 6497
rect 25686 6423 25742 6432
rect 25792 6254 25820 7414
rect 25872 6792 25924 6798
rect 25976 6746 26004 7919
rect 25924 6740 26004 6746
rect 25872 6734 26004 6740
rect 25884 6718 26004 6734
rect 26068 6644 26096 9318
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26160 8634 26188 8910
rect 26252 8634 26280 9415
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26344 7478 26372 9318
rect 26436 9178 26464 9318
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26516 7948 26568 7954
rect 26620 7936 26648 8842
rect 26712 8362 26740 9454
rect 27172 9450 27200 14334
rect 27264 13258 27292 16594
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27264 12442 27292 13194
rect 27356 12986 27384 18226
rect 27448 17134 27476 19382
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27448 16794 27476 17070
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27540 16114 27568 21422
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27896 21004 27948 21010
rect 27948 20964 28028 20992
rect 27896 20946 27948 20952
rect 27816 20806 27844 20946
rect 27804 20800 27856 20806
rect 27804 20742 27856 20748
rect 27607 20700 27915 20709
rect 27607 20698 27613 20700
rect 27669 20698 27693 20700
rect 27749 20698 27773 20700
rect 27829 20698 27853 20700
rect 27909 20698 27915 20700
rect 27669 20646 27671 20698
rect 27851 20646 27853 20698
rect 27607 20644 27613 20646
rect 27669 20644 27693 20646
rect 27749 20644 27773 20646
rect 27829 20644 27853 20646
rect 27909 20644 27915 20646
rect 27607 20635 27915 20644
rect 27607 19612 27915 19621
rect 27607 19610 27613 19612
rect 27669 19610 27693 19612
rect 27749 19610 27773 19612
rect 27829 19610 27853 19612
rect 27909 19610 27915 19612
rect 27669 19558 27671 19610
rect 27851 19558 27853 19610
rect 27607 19556 27613 19558
rect 27669 19556 27693 19558
rect 27749 19556 27773 19558
rect 27829 19556 27853 19558
rect 27909 19556 27915 19558
rect 27607 19547 27915 19556
rect 27607 18524 27915 18533
rect 27607 18522 27613 18524
rect 27669 18522 27693 18524
rect 27749 18522 27773 18524
rect 27829 18522 27853 18524
rect 27909 18522 27915 18524
rect 27669 18470 27671 18522
rect 27851 18470 27853 18522
rect 27607 18468 27613 18470
rect 27669 18468 27693 18470
rect 27749 18468 27773 18470
rect 27829 18468 27853 18470
rect 27909 18468 27915 18470
rect 27607 18459 27915 18468
rect 27802 18320 27858 18329
rect 27802 18255 27858 18264
rect 27816 18154 27844 18255
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27607 17436 27915 17445
rect 27607 17434 27613 17436
rect 27669 17434 27693 17436
rect 27749 17434 27773 17436
rect 27829 17434 27853 17436
rect 27909 17434 27915 17436
rect 27669 17382 27671 17434
rect 27851 17382 27853 17434
rect 27607 17380 27613 17382
rect 27669 17380 27693 17382
rect 27749 17380 27773 17382
rect 27829 17380 27853 17382
rect 27909 17380 27915 17382
rect 27607 17371 27915 17380
rect 28000 17338 28028 20964
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28092 19922 28120 20742
rect 28368 20262 28396 20878
rect 28460 20466 28488 21626
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28356 20256 28408 20262
rect 28356 20198 28408 20204
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 28552 19786 28580 20946
rect 28632 20392 28684 20398
rect 28828 20346 28856 21490
rect 29748 21486 29776 21927
rect 30010 21856 30066 21865
rect 30010 21791 30066 21800
rect 30286 21856 30342 21865
rect 30286 21791 30342 21800
rect 30024 21486 30052 21791
rect 30300 21486 30328 21791
rect 29000 21480 29052 21486
rect 29184 21480 29236 21486
rect 29052 21428 29132 21434
rect 29000 21422 29132 21428
rect 29184 21422 29236 21428
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 30288 21480 30340 21486
rect 30288 21422 30340 21428
rect 29012 21406 29132 21422
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 28632 20334 28684 20340
rect 28080 19780 28132 19786
rect 28080 19722 28132 19728
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28092 18358 28120 19722
rect 28644 19156 28672 20334
rect 28736 20318 28856 20346
rect 28736 20210 28764 20318
rect 28736 20182 28856 20210
rect 28552 19128 28672 19156
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 28080 18352 28132 18358
rect 28080 18294 28132 18300
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 27988 17332 28040 17338
rect 27988 17274 28040 17280
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27632 16522 27660 17070
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27607 16348 27915 16357
rect 27607 16346 27613 16348
rect 27669 16346 27693 16348
rect 27749 16346 27773 16348
rect 27829 16346 27853 16348
rect 27909 16346 27915 16348
rect 27669 16294 27671 16346
rect 27851 16294 27853 16346
rect 27607 16292 27613 16294
rect 27669 16292 27693 16294
rect 27749 16292 27773 16294
rect 27829 16292 27853 16294
rect 27909 16292 27915 16294
rect 27607 16283 27915 16292
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27436 15972 27488 15978
rect 27436 15914 27488 15920
rect 27448 15570 27476 15914
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27540 15706 27568 15846
rect 27710 15736 27766 15745
rect 27528 15700 27580 15706
rect 27710 15671 27766 15680
rect 27528 15642 27580 15648
rect 27724 15638 27752 15671
rect 27712 15632 27764 15638
rect 27712 15574 27764 15580
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27988 15564 28040 15570
rect 28092 15552 28120 17818
rect 28184 16114 28212 18566
rect 28354 18184 28410 18193
rect 28354 18119 28410 18128
rect 28368 17746 28396 18119
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28264 17264 28316 17270
rect 28264 17206 28316 17212
rect 28276 16658 28304 17206
rect 28368 17066 28396 17682
rect 28356 17060 28408 17066
rect 28356 17002 28408 17008
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28040 15524 28120 15552
rect 28264 15564 28316 15570
rect 27988 15506 28040 15512
rect 28264 15506 28316 15512
rect 27540 15162 27568 15506
rect 27607 15260 27915 15269
rect 27607 15258 27613 15260
rect 27669 15258 27693 15260
rect 27749 15258 27773 15260
rect 27829 15258 27853 15260
rect 27909 15258 27915 15260
rect 27669 15206 27671 15258
rect 27851 15206 27853 15258
rect 27607 15204 27613 15206
rect 27669 15204 27693 15206
rect 27749 15204 27773 15206
rect 27829 15204 27853 15206
rect 27909 15204 27915 15206
rect 27607 15195 27915 15204
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 28000 15026 28028 15506
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28080 14884 28132 14890
rect 28080 14826 28132 14832
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 27448 14074 27476 14486
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27607 14172 27915 14181
rect 27607 14170 27613 14172
rect 27669 14170 27693 14172
rect 27749 14170 27773 14172
rect 27829 14170 27853 14172
rect 27909 14170 27915 14172
rect 27669 14118 27671 14170
rect 27851 14118 27853 14170
rect 27607 14116 27613 14118
rect 27669 14116 27693 14118
rect 27749 14116 27773 14118
rect 27829 14116 27853 14118
rect 27909 14116 27915 14118
rect 27607 14107 27915 14116
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27712 13456 27764 13462
rect 27434 13424 27490 13433
rect 27712 13398 27764 13404
rect 27434 13359 27436 13368
rect 27488 13359 27490 13368
rect 27436 13330 27488 13336
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27448 12782 27476 13330
rect 27724 13326 27752 13398
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27607 13084 27915 13093
rect 27607 13082 27613 13084
rect 27669 13082 27693 13084
rect 27749 13082 27773 13084
rect 27829 13082 27853 13084
rect 27909 13082 27915 13084
rect 27669 13030 27671 13082
rect 27851 13030 27853 13082
rect 27607 13028 27613 13030
rect 27669 13028 27693 13030
rect 27749 13028 27773 13030
rect 27829 13028 27853 13030
rect 27909 13028 27915 13030
rect 27607 13019 27915 13028
rect 28000 12986 28028 14214
rect 28092 13462 28120 14826
rect 28080 13456 28132 13462
rect 28080 13398 28132 13404
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 28184 12918 28212 15098
rect 28276 14618 28304 15506
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28172 12912 28224 12918
rect 27526 12880 27582 12889
rect 28172 12854 28224 12860
rect 27526 12815 27528 12824
rect 27580 12815 27582 12824
rect 27528 12786 27580 12792
rect 28276 12782 28304 13874
rect 28368 13802 28396 16390
rect 28460 14906 28488 17750
rect 28552 17678 28580 19128
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28552 16776 28580 17614
rect 28644 17610 28672 18158
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28644 17202 28672 17546
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28552 16748 28672 16776
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28552 15366 28580 16594
rect 28644 16182 28672 16748
rect 28736 16697 28764 17682
rect 28722 16688 28778 16697
rect 28722 16623 28778 16632
rect 28828 16522 28856 20182
rect 29012 19310 29040 21286
rect 29104 21078 29132 21406
rect 29196 21146 29224 21422
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 29368 21344 29420 21350
rect 29368 21286 29420 21292
rect 29184 21140 29236 21146
rect 29184 21082 29236 21088
rect 29092 21072 29144 21078
rect 29092 21014 29144 21020
rect 29104 20602 29132 21014
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29184 20324 29236 20330
rect 29184 20266 29236 20272
rect 29196 20058 29224 20266
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 29000 19304 29052 19310
rect 28906 19272 28962 19281
rect 29000 19246 29052 19252
rect 28906 19207 28962 19216
rect 28920 18834 28948 19207
rect 29104 18986 29132 19382
rect 29380 19310 29408 21286
rect 29460 20596 29512 20602
rect 29460 20538 29512 20544
rect 29472 20058 29500 20538
rect 29552 20324 29604 20330
rect 29552 20266 29604 20272
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29012 18958 29132 18986
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28920 17882 28948 18566
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 28920 16522 28948 17138
rect 28816 16516 28868 16522
rect 28816 16458 28868 16464
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28460 14878 28580 14906
rect 28448 14816 28500 14822
rect 28448 14758 28500 14764
rect 28460 14385 28488 14758
rect 28552 14482 28580 14878
rect 28540 14476 28592 14482
rect 28540 14418 28592 14424
rect 28446 14376 28502 14385
rect 28446 14311 28502 14320
rect 28644 13938 28672 15506
rect 28736 14482 28764 15982
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28630 13832 28686 13841
rect 28356 13796 28408 13802
rect 28630 13767 28686 13776
rect 28356 13738 28408 13744
rect 28368 13462 28396 13738
rect 28356 13456 28408 13462
rect 28356 13398 28408 13404
rect 28644 13258 28672 13767
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 28264 12776 28316 12782
rect 28264 12718 28316 12724
rect 27252 12436 27304 12442
rect 29012 12434 29040 18958
rect 29196 18873 29224 19246
rect 29288 18970 29316 19246
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29182 18864 29238 18873
rect 29092 18828 29144 18834
rect 29182 18799 29238 18808
rect 29092 18770 29144 18776
rect 29104 17202 29132 18770
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 29184 17808 29236 17814
rect 29184 17750 29236 17756
rect 29196 17270 29224 17750
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29196 16658 29224 17206
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 29288 16454 29316 18362
rect 29472 17542 29500 19450
rect 29564 18426 29592 20266
rect 29656 19310 29684 21354
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 30300 20777 30328 21286
rect 30286 20768 30342 20777
rect 30286 20703 30342 20712
rect 29734 20496 29790 20505
rect 29734 20431 29790 20440
rect 30196 20460 30248 20466
rect 29748 19990 29776 20431
rect 30196 20402 30248 20408
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29932 19514 29960 20334
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29380 16658 29408 17070
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29276 16448 29328 16454
rect 29276 16390 29328 16396
rect 29380 16250 29408 16594
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29380 15162 29408 15506
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 29104 13394 29132 14418
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29472 13190 29500 17478
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29564 15706 29592 16594
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29656 15570 29684 16186
rect 29736 15972 29788 15978
rect 29736 15914 29788 15920
rect 29748 15609 29776 15914
rect 29734 15600 29790 15609
rect 29644 15564 29696 15570
rect 29734 15535 29736 15544
rect 29644 15506 29696 15512
rect 29788 15535 29790 15544
rect 29736 15506 29788 15512
rect 29656 14482 29684 15506
rect 29840 15502 29868 19246
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29932 17882 29960 18702
rect 30116 18222 30144 20198
rect 30208 19310 30236 20402
rect 30392 20346 30420 21966
rect 30840 21888 30892 21894
rect 30840 21830 30892 21836
rect 30852 21146 30880 21830
rect 31494 21244 31802 21253
rect 31494 21242 31500 21244
rect 31556 21242 31580 21244
rect 31636 21242 31660 21244
rect 31716 21242 31740 21244
rect 31796 21242 31802 21244
rect 31556 21190 31558 21242
rect 31738 21190 31740 21242
rect 31494 21188 31500 21190
rect 31556 21188 31580 21190
rect 31636 21188 31660 21190
rect 31716 21188 31740 21190
rect 31796 21188 31802 21190
rect 31494 21179 31802 21188
rect 30840 21140 30892 21146
rect 30840 21082 30892 21088
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30484 20602 30512 20742
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 30576 20534 30604 20878
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30852 20466 30880 21082
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30748 20392 30800 20398
rect 30288 20324 30340 20330
rect 30392 20318 30512 20346
rect 30748 20334 30800 20340
rect 30288 20266 30340 20272
rect 30300 19446 30328 20266
rect 30484 19922 30512 20318
rect 30760 20074 30788 20334
rect 30760 20058 30880 20074
rect 30748 20052 30880 20058
rect 30800 20046 30880 20052
rect 30748 19994 30800 20000
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30208 18426 30236 19246
rect 30484 18426 30512 19858
rect 30656 19304 30708 19310
rect 30576 19264 30656 19292
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30012 18148 30064 18154
rect 30012 18090 30064 18096
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 14618 29868 15438
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 30024 14482 30052 18090
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30194 17912 30250 17921
rect 30194 17847 30250 17856
rect 30208 17746 30236 17847
rect 30484 17746 30512 18022
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30196 16992 30248 16998
rect 30196 16934 30248 16940
rect 30208 16250 30236 16934
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 30208 15570 30236 16050
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30208 15162 30236 15506
rect 30196 15156 30248 15162
rect 30196 15098 30248 15104
rect 30104 14612 30156 14618
rect 30104 14554 30156 14560
rect 30116 14521 30144 14554
rect 30102 14512 30158 14521
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 30012 14476 30064 14482
rect 30102 14447 30158 14456
rect 30012 14418 30064 14424
rect 30116 14414 30144 14447
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29828 14272 29880 14278
rect 29828 14214 29880 14220
rect 29840 13394 29868 14214
rect 30208 13870 30236 15098
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29460 13184 29512 13190
rect 29460 13126 29512 13132
rect 29840 12986 29868 13330
rect 30300 12986 30328 17546
rect 30472 17196 30524 17202
rect 30472 17138 30524 17144
rect 30380 17060 30432 17066
rect 30380 17002 30432 17008
rect 30392 16658 30420 17002
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30392 15638 30420 15982
rect 30484 15910 30512 17138
rect 30576 16998 30604 19264
rect 30656 19246 30708 19252
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30668 18970 30696 19110
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30656 18216 30708 18222
rect 30656 18158 30708 18164
rect 30668 17338 30696 18158
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30576 16794 30604 16934
rect 30564 16788 30616 16794
rect 30564 16730 30616 16736
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30380 15632 30432 15638
rect 30380 15574 30432 15580
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30392 14550 30420 15438
rect 30484 14890 30512 15846
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30576 14958 30604 15506
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30472 14884 30524 14890
rect 30472 14826 30524 14832
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13870 30420 14214
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30392 12782 30420 13806
rect 30484 13530 30512 14554
rect 30576 14074 30604 14894
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30668 12986 30696 16594
rect 30760 16046 30788 19858
rect 30852 19378 30880 20046
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30840 17264 30892 17270
rect 30840 17206 30892 17212
rect 30748 16040 30800 16046
rect 30748 15982 30800 15988
rect 30852 15162 30880 17206
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30852 14482 30880 15098
rect 30944 14618 30972 20946
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 31036 19990 31064 20334
rect 31494 20156 31802 20165
rect 31494 20154 31500 20156
rect 31556 20154 31580 20156
rect 31636 20154 31660 20156
rect 31716 20154 31740 20156
rect 31796 20154 31802 20156
rect 31556 20102 31558 20154
rect 31738 20102 31740 20154
rect 31494 20100 31500 20102
rect 31556 20100 31580 20102
rect 31636 20100 31660 20102
rect 31716 20100 31740 20102
rect 31796 20100 31802 20102
rect 31494 20091 31802 20100
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 31036 14482 31064 19314
rect 31494 19068 31802 19077
rect 31494 19066 31500 19068
rect 31556 19066 31580 19068
rect 31636 19066 31660 19068
rect 31716 19066 31740 19068
rect 31796 19066 31802 19068
rect 31556 19014 31558 19066
rect 31738 19014 31740 19066
rect 31494 19012 31500 19014
rect 31556 19012 31580 19014
rect 31636 19012 31660 19014
rect 31716 19012 31740 19014
rect 31796 19012 31802 19014
rect 31494 19003 31802 19012
rect 31494 17980 31802 17989
rect 31494 17978 31500 17980
rect 31556 17978 31580 17980
rect 31636 17978 31660 17980
rect 31716 17978 31740 17980
rect 31796 17978 31802 17980
rect 31556 17926 31558 17978
rect 31738 17926 31740 17978
rect 31494 17924 31500 17926
rect 31556 17924 31580 17926
rect 31636 17924 31660 17926
rect 31716 17924 31740 17926
rect 31796 17924 31802 17926
rect 31494 17915 31802 17924
rect 31494 16892 31802 16901
rect 31494 16890 31500 16892
rect 31556 16890 31580 16892
rect 31636 16890 31660 16892
rect 31716 16890 31740 16892
rect 31796 16890 31802 16892
rect 31556 16838 31558 16890
rect 31738 16838 31740 16890
rect 31494 16836 31500 16838
rect 31556 16836 31580 16838
rect 31636 16836 31660 16838
rect 31716 16836 31740 16838
rect 31796 16836 31802 16838
rect 31494 16827 31802 16836
rect 31494 15804 31802 15813
rect 31494 15802 31500 15804
rect 31556 15802 31580 15804
rect 31636 15802 31660 15804
rect 31716 15802 31740 15804
rect 31796 15802 31802 15804
rect 31556 15750 31558 15802
rect 31738 15750 31740 15802
rect 31494 15748 31500 15750
rect 31556 15748 31580 15750
rect 31636 15748 31660 15750
rect 31716 15748 31740 15750
rect 31796 15748 31802 15750
rect 31494 15739 31802 15748
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31128 14618 31156 14962
rect 31494 14716 31802 14725
rect 31494 14714 31500 14716
rect 31556 14714 31580 14716
rect 31636 14714 31660 14716
rect 31716 14714 31740 14716
rect 31796 14714 31802 14716
rect 31556 14662 31558 14714
rect 31738 14662 31740 14714
rect 31494 14660 31500 14662
rect 31556 14660 31580 14662
rect 31636 14660 31660 14662
rect 31716 14660 31740 14662
rect 31796 14660 31802 14662
rect 31494 14651 31802 14660
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 30852 13530 30880 14418
rect 31036 13530 31064 14418
rect 31494 13628 31802 13637
rect 31494 13626 31500 13628
rect 31556 13626 31580 13628
rect 31636 13626 31660 13628
rect 31716 13626 31740 13628
rect 31796 13626 31802 13628
rect 31556 13574 31558 13626
rect 31738 13574 31740 13626
rect 31494 13572 31500 13574
rect 31556 13572 31580 13574
rect 31636 13572 31660 13574
rect 31716 13572 31740 13574
rect 31796 13572 31802 13574
rect 31494 13563 31802 13572
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 31494 12540 31802 12549
rect 31494 12538 31500 12540
rect 31556 12538 31580 12540
rect 31636 12538 31660 12540
rect 31716 12538 31740 12540
rect 31796 12538 31802 12540
rect 31556 12486 31558 12538
rect 31738 12486 31740 12538
rect 31494 12484 31500 12486
rect 31556 12484 31580 12486
rect 31636 12484 31660 12486
rect 31716 12484 31740 12486
rect 31796 12484 31802 12486
rect 31494 12475 31802 12484
rect 27252 12378 27304 12384
rect 28920 12406 29040 12434
rect 27607 11996 27915 12005
rect 27607 11994 27613 11996
rect 27669 11994 27693 11996
rect 27749 11994 27773 11996
rect 27829 11994 27853 11996
rect 27909 11994 27915 11996
rect 27669 11942 27671 11994
rect 27851 11942 27853 11994
rect 27607 11940 27613 11942
rect 27669 11940 27693 11942
rect 27749 11940 27773 11942
rect 27829 11940 27853 11942
rect 27909 11940 27915 11942
rect 27607 11931 27915 11940
rect 27528 11552 27580 11558
rect 27528 11494 27580 11500
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 27540 10538 27568 11494
rect 28644 11218 28672 11494
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 27607 10908 27915 10917
rect 27607 10906 27613 10908
rect 27669 10906 27693 10908
rect 27749 10906 27773 10908
rect 27829 10906 27853 10908
rect 27909 10906 27915 10908
rect 27669 10854 27671 10906
rect 27851 10854 27853 10906
rect 27607 10852 27613 10854
rect 27669 10852 27693 10854
rect 27749 10852 27773 10854
rect 27829 10852 27853 10854
rect 27909 10852 27915 10854
rect 27607 10843 27915 10852
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27712 10532 27764 10538
rect 27712 10474 27764 10480
rect 27540 10146 27568 10474
rect 27724 10266 27752 10474
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27448 10118 27568 10146
rect 27618 10160 27674 10169
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26804 8838 26832 9318
rect 27448 9110 27476 10118
rect 27618 10095 27674 10104
rect 27632 10062 27660 10095
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27607 9820 27915 9829
rect 27607 9818 27613 9820
rect 27669 9818 27693 9820
rect 27749 9818 27773 9820
rect 27829 9818 27853 9820
rect 27909 9818 27915 9820
rect 27669 9766 27671 9818
rect 27851 9766 27853 9818
rect 27607 9764 27613 9766
rect 27669 9764 27693 9766
rect 27749 9764 27773 9766
rect 27829 9764 27853 9766
rect 27909 9764 27915 9766
rect 27607 9755 27915 9764
rect 27802 9616 27858 9625
rect 28184 9586 28212 11086
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28828 10198 28856 10542
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 28920 9586 28948 12406
rect 29734 12200 29790 12209
rect 29734 12135 29790 12144
rect 29748 11354 29776 12135
rect 29918 11792 29974 11801
rect 29918 11727 29974 11736
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29932 11218 29960 11727
rect 31494 11452 31802 11461
rect 31494 11450 31500 11452
rect 31556 11450 31580 11452
rect 31636 11450 31660 11452
rect 31716 11450 31740 11452
rect 31796 11450 31802 11452
rect 31556 11398 31558 11450
rect 31738 11398 31740 11450
rect 31494 11396 31500 11398
rect 31556 11396 31580 11398
rect 31636 11396 31660 11398
rect 31716 11396 31740 11398
rect 31796 11396 31802 11398
rect 31494 11387 31802 11396
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 30196 11008 30248 11014
rect 30196 10950 30248 10956
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29000 10532 29052 10538
rect 29000 10474 29052 10480
rect 29012 10266 29040 10474
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 27802 9551 27858 9560
rect 28172 9580 28224 9586
rect 27816 9382 27844 9551
rect 28172 9522 28224 9528
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 27436 9104 27488 9110
rect 27436 9046 27488 9052
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 27540 8634 27568 9318
rect 28368 9178 28396 9318
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 29104 9110 29132 10542
rect 29564 10198 29592 10950
rect 30208 10606 30236 10950
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 29552 10192 29604 10198
rect 29552 10134 29604 10140
rect 30208 9722 30236 10542
rect 31494 10364 31802 10373
rect 31494 10362 31500 10364
rect 31556 10362 31580 10364
rect 31636 10362 31660 10364
rect 31716 10362 31740 10364
rect 31796 10362 31802 10364
rect 31556 10310 31558 10362
rect 31738 10310 31740 10362
rect 31494 10308 31500 10310
rect 31556 10308 31580 10310
rect 31636 10308 31660 10310
rect 31716 10308 31740 10310
rect 31796 10308 31802 10310
rect 31494 10299 31802 10308
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 31494 9276 31802 9285
rect 31494 9274 31500 9276
rect 31556 9274 31580 9276
rect 31636 9274 31660 9276
rect 31716 9274 31740 9276
rect 31796 9274 31802 9276
rect 31556 9222 31558 9274
rect 31738 9222 31740 9274
rect 31494 9220 31500 9222
rect 31556 9220 31580 9222
rect 31636 9220 31660 9222
rect 31716 9220 31740 9222
rect 31796 9220 31802 9222
rect 31494 9211 31802 9220
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 27607 8732 27915 8741
rect 27607 8730 27613 8732
rect 27669 8730 27693 8732
rect 27749 8730 27773 8732
rect 27829 8730 27853 8732
rect 27909 8730 27915 8732
rect 27669 8678 27671 8730
rect 27851 8678 27853 8730
rect 27607 8676 27613 8678
rect 27669 8676 27693 8678
rect 27749 8676 27773 8678
rect 27829 8676 27853 8678
rect 27909 8676 27915 8678
rect 27607 8667 27915 8676
rect 28644 8634 28672 8910
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 26700 8356 26752 8362
rect 26700 8298 26752 8304
rect 26568 7908 26648 7936
rect 26516 7890 26568 7896
rect 26332 7472 26384 7478
rect 26384 7432 26464 7460
rect 26332 7414 26384 7420
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 26160 6866 26188 7142
rect 26252 6866 26280 7278
rect 26332 6996 26384 7002
rect 26332 6938 26384 6944
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 26344 6798 26372 6938
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26148 6656 26200 6662
rect 26068 6616 26148 6644
rect 26148 6598 26200 6604
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 25596 6248 25648 6254
rect 25596 6190 25648 6196
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 25608 6118 25636 6190
rect 25596 6112 25648 6118
rect 25700 6089 25728 6190
rect 25596 6054 25648 6060
rect 25686 6080 25742 6089
rect 25686 6015 25742 6024
rect 25596 5772 25648 5778
rect 25516 5732 25596 5760
rect 25596 5714 25648 5720
rect 25504 5568 25556 5574
rect 25502 5536 25504 5545
rect 25556 5536 25558 5545
rect 25502 5471 25558 5480
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 25332 4146 25360 4558
rect 25608 4554 25636 5714
rect 25792 5370 25820 6190
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25792 4729 25820 4762
rect 25778 4720 25834 4729
rect 25688 4684 25740 4690
rect 25778 4655 25834 4664
rect 25688 4626 25740 4632
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25504 4480 25556 4486
rect 25504 4422 25556 4428
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25226 3496 25282 3505
rect 25226 3431 25282 3440
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 24768 2576 24820 2582
rect 24952 2576 25004 2582
rect 24820 2536 24900 2564
rect 24768 2518 24820 2524
rect 24768 2440 24820 2446
rect 24688 2400 24768 2428
rect 24768 2382 24820 2388
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 24400 2100 24452 2106
rect 24400 2042 24452 2048
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 23480 2032 23532 2038
rect 23480 1974 23532 1980
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 24688 1714 24716 2246
rect 24780 1892 24808 2382
rect 24872 1970 24900 2536
rect 24952 2518 25004 2524
rect 25228 2508 25280 2514
rect 25332 2496 25360 2858
rect 25424 2650 25452 4422
rect 25516 4078 25544 4422
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25594 4040 25650 4049
rect 25594 3975 25596 3984
rect 25648 3975 25650 3984
rect 25596 3946 25648 3952
rect 25700 3602 25728 4626
rect 25884 4282 25912 6394
rect 25964 6384 26016 6390
rect 25964 6326 26016 6332
rect 25976 5778 26004 6326
rect 26160 5778 26188 6598
rect 26252 6458 26280 6598
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26252 5953 26280 6054
rect 26238 5944 26294 5953
rect 26238 5879 26240 5888
rect 26292 5879 26294 5888
rect 26240 5850 26292 5856
rect 25964 5772 26016 5778
rect 25964 5714 26016 5720
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 25976 5370 26004 5510
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25962 5128 26018 5137
rect 25962 5063 25964 5072
rect 26016 5063 26018 5072
rect 25964 5034 26016 5040
rect 26068 4468 26096 5510
rect 26344 4826 26372 6598
rect 26436 5914 26464 7432
rect 26528 7410 26556 7890
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 26700 7268 26752 7274
rect 26620 7228 26700 7256
rect 26620 7002 26648 7228
rect 26700 7210 26752 7216
rect 26620 6996 26692 7002
rect 26620 6944 26640 6996
rect 26620 6938 26692 6944
rect 26620 6118 26648 6938
rect 26804 6866 26832 7346
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26698 6488 26754 6497
rect 26698 6423 26754 6432
rect 26712 6254 26740 6423
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26424 5908 26476 5914
rect 26424 5850 26476 5856
rect 26422 5808 26478 5817
rect 26422 5743 26478 5752
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26344 4690 26372 4762
rect 26332 4684 26384 4690
rect 26332 4626 26384 4632
rect 26332 4548 26384 4554
rect 26436 4536 26464 5743
rect 26516 5704 26568 5710
rect 26514 5672 26516 5681
rect 26568 5672 26570 5681
rect 26712 5642 26740 6190
rect 26514 5607 26570 5616
rect 26608 5636 26660 5642
rect 26608 5578 26660 5584
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26528 5370 26556 5510
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26528 4758 26556 5306
rect 26620 5166 26648 5578
rect 26712 5370 26740 5578
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26700 5092 26752 5098
rect 26700 5034 26752 5040
rect 26516 4752 26568 4758
rect 26516 4694 26568 4700
rect 26516 4548 26568 4554
rect 26436 4508 26516 4536
rect 26332 4490 26384 4496
rect 26516 4490 26568 4496
rect 26240 4480 26292 4486
rect 26068 4440 26240 4468
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 25884 3602 25912 4218
rect 26068 3738 26096 4440
rect 26240 4422 26292 4428
rect 26344 4128 26372 4490
rect 26712 4486 26740 5034
rect 26896 4758 26924 7142
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27172 6254 27200 6598
rect 27160 6248 27212 6254
rect 27160 6190 27212 6196
rect 27344 6248 27396 6254
rect 27344 6190 27396 6196
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 26988 5778 27016 6054
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 26988 5030 27016 5714
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 27080 5545 27108 5646
rect 27066 5536 27122 5545
rect 27066 5471 27122 5480
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26884 4752 26936 4758
rect 26882 4720 26884 4729
rect 26936 4720 26938 4729
rect 26792 4684 26844 4690
rect 26882 4655 26938 4664
rect 26792 4626 26844 4632
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26424 4140 26476 4146
rect 26344 4100 26424 4128
rect 26424 4082 26476 4088
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 26528 3602 26556 4014
rect 26700 4004 26752 4010
rect 26700 3946 26752 3952
rect 26712 3738 26740 3946
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 26804 3534 26832 4626
rect 26882 4584 26938 4593
rect 26882 4519 26938 4528
rect 26896 4078 26924 4519
rect 26976 4480 27028 4486
rect 26976 4422 27028 4428
rect 26988 4078 27016 4422
rect 27080 4078 27108 5471
rect 27158 5264 27214 5273
rect 27158 5199 27214 5208
rect 27172 5030 27200 5199
rect 27356 5098 27384 6190
rect 27344 5092 27396 5098
rect 27344 5034 27396 5040
rect 27160 5024 27212 5030
rect 27212 4984 27292 5012
rect 27160 4966 27212 4972
rect 27264 4078 27292 4984
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26976 4072 27028 4078
rect 26976 4014 27028 4020
rect 27068 4072 27120 4078
rect 27160 4072 27212 4078
rect 27068 4014 27120 4020
rect 27158 4040 27160 4049
rect 27252 4072 27304 4078
rect 27212 4040 27214 4049
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26896 3466 26924 3878
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 26884 3460 26936 3466
rect 26884 3402 26936 3408
rect 25700 3194 25728 3402
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 26988 3126 27016 4014
rect 27252 4014 27304 4020
rect 27158 3975 27214 3984
rect 27448 3602 27476 8502
rect 28172 8424 28224 8430
rect 28172 8366 28224 8372
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 27607 7644 27915 7653
rect 27607 7642 27613 7644
rect 27669 7642 27693 7644
rect 27749 7642 27773 7644
rect 27829 7642 27853 7644
rect 27909 7642 27915 7644
rect 27669 7590 27671 7642
rect 27851 7590 27853 7642
rect 27607 7588 27613 7590
rect 27669 7588 27693 7590
rect 27749 7588 27773 7590
rect 27829 7588 27853 7590
rect 27909 7588 27915 7590
rect 27607 7579 27915 7588
rect 28000 7206 28028 8230
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 28092 7002 28120 7822
rect 28080 6996 28132 7002
rect 28080 6938 28132 6944
rect 27607 6556 27915 6565
rect 27607 6554 27613 6556
rect 27669 6554 27693 6556
rect 27749 6554 27773 6556
rect 27829 6554 27853 6556
rect 27909 6554 27915 6556
rect 27669 6502 27671 6554
rect 27851 6502 27853 6554
rect 27607 6500 27613 6502
rect 27669 6500 27693 6502
rect 27749 6500 27773 6502
rect 27829 6500 27853 6502
rect 27909 6500 27915 6502
rect 27607 6491 27915 6500
rect 28184 6458 28212 8366
rect 29104 8090 29132 9046
rect 31494 8188 31802 8197
rect 31494 8186 31500 8188
rect 31556 8186 31580 8188
rect 31636 8186 31660 8188
rect 31716 8186 31740 8188
rect 31796 8186 31802 8188
rect 31556 8134 31558 8186
rect 31738 8134 31740 8186
rect 31494 8132 31500 8134
rect 31556 8132 31580 8134
rect 31636 8132 31660 8134
rect 31716 8132 31740 8134
rect 31796 8132 31802 8134
rect 31494 8123 31802 8132
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 28276 7478 28304 8026
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28354 7848 28410 7857
rect 28354 7783 28356 7792
rect 28408 7783 28410 7792
rect 28356 7754 28408 7760
rect 28264 7472 28316 7478
rect 28264 7414 28316 7420
rect 28276 6866 28304 7414
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28368 6474 28396 7754
rect 28540 7744 28592 7750
rect 28540 7686 28592 7692
rect 28552 6934 28580 7686
rect 28540 6928 28592 6934
rect 28540 6870 28592 6876
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28368 6458 28488 6474
rect 28644 6458 28672 6598
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28356 6452 28488 6458
rect 28408 6446 28488 6452
rect 28356 6394 28408 6400
rect 28080 6248 28132 6254
rect 27618 6216 27674 6225
rect 28080 6190 28132 6196
rect 27618 6151 27620 6160
rect 27672 6151 27674 6160
rect 27988 6180 28040 6186
rect 27620 6122 27672 6128
rect 27988 6122 28040 6128
rect 27607 5468 27915 5477
rect 27607 5466 27613 5468
rect 27669 5466 27693 5468
rect 27749 5466 27773 5468
rect 27829 5466 27853 5468
rect 27909 5466 27915 5468
rect 27669 5414 27671 5466
rect 27851 5414 27853 5466
rect 27607 5412 27613 5414
rect 27669 5412 27693 5414
rect 27749 5412 27773 5414
rect 27829 5412 27853 5414
rect 27909 5412 27915 5414
rect 27607 5403 27915 5412
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27632 4593 27660 4966
rect 27618 4584 27674 4593
rect 27528 4548 27580 4554
rect 27618 4519 27674 4528
rect 27528 4490 27580 4496
rect 27540 4010 27568 4490
rect 27607 4380 27915 4389
rect 27607 4378 27613 4380
rect 27669 4378 27693 4380
rect 27749 4378 27773 4380
rect 27829 4378 27853 4380
rect 27909 4378 27915 4380
rect 27669 4326 27671 4378
rect 27851 4326 27853 4378
rect 27607 4324 27613 4326
rect 27669 4324 27693 4326
rect 27749 4324 27773 4326
rect 27829 4324 27853 4326
rect 27909 4324 27915 4326
rect 27607 4315 27915 4324
rect 28000 4078 28028 6122
rect 28092 5846 28120 6190
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 28080 5840 28132 5846
rect 28080 5782 28132 5788
rect 28092 5234 28120 5782
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28368 5166 28396 6122
rect 28460 5778 28488 6446
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 28736 6254 28764 7890
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28816 7268 28868 7274
rect 28816 7210 28868 7216
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 28828 5914 28856 7210
rect 29012 7002 29040 7482
rect 31494 7100 31802 7109
rect 31494 7098 31500 7100
rect 31556 7098 31580 7100
rect 31636 7098 31660 7100
rect 31716 7098 31740 7100
rect 31796 7098 31802 7100
rect 31556 7046 31558 7098
rect 31738 7046 31740 7098
rect 31494 7044 31500 7046
rect 31556 7044 31580 7046
rect 31636 7044 31660 7046
rect 31716 7044 31740 7046
rect 31796 7044 31802 7046
rect 31494 7035 31802 7044
rect 29000 6996 29052 7002
rect 29000 6938 29052 6944
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28460 5574 28488 5714
rect 29012 5710 29040 6054
rect 29380 5914 29408 6190
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 29656 5778 29684 6054
rect 31494 6012 31802 6021
rect 31494 6010 31500 6012
rect 31556 6010 31580 6012
rect 31636 6010 31660 6012
rect 31716 6010 31740 6012
rect 31796 6010 31802 6012
rect 31556 5958 31558 6010
rect 31738 5958 31740 6010
rect 31494 5956 31500 5958
rect 31556 5956 31580 5958
rect 31636 5956 31660 5958
rect 31716 5956 31740 5958
rect 31796 5956 31802 5958
rect 31494 5947 31802 5956
rect 29644 5772 29696 5778
rect 29644 5714 29696 5720
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28632 5568 28684 5574
rect 28632 5510 28684 5516
rect 28644 5370 28672 5510
rect 28632 5364 28684 5370
rect 28632 5306 28684 5312
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28080 5092 28132 5098
rect 28080 5034 28132 5040
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27436 3596 27488 3602
rect 27436 3538 27488 3544
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27172 3194 27200 3470
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 26976 3120 27028 3126
rect 26976 3062 27028 3068
rect 27448 3058 27476 3538
rect 27607 3292 27915 3301
rect 27607 3290 27613 3292
rect 27669 3290 27693 3292
rect 27749 3290 27773 3292
rect 27829 3290 27853 3292
rect 27909 3290 27915 3292
rect 27669 3238 27671 3290
rect 27851 3238 27853 3290
rect 27607 3236 27613 3238
rect 27669 3236 27693 3238
rect 27749 3236 27773 3238
rect 27829 3236 27853 3238
rect 27909 3236 27915 3238
rect 27607 3227 27915 3236
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25280 2468 25360 2496
rect 25228 2450 25280 2456
rect 25332 2106 25360 2468
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25516 2106 25544 2450
rect 25608 2446 25636 2926
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 26436 2514 26464 2790
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25320 2100 25372 2106
rect 25320 2042 25372 2048
rect 25504 2100 25556 2106
rect 25504 2042 25556 2048
rect 25700 2038 25728 2450
rect 25976 2106 26004 2450
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 25964 2100 26016 2106
rect 25964 2042 26016 2048
rect 26160 2038 26188 2382
rect 26516 2372 26568 2378
rect 26516 2314 26568 2320
rect 25688 2032 25740 2038
rect 25688 1974 25740 1980
rect 26148 2032 26200 2038
rect 26148 1974 26200 1980
rect 24860 1964 24912 1970
rect 24860 1906 24912 1912
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 24768 1886 24820 1892
rect 24768 1828 24820 1834
rect 24860 1828 24912 1834
rect 24860 1770 24912 1776
rect 24872 1714 24900 1770
rect 24688 1686 24900 1714
rect 23720 1660 24028 1669
rect 23720 1658 23726 1660
rect 23782 1658 23806 1660
rect 23862 1658 23886 1660
rect 23942 1658 23966 1660
rect 24022 1658 24028 1660
rect 23782 1606 23784 1658
rect 23964 1606 23966 1658
rect 23720 1604 23726 1606
rect 23782 1604 23806 1606
rect 23862 1604 23886 1606
rect 23942 1604 23966 1606
rect 24022 1604 24028 1606
rect 23720 1595 24028 1604
rect 26252 1562 26280 1906
rect 26528 1834 26556 2314
rect 26620 2106 26648 2586
rect 27356 2378 27384 2790
rect 27344 2372 27396 2378
rect 27344 2314 27396 2320
rect 27607 2204 27915 2213
rect 27607 2202 27613 2204
rect 27669 2202 27693 2204
rect 27749 2202 27773 2204
rect 27829 2202 27853 2204
rect 27909 2202 27915 2204
rect 27669 2150 27671 2202
rect 27851 2150 27853 2202
rect 27607 2148 27613 2150
rect 27669 2148 27693 2150
rect 27749 2148 27773 2150
rect 27829 2148 27853 2150
rect 27909 2148 27915 2150
rect 27607 2139 27915 2148
rect 26608 2100 26660 2106
rect 26608 2042 26660 2048
rect 28000 1970 28028 4014
rect 28092 4010 28120 5034
rect 28264 5024 28316 5030
rect 28264 4966 28316 4972
rect 28080 4004 28132 4010
rect 28080 3946 28132 3952
rect 28172 4004 28224 4010
rect 28172 3946 28224 3952
rect 28184 3738 28212 3946
rect 28276 3777 28304 4966
rect 28262 3768 28318 3777
rect 28172 3732 28224 3738
rect 28262 3703 28318 3712
rect 28172 3674 28224 3680
rect 28644 3097 28672 5306
rect 29104 5166 29132 5578
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 5166 29592 5510
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 29644 5024 29696 5030
rect 29644 4966 29696 4972
rect 29656 4486 29684 4966
rect 31494 4924 31802 4933
rect 31494 4922 31500 4924
rect 31556 4922 31580 4924
rect 31636 4922 31660 4924
rect 31716 4922 31740 4924
rect 31796 4922 31802 4924
rect 31556 4870 31558 4922
rect 31738 4870 31740 4922
rect 31494 4868 31500 4870
rect 31556 4868 31580 4870
rect 31636 4868 31660 4870
rect 31716 4868 31740 4870
rect 31796 4868 31802 4870
rect 31494 4859 31802 4868
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 31494 3836 31802 3845
rect 31494 3834 31500 3836
rect 31556 3834 31580 3836
rect 31636 3834 31660 3836
rect 31716 3834 31740 3836
rect 31796 3834 31802 3836
rect 31556 3782 31558 3834
rect 31738 3782 31740 3834
rect 31494 3780 31500 3782
rect 31556 3780 31580 3782
rect 31636 3780 31660 3782
rect 31716 3780 31740 3782
rect 31796 3780 31802 3782
rect 31494 3771 31802 3780
rect 28630 3088 28686 3097
rect 28630 3023 28686 3032
rect 31494 2748 31802 2757
rect 31494 2746 31500 2748
rect 31556 2746 31580 2748
rect 31636 2746 31660 2748
rect 31716 2746 31740 2748
rect 31796 2746 31802 2748
rect 31556 2694 31558 2746
rect 31738 2694 31740 2746
rect 31494 2692 31500 2694
rect 31556 2692 31580 2694
rect 31636 2692 31660 2694
rect 31716 2692 31740 2694
rect 31796 2692 31802 2694
rect 31494 2683 31802 2692
rect 27988 1964 28040 1970
rect 27988 1906 28040 1912
rect 26516 1828 26568 1834
rect 26516 1770 26568 1776
rect 31494 1660 31802 1669
rect 31494 1658 31500 1660
rect 31556 1658 31580 1660
rect 31636 1658 31660 1660
rect 31716 1658 31740 1660
rect 31796 1658 31802 1660
rect 31556 1606 31558 1658
rect 31738 1606 31740 1658
rect 31494 1604 31500 1606
rect 31556 1604 31580 1606
rect 31636 1604 31660 1606
rect 31716 1604 31740 1606
rect 31796 1604 31802 1606
rect 31494 1595 31802 1604
rect 26240 1556 26292 1562
rect 26240 1498 26292 1504
rect 21824 1488 21876 1494
rect 21824 1430 21876 1436
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 19708 1420 19760 1426
rect 19708 1362 19760 1368
rect 19064 1352 19116 1358
rect 19064 1294 19116 1300
rect 4285 1116 4593 1125
rect 4285 1114 4291 1116
rect 4347 1114 4371 1116
rect 4427 1114 4451 1116
rect 4507 1114 4531 1116
rect 4587 1114 4593 1116
rect 4347 1062 4349 1114
rect 4529 1062 4531 1114
rect 4285 1060 4291 1062
rect 4347 1060 4371 1062
rect 4427 1060 4451 1062
rect 4507 1060 4531 1062
rect 4587 1060 4593 1062
rect 4285 1051 4593 1060
rect 12059 1116 12367 1125
rect 12059 1114 12065 1116
rect 12121 1114 12145 1116
rect 12201 1114 12225 1116
rect 12281 1114 12305 1116
rect 12361 1114 12367 1116
rect 12121 1062 12123 1114
rect 12303 1062 12305 1114
rect 12059 1060 12065 1062
rect 12121 1060 12145 1062
rect 12201 1060 12225 1062
rect 12281 1060 12305 1062
rect 12361 1060 12367 1062
rect 12059 1051 12367 1060
rect 19833 1116 20141 1125
rect 19833 1114 19839 1116
rect 19895 1114 19919 1116
rect 19975 1114 19999 1116
rect 20055 1114 20079 1116
rect 20135 1114 20141 1116
rect 19895 1062 19897 1114
rect 20077 1062 20079 1114
rect 19833 1060 19839 1062
rect 19895 1060 19919 1062
rect 19975 1060 19999 1062
rect 20055 1060 20079 1062
rect 20135 1060 20141 1062
rect 19833 1051 20141 1060
rect 27607 1116 27915 1125
rect 27607 1114 27613 1116
rect 27669 1114 27693 1116
rect 27749 1114 27773 1116
rect 27829 1114 27853 1116
rect 27909 1114 27915 1116
rect 27669 1062 27671 1114
rect 27851 1062 27853 1114
rect 27607 1060 27613 1062
rect 27669 1060 27693 1062
rect 27749 1060 27773 1062
rect 27829 1060 27853 1062
rect 27909 1060 27915 1062
rect 27607 1051 27915 1060
rect 8172 572 8480 581
rect 8172 570 8178 572
rect 8234 570 8258 572
rect 8314 570 8338 572
rect 8394 570 8418 572
rect 8474 570 8480 572
rect 8234 518 8236 570
rect 8416 518 8418 570
rect 8172 516 8178 518
rect 8234 516 8258 518
rect 8314 516 8338 518
rect 8394 516 8418 518
rect 8474 516 8480 518
rect 8172 507 8480 516
rect 15946 572 16254 581
rect 15946 570 15952 572
rect 16008 570 16032 572
rect 16088 570 16112 572
rect 16168 570 16192 572
rect 16248 570 16254 572
rect 16008 518 16010 570
rect 16190 518 16192 570
rect 15946 516 15952 518
rect 16008 516 16032 518
rect 16088 516 16112 518
rect 16168 516 16192 518
rect 16248 516 16254 518
rect 15946 507 16254 516
rect 23720 572 24028 581
rect 23720 570 23726 572
rect 23782 570 23806 572
rect 23862 570 23886 572
rect 23942 570 23966 572
rect 24022 570 24028 572
rect 23782 518 23784 570
rect 23964 518 23966 570
rect 23720 516 23726 518
rect 23782 516 23806 518
rect 23862 516 23886 518
rect 23942 516 23966 518
rect 24022 516 24028 518
rect 23720 507 24028 516
rect 31494 572 31802 581
rect 31494 570 31500 572
rect 31556 570 31580 572
rect 31636 570 31660 572
rect 31716 570 31740 572
rect 31796 570 31802 572
rect 31556 518 31558 570
rect 31738 518 31740 570
rect 31494 516 31500 518
rect 31556 516 31580 518
rect 31636 516 31660 518
rect 31716 516 31740 518
rect 31796 516 31802 518
rect 31494 507 31802 516
<< via2 >>
rect 4526 21936 4582 21992
rect 1306 21256 1362 21312
rect 2134 21140 2190 21176
rect 2134 21120 2136 21140
rect 2136 21120 2188 21140
rect 2188 21120 2190 21140
rect 1582 20712 1638 20768
rect 2502 18808 2558 18864
rect 3330 20712 3386 20768
rect 3974 21140 4030 21176
rect 4291 21786 4347 21788
rect 4371 21786 4427 21788
rect 4451 21786 4507 21788
rect 4531 21786 4587 21788
rect 4291 21734 4337 21786
rect 4337 21734 4347 21786
rect 4371 21734 4401 21786
rect 4401 21734 4413 21786
rect 4413 21734 4427 21786
rect 4451 21734 4465 21786
rect 4465 21734 4477 21786
rect 4477 21734 4507 21786
rect 4531 21734 4541 21786
rect 4541 21734 4587 21786
rect 4291 21732 4347 21734
rect 4371 21732 4427 21734
rect 4451 21732 4507 21734
rect 4531 21732 4587 21734
rect 3974 21120 3976 21140
rect 3976 21120 4028 21140
rect 4028 21120 4030 21140
rect 4291 20698 4347 20700
rect 4371 20698 4427 20700
rect 4451 20698 4507 20700
rect 4531 20698 4587 20700
rect 4291 20646 4337 20698
rect 4337 20646 4347 20698
rect 4371 20646 4401 20698
rect 4401 20646 4413 20698
rect 4413 20646 4427 20698
rect 4451 20646 4465 20698
rect 4465 20646 4477 20698
rect 4477 20646 4507 20698
rect 4531 20646 4541 20698
rect 4541 20646 4587 20698
rect 4291 20644 4347 20646
rect 4371 20644 4427 20646
rect 4451 20644 4507 20646
rect 4531 20644 4587 20646
rect 4986 21564 4988 21584
rect 4988 21564 5040 21584
rect 5040 21564 5042 21584
rect 4986 21528 5042 21564
rect 12530 21936 12586 21992
rect 7010 21800 7066 21856
rect 8850 21800 8906 21856
rect 2686 17992 2742 18048
rect 1030 7384 1086 7440
rect 1766 6840 1822 6896
rect 3790 18148 3846 18184
rect 3790 18128 3792 18148
rect 3792 18128 3844 18148
rect 3844 18128 3846 18148
rect 4291 19610 4347 19612
rect 4371 19610 4427 19612
rect 4451 19610 4507 19612
rect 4531 19610 4587 19612
rect 4291 19558 4337 19610
rect 4337 19558 4347 19610
rect 4371 19558 4401 19610
rect 4401 19558 4413 19610
rect 4413 19558 4427 19610
rect 4451 19558 4465 19610
rect 4465 19558 4477 19610
rect 4477 19558 4507 19610
rect 4531 19558 4541 19610
rect 4541 19558 4587 19610
rect 4291 19556 4347 19558
rect 4371 19556 4427 19558
rect 4451 19556 4507 19558
rect 4531 19556 4587 19558
rect 4250 19352 4306 19408
rect 4342 18808 4398 18864
rect 4250 18692 4306 18728
rect 4250 18672 4252 18692
rect 4252 18672 4304 18692
rect 4304 18672 4306 18692
rect 4291 18522 4347 18524
rect 4371 18522 4427 18524
rect 4451 18522 4507 18524
rect 4531 18522 4587 18524
rect 4291 18470 4337 18522
rect 4337 18470 4347 18522
rect 4371 18470 4401 18522
rect 4401 18470 4413 18522
rect 4413 18470 4427 18522
rect 4451 18470 4465 18522
rect 4465 18470 4477 18522
rect 4477 18470 4507 18522
rect 4531 18470 4541 18522
rect 4541 18470 4587 18522
rect 4291 18468 4347 18470
rect 4371 18468 4427 18470
rect 4451 18468 4507 18470
rect 4531 18468 4587 18470
rect 3974 17992 4030 18048
rect 2042 8064 2098 8120
rect 1950 6704 2006 6760
rect 4434 18148 4490 18184
rect 6182 21292 6184 21312
rect 6184 21292 6236 21312
rect 6236 21292 6238 21312
rect 6182 21256 6238 21292
rect 4434 18128 4436 18148
rect 4436 18128 4488 18148
rect 4488 18128 4490 18148
rect 4291 17434 4347 17436
rect 4371 17434 4427 17436
rect 4451 17434 4507 17436
rect 4531 17434 4587 17436
rect 4291 17382 4337 17434
rect 4337 17382 4347 17434
rect 4371 17382 4401 17434
rect 4401 17382 4413 17434
rect 4413 17382 4427 17434
rect 4451 17382 4465 17434
rect 4465 17382 4477 17434
rect 4477 17382 4507 17434
rect 4531 17382 4541 17434
rect 4541 17382 4587 17434
rect 4291 17380 4347 17382
rect 4371 17380 4427 17382
rect 4451 17380 4507 17382
rect 4531 17380 4587 17382
rect 4291 16346 4347 16348
rect 4371 16346 4427 16348
rect 4451 16346 4507 16348
rect 4531 16346 4587 16348
rect 4291 16294 4337 16346
rect 4337 16294 4347 16346
rect 4371 16294 4401 16346
rect 4401 16294 4413 16346
rect 4413 16294 4427 16346
rect 4451 16294 4465 16346
rect 4465 16294 4477 16346
rect 4477 16294 4507 16346
rect 4531 16294 4541 16346
rect 4541 16294 4587 16346
rect 4291 16292 4347 16294
rect 4371 16292 4427 16294
rect 4451 16292 4507 16294
rect 4531 16292 4587 16294
rect 4291 15258 4347 15260
rect 4371 15258 4427 15260
rect 4451 15258 4507 15260
rect 4531 15258 4587 15260
rect 4291 15206 4337 15258
rect 4337 15206 4347 15258
rect 4371 15206 4401 15258
rect 4401 15206 4413 15258
rect 4413 15206 4427 15258
rect 4451 15206 4465 15258
rect 4465 15206 4477 15258
rect 4477 15206 4507 15258
rect 4531 15206 4541 15258
rect 4541 15206 4587 15258
rect 4291 15204 4347 15206
rect 4371 15204 4427 15206
rect 4451 15204 4507 15206
rect 4531 15204 4587 15206
rect 4291 14170 4347 14172
rect 4371 14170 4427 14172
rect 4451 14170 4507 14172
rect 4531 14170 4587 14172
rect 4291 14118 4337 14170
rect 4337 14118 4347 14170
rect 4371 14118 4401 14170
rect 4401 14118 4413 14170
rect 4413 14118 4427 14170
rect 4451 14118 4465 14170
rect 4465 14118 4477 14170
rect 4477 14118 4507 14170
rect 4531 14118 4541 14170
rect 4541 14118 4587 14170
rect 4291 14116 4347 14118
rect 4371 14116 4427 14118
rect 4451 14116 4507 14118
rect 4531 14116 4587 14118
rect 4291 13082 4347 13084
rect 4371 13082 4427 13084
rect 4451 13082 4507 13084
rect 4531 13082 4587 13084
rect 4291 13030 4337 13082
rect 4337 13030 4347 13082
rect 4371 13030 4401 13082
rect 4401 13030 4413 13082
rect 4413 13030 4427 13082
rect 4451 13030 4465 13082
rect 4465 13030 4477 13082
rect 4477 13030 4507 13082
rect 4531 13030 4541 13082
rect 4541 13030 4587 13082
rect 4291 13028 4347 13030
rect 4371 13028 4427 13030
rect 4451 13028 4507 13030
rect 4531 13028 4587 13030
rect 5446 18264 5502 18320
rect 5078 17176 5134 17232
rect 3238 8880 3294 8936
rect 2870 8064 2926 8120
rect 4066 10648 4122 10704
rect 4291 11994 4347 11996
rect 4371 11994 4427 11996
rect 4451 11994 4507 11996
rect 4531 11994 4587 11996
rect 4291 11942 4337 11994
rect 4337 11942 4347 11994
rect 4371 11942 4401 11994
rect 4401 11942 4413 11994
rect 4413 11942 4427 11994
rect 4451 11942 4465 11994
rect 4465 11942 4477 11994
rect 4477 11942 4507 11994
rect 4531 11942 4541 11994
rect 4541 11942 4587 11994
rect 4291 11940 4347 11942
rect 4371 11940 4427 11942
rect 4451 11940 4507 11942
rect 4531 11940 4587 11942
rect 4291 10906 4347 10908
rect 4371 10906 4427 10908
rect 4451 10906 4507 10908
rect 4531 10906 4587 10908
rect 4291 10854 4337 10906
rect 4337 10854 4347 10906
rect 4371 10854 4401 10906
rect 4401 10854 4413 10906
rect 4413 10854 4427 10906
rect 4451 10854 4465 10906
rect 4465 10854 4477 10906
rect 4477 10854 4507 10906
rect 4531 10854 4541 10906
rect 4541 10854 4587 10906
rect 4291 10852 4347 10854
rect 4371 10852 4427 10854
rect 4451 10852 4507 10854
rect 4531 10852 4587 10854
rect 4291 9818 4347 9820
rect 4371 9818 4427 9820
rect 4451 9818 4507 9820
rect 4531 9818 4587 9820
rect 4291 9766 4337 9818
rect 4337 9766 4347 9818
rect 4371 9766 4401 9818
rect 4401 9766 4413 9818
rect 4413 9766 4427 9818
rect 4451 9766 4465 9818
rect 4465 9766 4477 9818
rect 4477 9766 4507 9818
rect 4531 9766 4541 9818
rect 4541 9766 4587 9818
rect 4291 9764 4347 9766
rect 4371 9764 4427 9766
rect 4451 9764 4507 9766
rect 4531 9764 4587 9766
rect 4710 9152 4766 9208
rect 5170 12824 5226 12880
rect 5446 17620 5448 17640
rect 5448 17620 5500 17640
rect 5500 17620 5502 17640
rect 5446 17584 5502 17620
rect 5354 16088 5410 16144
rect 5906 18672 5962 18728
rect 6458 21140 6514 21176
rect 6458 21120 6460 21140
rect 6460 21120 6512 21140
rect 6512 21120 6514 21140
rect 6366 20712 6422 20768
rect 6550 19488 6606 19544
rect 6642 19236 6698 19272
rect 6642 19216 6644 19236
rect 6644 19216 6696 19236
rect 6696 19216 6698 19236
rect 5354 12280 5410 12336
rect 4291 8730 4347 8732
rect 4371 8730 4427 8732
rect 4451 8730 4507 8732
rect 4531 8730 4587 8732
rect 4291 8678 4337 8730
rect 4337 8678 4347 8730
rect 4371 8678 4401 8730
rect 4401 8678 4413 8730
rect 4413 8678 4427 8730
rect 4451 8678 4465 8730
rect 4465 8678 4477 8730
rect 4477 8678 4507 8730
rect 4531 8678 4541 8730
rect 4541 8678 4587 8730
rect 4291 8676 4347 8678
rect 4371 8676 4427 8678
rect 4451 8676 4507 8678
rect 4531 8676 4587 8678
rect 4066 8064 4122 8120
rect 3882 6976 3938 7032
rect 4291 7642 4347 7644
rect 4371 7642 4427 7644
rect 4451 7642 4507 7644
rect 4531 7642 4587 7644
rect 4291 7590 4337 7642
rect 4337 7590 4347 7642
rect 4371 7590 4401 7642
rect 4401 7590 4413 7642
rect 4413 7590 4427 7642
rect 4451 7590 4465 7642
rect 4465 7590 4477 7642
rect 4477 7590 4507 7642
rect 4531 7590 4541 7642
rect 4541 7590 4587 7642
rect 4291 7588 4347 7590
rect 4371 7588 4427 7590
rect 4451 7588 4507 7590
rect 4531 7588 4587 7590
rect 3974 6180 4030 6216
rect 3974 6160 3976 6180
rect 3976 6160 4028 6180
rect 4028 6160 4030 6180
rect 4526 6740 4528 6760
rect 4528 6740 4580 6760
rect 4580 6740 4582 6760
rect 4526 6704 4582 6740
rect 4291 6554 4347 6556
rect 4371 6554 4427 6556
rect 4451 6554 4507 6556
rect 4531 6554 4587 6556
rect 4291 6502 4337 6554
rect 4337 6502 4347 6554
rect 4371 6502 4401 6554
rect 4401 6502 4413 6554
rect 4413 6502 4427 6554
rect 4451 6502 4465 6554
rect 4465 6502 4477 6554
rect 4477 6502 4507 6554
rect 4531 6502 4541 6554
rect 4541 6502 4587 6554
rect 4291 6500 4347 6502
rect 4371 6500 4427 6502
rect 4451 6500 4507 6502
rect 4531 6500 4587 6502
rect 4291 5466 4347 5468
rect 4371 5466 4427 5468
rect 4451 5466 4507 5468
rect 4531 5466 4587 5468
rect 4291 5414 4337 5466
rect 4337 5414 4347 5466
rect 4371 5414 4401 5466
rect 4401 5414 4413 5466
rect 4413 5414 4427 5466
rect 4451 5414 4465 5466
rect 4465 5414 4477 5466
rect 4477 5414 4507 5466
rect 4531 5414 4541 5466
rect 4541 5414 4587 5466
rect 4291 5412 4347 5414
rect 4371 5412 4427 5414
rect 4451 5412 4507 5414
rect 4531 5412 4587 5414
rect 5262 11056 5318 11112
rect 5170 9560 5226 9616
rect 5170 8880 5226 8936
rect 4986 6568 5042 6624
rect 6458 18128 6514 18184
rect 5722 9016 5778 9072
rect 5630 8336 5686 8392
rect 5446 7792 5502 7848
rect 5446 7692 5448 7712
rect 5448 7692 5500 7712
rect 5500 7692 5502 7712
rect 5446 7656 5502 7692
rect 5446 7112 5502 7168
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 7930 20576 7986 20632
rect 8666 20596 8722 20632
rect 8666 20576 8668 20596
rect 8668 20576 8720 20596
rect 8720 20576 8722 20596
rect 7838 20460 7894 20496
rect 7838 20440 7840 20460
rect 7840 20440 7892 20460
rect 7892 20440 7894 20460
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 6642 16632 6698 16688
rect 6182 9560 6238 9616
rect 5906 7928 5962 7984
rect 5446 6840 5502 6896
rect 5446 6724 5502 6760
rect 5446 6704 5448 6724
rect 5448 6704 5500 6724
rect 5500 6704 5502 6724
rect 5814 6432 5870 6488
rect 4291 4378 4347 4380
rect 4371 4378 4427 4380
rect 4451 4378 4507 4380
rect 4531 4378 4587 4380
rect 4291 4326 4337 4378
rect 4337 4326 4347 4378
rect 4371 4326 4401 4378
rect 4401 4326 4413 4378
rect 4413 4326 4427 4378
rect 4451 4326 4465 4378
rect 4465 4326 4477 4378
rect 4477 4326 4507 4378
rect 4531 4326 4541 4378
rect 4541 4326 4587 4378
rect 4291 4324 4347 4326
rect 4371 4324 4427 4326
rect 4451 4324 4507 4326
rect 4531 4324 4587 4326
rect 6090 9424 6146 9480
rect 6090 8744 6146 8800
rect 6550 10512 6606 10568
rect 7102 11600 7158 11656
rect 7654 18264 7710 18320
rect 7838 17484 7840 17504
rect 7840 17484 7892 17504
rect 7892 17484 7894 17504
rect 7838 17448 7894 17484
rect 6918 9968 6974 10024
rect 6458 8064 6514 8120
rect 6734 8472 6790 8528
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 8574 17992 8630 18048
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 8114 17720 8170 17776
rect 7654 13776 7710 13832
rect 8482 17040 8538 17096
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 8482 16360 8538 16416
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 8390 15136 8446 15192
rect 8574 15136 8630 15192
rect 7930 12688 7986 12744
rect 7746 10684 7748 10704
rect 7748 10684 7800 10704
rect 7800 10684 7802 10704
rect 7746 10648 7802 10684
rect 7378 9560 7434 9616
rect 7194 9152 7250 9208
rect 7102 8900 7158 8936
rect 7102 8880 7104 8900
rect 7104 8880 7156 8900
rect 7156 8880 7158 8900
rect 6090 5752 6146 5808
rect 4291 3290 4347 3292
rect 4371 3290 4427 3292
rect 4451 3290 4507 3292
rect 4531 3290 4587 3292
rect 4291 3238 4337 3290
rect 4337 3238 4347 3290
rect 4371 3238 4401 3290
rect 4401 3238 4413 3290
rect 4413 3238 4427 3290
rect 4451 3238 4465 3290
rect 4465 3238 4477 3290
rect 4477 3238 4507 3290
rect 4531 3238 4541 3290
rect 4541 3238 4587 3290
rect 4291 3236 4347 3238
rect 4371 3236 4427 3238
rect 4451 3236 4507 3238
rect 4531 3236 4587 3238
rect 6734 7248 6790 7304
rect 6642 6568 6698 6624
rect 7010 7948 7066 7984
rect 7010 7928 7012 7948
rect 7012 7928 7064 7948
rect 7064 7928 7066 7948
rect 7286 8336 7342 8392
rect 6918 5908 6974 5944
rect 6918 5888 6920 5908
rect 6920 5888 6972 5908
rect 6972 5888 6974 5908
rect 7286 7112 7342 7168
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 12065 21786 12121 21788
rect 12145 21786 12201 21788
rect 12225 21786 12281 21788
rect 12305 21786 12361 21788
rect 12065 21734 12111 21786
rect 12111 21734 12121 21786
rect 12145 21734 12175 21786
rect 12175 21734 12187 21786
rect 12187 21734 12201 21786
rect 12225 21734 12239 21786
rect 12239 21734 12251 21786
rect 12251 21734 12281 21786
rect 12305 21734 12315 21786
rect 12315 21734 12361 21786
rect 12065 21732 12121 21734
rect 12145 21732 12201 21734
rect 12225 21732 12281 21734
rect 12305 21732 12361 21734
rect 13358 21664 13414 21720
rect 10414 20984 10470 21040
rect 10322 20712 10378 20768
rect 10782 19896 10838 19952
rect 10138 19624 10194 19680
rect 9494 19352 9550 19408
rect 10046 19352 10102 19408
rect 9126 18672 9182 18728
rect 9034 18264 9090 18320
rect 8574 13912 8630 13968
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8390 13232 8446 13288
rect 8114 13096 8170 13152
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8942 14900 8944 14920
rect 8944 14900 8996 14920
rect 8996 14900 8998 14920
rect 8942 14864 8998 14900
rect 9218 17312 9274 17368
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8206 10140 8208 10160
rect 8208 10140 8260 10160
rect 8260 10140 8262 10160
rect 8206 10104 8262 10140
rect 8298 9968 8354 10024
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8022 9152 8078 9208
rect 8666 10648 8722 10704
rect 8114 8900 8170 8936
rect 8114 8880 8116 8900
rect 8116 8880 8168 8900
rect 8168 8880 8170 8900
rect 8482 8880 8538 8936
rect 7930 8744 7986 8800
rect 7930 8608 7986 8664
rect 8390 8492 8446 8528
rect 8390 8472 8392 8492
rect 8392 8472 8444 8492
rect 8444 8472 8446 8492
rect 8390 8356 8446 8392
rect 8390 8336 8392 8356
rect 8392 8336 8444 8356
rect 8444 8336 8446 8356
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 9310 16904 9366 16960
rect 9402 16768 9458 16824
rect 9954 18264 10010 18320
rect 10690 19216 10746 19272
rect 11150 19488 11206 19544
rect 11150 18944 11206 19000
rect 10138 17856 10194 17912
rect 10138 17740 10194 17776
rect 10138 17720 10140 17740
rect 10140 17720 10192 17740
rect 10192 17720 10194 17740
rect 11058 18692 11114 18728
rect 11058 18672 11060 18692
rect 11060 18672 11112 18692
rect 11112 18672 11114 18692
rect 10506 17312 10562 17368
rect 10874 17992 10930 18048
rect 9310 15136 9366 15192
rect 9678 15544 9734 15600
rect 9954 15408 10010 15464
rect 9770 14728 9826 14784
rect 9954 14320 10010 14376
rect 9126 12144 9182 12200
rect 9034 11600 9090 11656
rect 9954 13812 9956 13832
rect 9956 13812 10008 13832
rect 10008 13812 10010 13832
rect 9954 13776 10010 13812
rect 9954 13640 10010 13696
rect 8942 10920 8998 10976
rect 10966 17448 11022 17504
rect 10874 17176 10930 17232
rect 11150 17856 11206 17912
rect 10598 16652 10654 16688
rect 10598 16632 10600 16652
rect 10600 16632 10652 16652
rect 10652 16632 10654 16652
rect 10690 16360 10746 16416
rect 10966 16904 11022 16960
rect 10414 16088 10470 16144
rect 10138 13912 10194 13968
rect 10782 14864 10838 14920
rect 11242 17720 11298 17776
rect 11426 20884 11428 20904
rect 11428 20884 11480 20904
rect 11480 20884 11482 20904
rect 11426 20848 11482 20884
rect 11426 19252 11428 19272
rect 11428 19252 11480 19272
rect 11480 19252 11482 19272
rect 11426 19216 11482 19252
rect 11610 19080 11666 19136
rect 11518 18808 11574 18864
rect 11058 15136 11114 15192
rect 10966 15000 11022 15056
rect 10506 13776 10562 13832
rect 9954 12688 10010 12744
rect 10138 13268 10140 13288
rect 10140 13268 10192 13288
rect 10192 13268 10194 13288
rect 10138 13232 10194 13268
rect 10506 13132 10508 13152
rect 10508 13132 10560 13152
rect 10560 13132 10562 13152
rect 8850 9444 8906 9480
rect 8850 9424 8852 9444
rect 8852 9424 8904 9444
rect 8904 9424 8906 9444
rect 8850 8472 8906 8528
rect 8022 7792 8078 7848
rect 8206 7792 8262 7848
rect 7838 6296 7894 6352
rect 7746 6024 7802 6080
rect 8574 7928 8630 7984
rect 9034 8064 9090 8120
rect 8942 7928 8998 7984
rect 8666 7812 8722 7848
rect 8666 7792 8668 7812
rect 8668 7792 8720 7812
rect 8720 7792 8722 7812
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 8206 6704 8262 6760
rect 8482 6704 8538 6760
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 8758 6976 8814 7032
rect 9678 11076 9734 11112
rect 9678 11056 9680 11076
rect 9680 11056 9732 11076
rect 9732 11056 9734 11076
rect 9494 8780 9496 8800
rect 9496 8780 9548 8800
rect 9548 8780 9550 8800
rect 9494 8744 9550 8780
rect 10506 13096 10562 13132
rect 10782 13812 10784 13832
rect 10784 13812 10836 13832
rect 10836 13812 10838 13832
rect 10782 13776 10838 13812
rect 11242 13912 11298 13968
rect 11610 16088 11666 16144
rect 12346 21004 12402 21040
rect 12346 20984 12348 21004
rect 12348 20984 12400 21004
rect 12400 20984 12402 21004
rect 11794 20596 11850 20632
rect 11794 20576 11796 20596
rect 11796 20576 11848 20596
rect 11848 20576 11850 20596
rect 12065 20698 12121 20700
rect 12145 20698 12201 20700
rect 12225 20698 12281 20700
rect 12305 20698 12361 20700
rect 12065 20646 12111 20698
rect 12111 20646 12121 20698
rect 12145 20646 12175 20698
rect 12175 20646 12187 20698
rect 12187 20646 12201 20698
rect 12225 20646 12239 20698
rect 12239 20646 12251 20698
rect 12251 20646 12281 20698
rect 12305 20646 12315 20698
rect 12315 20646 12361 20698
rect 12065 20644 12121 20646
rect 12145 20644 12201 20646
rect 12225 20644 12281 20646
rect 12305 20644 12361 20646
rect 13726 22072 13782 22128
rect 13726 21936 13782 21992
rect 13542 21528 13598 21584
rect 13266 21256 13322 21312
rect 11794 17992 11850 18048
rect 12065 19610 12121 19612
rect 12145 19610 12201 19612
rect 12225 19610 12281 19612
rect 12305 19610 12361 19612
rect 12065 19558 12111 19610
rect 12111 19558 12121 19610
rect 12145 19558 12175 19610
rect 12175 19558 12187 19610
rect 12187 19558 12201 19610
rect 12225 19558 12239 19610
rect 12239 19558 12251 19610
rect 12251 19558 12281 19610
rect 12305 19558 12315 19610
rect 12315 19558 12361 19610
rect 12065 19556 12121 19558
rect 12145 19556 12201 19558
rect 12225 19556 12281 19558
rect 12305 19556 12361 19558
rect 12065 18522 12121 18524
rect 12145 18522 12201 18524
rect 12225 18522 12281 18524
rect 12305 18522 12361 18524
rect 12065 18470 12111 18522
rect 12111 18470 12121 18522
rect 12145 18470 12175 18522
rect 12175 18470 12187 18522
rect 12187 18470 12201 18522
rect 12225 18470 12239 18522
rect 12239 18470 12251 18522
rect 12251 18470 12281 18522
rect 12305 18470 12315 18522
rect 12315 18470 12361 18522
rect 12065 18468 12121 18470
rect 12145 18468 12201 18470
rect 12225 18468 12281 18470
rect 12305 18468 12361 18470
rect 11978 17856 12034 17912
rect 12065 17434 12121 17436
rect 12145 17434 12201 17436
rect 12225 17434 12281 17436
rect 12305 17434 12361 17436
rect 12065 17382 12111 17434
rect 12111 17382 12121 17434
rect 12145 17382 12175 17434
rect 12175 17382 12187 17434
rect 12187 17382 12201 17434
rect 12225 17382 12239 17434
rect 12239 17382 12251 17434
rect 12251 17382 12281 17434
rect 12305 17382 12315 17434
rect 12315 17382 12361 17434
rect 12065 17380 12121 17382
rect 12145 17380 12201 17382
rect 12225 17380 12281 17382
rect 12305 17380 12361 17382
rect 11978 17060 12034 17096
rect 11978 17040 11980 17060
rect 11980 17040 12032 17060
rect 12032 17040 12034 17060
rect 11978 16904 12034 16960
rect 11794 16632 11850 16688
rect 12070 16496 12126 16552
rect 12065 16346 12121 16348
rect 12145 16346 12201 16348
rect 12225 16346 12281 16348
rect 12305 16346 12361 16348
rect 12065 16294 12111 16346
rect 12111 16294 12121 16346
rect 12145 16294 12175 16346
rect 12175 16294 12187 16346
rect 12187 16294 12201 16346
rect 12225 16294 12239 16346
rect 12239 16294 12251 16346
rect 12251 16294 12281 16346
rect 12305 16294 12315 16346
rect 12315 16294 12361 16346
rect 12065 16292 12121 16294
rect 12145 16292 12201 16294
rect 12225 16292 12281 16294
rect 12305 16292 12361 16294
rect 11886 14864 11942 14920
rect 11518 14728 11574 14784
rect 12065 15258 12121 15260
rect 12145 15258 12201 15260
rect 12225 15258 12281 15260
rect 12305 15258 12361 15260
rect 12065 15206 12111 15258
rect 12111 15206 12121 15258
rect 12145 15206 12175 15258
rect 12175 15206 12187 15258
rect 12187 15206 12201 15258
rect 12225 15206 12239 15258
rect 12239 15206 12251 15258
rect 12251 15206 12281 15258
rect 12305 15206 12315 15258
rect 12315 15206 12361 15258
rect 12065 15204 12121 15206
rect 12145 15204 12201 15206
rect 12225 15204 12281 15206
rect 12305 15204 12361 15206
rect 11334 13640 11390 13696
rect 10874 12824 10930 12880
rect 10782 12724 10784 12744
rect 10784 12724 10836 12744
rect 10836 12724 10838 12744
rect 10782 12688 10838 12724
rect 10690 12280 10746 12336
rect 9954 12008 10010 12064
rect 10046 11736 10102 11792
rect 10138 10376 10194 10432
rect 10322 10920 10378 10976
rect 9954 8880 10010 8936
rect 9218 6024 9274 6080
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 9586 8064 9642 8120
rect 9862 8064 9918 8120
rect 9770 7928 9826 7984
rect 10138 9324 10140 9344
rect 10140 9324 10192 9344
rect 10192 9324 10194 9344
rect 10138 9288 10194 9324
rect 11150 12552 11206 12608
rect 11058 12008 11114 12064
rect 10506 10920 10562 10976
rect 10506 10376 10562 10432
rect 10414 8880 10470 8936
rect 9770 7656 9826 7712
rect 9954 7520 10010 7576
rect 10230 8064 10286 8120
rect 9770 6704 9826 6760
rect 9770 6024 9826 6080
rect 9586 5752 9642 5808
rect 10230 7284 10232 7304
rect 10232 7284 10284 7304
rect 10284 7284 10286 7304
rect 10230 7248 10286 7284
rect 10414 6840 10470 6896
rect 10322 6568 10378 6624
rect 10322 5888 10378 5944
rect 10322 5480 10378 5536
rect 10322 4936 10378 4992
rect 10414 4800 10470 4856
rect 12065 14170 12121 14172
rect 12145 14170 12201 14172
rect 12225 14170 12281 14172
rect 12305 14170 12361 14172
rect 12065 14118 12111 14170
rect 12111 14118 12121 14170
rect 12145 14118 12175 14170
rect 12175 14118 12187 14170
rect 12187 14118 12201 14170
rect 12225 14118 12239 14170
rect 12239 14118 12251 14170
rect 12251 14118 12281 14170
rect 12305 14118 12315 14170
rect 12315 14118 12361 14170
rect 12065 14116 12121 14118
rect 12145 14116 12201 14118
rect 12225 14116 12281 14118
rect 12305 14116 12361 14118
rect 11886 13776 11942 13832
rect 11794 13640 11850 13696
rect 12530 14864 12586 14920
rect 12714 14320 12770 14376
rect 11794 13232 11850 13288
rect 12065 13082 12121 13084
rect 12145 13082 12201 13084
rect 12225 13082 12281 13084
rect 12305 13082 12361 13084
rect 12065 13030 12111 13082
rect 12111 13030 12121 13082
rect 12145 13030 12175 13082
rect 12175 13030 12187 13082
rect 12187 13030 12201 13082
rect 12225 13030 12239 13082
rect 12239 13030 12251 13082
rect 12251 13030 12281 13082
rect 12305 13030 12315 13082
rect 12315 13030 12361 13082
rect 12065 13028 12121 13030
rect 12145 13028 12201 13030
rect 12225 13028 12281 13030
rect 12305 13028 12361 13030
rect 11702 11636 11704 11656
rect 11704 11636 11756 11656
rect 11756 11636 11758 11656
rect 11702 11600 11758 11636
rect 10874 10784 10930 10840
rect 10966 10412 10968 10432
rect 10968 10412 11020 10432
rect 11020 10412 11022 10432
rect 10966 10376 11022 10412
rect 11518 11212 11574 11248
rect 11518 11192 11520 11212
rect 11520 11192 11572 11212
rect 11572 11192 11574 11212
rect 11334 11092 11336 11112
rect 11336 11092 11388 11112
rect 11388 11092 11390 11112
rect 11334 11056 11390 11092
rect 11334 10648 11390 10704
rect 10874 9832 10930 9888
rect 12065 11994 12121 11996
rect 12145 11994 12201 11996
rect 12225 11994 12281 11996
rect 12305 11994 12361 11996
rect 12065 11942 12111 11994
rect 12111 11942 12121 11994
rect 12145 11942 12175 11994
rect 12175 11942 12187 11994
rect 12187 11942 12201 11994
rect 12225 11942 12239 11994
rect 12239 11942 12251 11994
rect 12251 11942 12281 11994
rect 12305 11942 12315 11994
rect 12315 11942 12361 11994
rect 12065 11940 12121 11942
rect 12145 11940 12201 11942
rect 12225 11940 12281 11942
rect 12305 11940 12361 11942
rect 12070 11736 12126 11792
rect 11794 10920 11850 10976
rect 12438 11464 12494 11520
rect 11886 9832 11942 9888
rect 12065 10906 12121 10908
rect 12145 10906 12201 10908
rect 12225 10906 12281 10908
rect 12305 10906 12361 10908
rect 12065 10854 12111 10906
rect 12111 10854 12121 10906
rect 12145 10854 12175 10906
rect 12175 10854 12187 10906
rect 12187 10854 12201 10906
rect 12225 10854 12239 10906
rect 12239 10854 12251 10906
rect 12251 10854 12281 10906
rect 12305 10854 12315 10906
rect 12315 10854 12361 10906
rect 12065 10852 12121 10854
rect 12145 10852 12201 10854
rect 12225 10852 12281 10854
rect 12305 10852 12361 10854
rect 13266 19352 13322 19408
rect 12990 18400 13046 18456
rect 13358 18264 13414 18320
rect 13358 18128 13414 18184
rect 13818 21800 13874 21856
rect 14738 21528 14794 21584
rect 14186 21292 14188 21312
rect 14188 21292 14240 21312
rect 14240 21292 14242 21312
rect 14186 21256 14242 21292
rect 13726 20576 13782 20632
rect 13910 19252 13912 19272
rect 13912 19252 13964 19272
rect 13964 19252 13966 19272
rect 13910 19216 13966 19252
rect 13726 18944 13782 19000
rect 13542 17740 13598 17776
rect 13542 17720 13544 17740
rect 13544 17720 13596 17740
rect 13596 17720 13598 17740
rect 13542 16632 13598 16688
rect 13082 12552 13138 12608
rect 12990 11736 13046 11792
rect 12714 11328 12770 11384
rect 12162 10240 12218 10296
rect 12162 9968 12218 10024
rect 12346 9988 12402 10024
rect 12346 9968 12348 9988
rect 12348 9968 12400 9988
rect 12400 9968 12402 9988
rect 12065 9818 12121 9820
rect 12145 9818 12201 9820
rect 12225 9818 12281 9820
rect 12305 9818 12361 9820
rect 12065 9766 12111 9818
rect 12111 9766 12121 9818
rect 12145 9766 12175 9818
rect 12175 9766 12187 9818
rect 12187 9766 12201 9818
rect 12225 9766 12239 9818
rect 12239 9766 12251 9818
rect 12251 9766 12281 9818
rect 12305 9766 12315 9818
rect 12315 9766 12361 9818
rect 12065 9764 12121 9766
rect 12145 9764 12201 9766
rect 12225 9764 12281 9766
rect 12305 9764 12361 9766
rect 10690 9152 10746 9208
rect 10690 8780 10692 8800
rect 10692 8780 10744 8800
rect 10744 8780 10746 8800
rect 10690 8744 10746 8780
rect 10690 8508 10692 8528
rect 10692 8508 10744 8528
rect 10744 8508 10746 8528
rect 10690 8472 10746 8508
rect 11058 9288 11114 9344
rect 11058 8744 11114 8800
rect 11058 8608 11114 8664
rect 10782 7656 10838 7712
rect 10966 7656 11022 7712
rect 10690 7384 10746 7440
rect 10690 6180 10746 6216
rect 10690 6160 10692 6180
rect 10692 6160 10744 6180
rect 10744 6160 10746 6180
rect 10598 5072 10654 5128
rect 10782 5752 10838 5808
rect 11426 8744 11482 8800
rect 11242 8336 11298 8392
rect 12254 9560 12310 9616
rect 12070 8880 12126 8936
rect 12065 8730 12121 8732
rect 12145 8730 12201 8732
rect 12225 8730 12281 8732
rect 12305 8730 12361 8732
rect 12065 8678 12111 8730
rect 12111 8678 12121 8730
rect 12145 8678 12175 8730
rect 12175 8678 12187 8730
rect 12187 8678 12201 8730
rect 12225 8678 12239 8730
rect 12239 8678 12251 8730
rect 12251 8678 12281 8730
rect 12305 8678 12315 8730
rect 12315 8678 12361 8730
rect 12065 8676 12121 8678
rect 12145 8676 12201 8678
rect 12225 8676 12281 8678
rect 12305 8676 12361 8678
rect 12806 9832 12862 9888
rect 12714 9172 12770 9208
rect 12714 9152 12716 9172
rect 12716 9152 12768 9172
rect 12768 9152 12770 9172
rect 15106 21412 15162 21448
rect 15106 21392 15108 21412
rect 15108 21392 15160 21412
rect 15160 21392 15162 21412
rect 15106 20848 15162 20904
rect 14094 17584 14150 17640
rect 13634 12144 13690 12200
rect 13726 11464 13782 11520
rect 13726 11328 13782 11384
rect 14278 18536 14334 18592
rect 14094 14220 14096 14240
rect 14096 14220 14148 14240
rect 14148 14220 14150 14240
rect 14094 14184 14150 14220
rect 14646 18400 14702 18456
rect 14646 17992 14702 18048
rect 14646 17312 14702 17368
rect 14462 16360 14518 16416
rect 14738 16088 14794 16144
rect 15106 19760 15162 19816
rect 15750 21392 15806 21448
rect 19839 21786 19895 21788
rect 19919 21786 19975 21788
rect 19999 21786 20055 21788
rect 20079 21786 20135 21788
rect 19839 21734 19885 21786
rect 19885 21734 19895 21786
rect 19919 21734 19949 21786
rect 19949 21734 19961 21786
rect 19961 21734 19975 21786
rect 19999 21734 20013 21786
rect 20013 21734 20025 21786
rect 20025 21734 20055 21786
rect 20079 21734 20089 21786
rect 20089 21734 20135 21786
rect 19839 21732 19895 21734
rect 19919 21732 19975 21734
rect 19999 21732 20055 21734
rect 20079 21732 20135 21734
rect 15952 21242 16008 21244
rect 16032 21242 16088 21244
rect 16112 21242 16168 21244
rect 16192 21242 16248 21244
rect 15952 21190 15998 21242
rect 15998 21190 16008 21242
rect 16032 21190 16062 21242
rect 16062 21190 16074 21242
rect 16074 21190 16088 21242
rect 16112 21190 16126 21242
rect 16126 21190 16138 21242
rect 16138 21190 16168 21242
rect 16192 21190 16202 21242
rect 16202 21190 16248 21242
rect 15952 21188 16008 21190
rect 16032 21188 16088 21190
rect 16112 21188 16168 21190
rect 16192 21188 16248 21190
rect 15934 20440 15990 20496
rect 15290 19080 15346 19136
rect 15198 18944 15254 19000
rect 15290 17312 15346 17368
rect 13450 10920 13506 10976
rect 13358 10648 13414 10704
rect 13174 10376 13230 10432
rect 13634 10376 13690 10432
rect 13542 10104 13598 10160
rect 14462 12280 14518 12336
rect 11518 8200 11574 8256
rect 11610 7248 11666 7304
rect 12065 7642 12121 7644
rect 12145 7642 12201 7644
rect 12225 7642 12281 7644
rect 12305 7642 12361 7644
rect 12065 7590 12111 7642
rect 12111 7590 12121 7642
rect 12145 7590 12175 7642
rect 12175 7590 12187 7642
rect 12187 7590 12201 7642
rect 12225 7590 12239 7642
rect 12239 7590 12251 7642
rect 12251 7590 12281 7642
rect 12305 7590 12315 7642
rect 12315 7590 12361 7642
rect 12065 7588 12121 7590
rect 12145 7588 12201 7590
rect 12225 7588 12281 7590
rect 12305 7588 12361 7590
rect 11794 6840 11850 6896
rect 11242 6432 11298 6488
rect 11334 5480 11390 5536
rect 11610 5752 11666 5808
rect 12065 6554 12121 6556
rect 12145 6554 12201 6556
rect 12225 6554 12281 6556
rect 12305 6554 12361 6556
rect 12065 6502 12111 6554
rect 12111 6502 12121 6554
rect 12145 6502 12175 6554
rect 12175 6502 12187 6554
rect 12187 6502 12201 6554
rect 12225 6502 12239 6554
rect 12239 6502 12251 6554
rect 12251 6502 12281 6554
rect 12305 6502 12315 6554
rect 12315 6502 12361 6554
rect 12065 6500 12121 6502
rect 12145 6500 12201 6502
rect 12225 6500 12281 6502
rect 12305 6500 12361 6502
rect 12438 6432 12494 6488
rect 12065 5466 12121 5468
rect 12145 5466 12201 5468
rect 12225 5466 12281 5468
rect 12305 5466 12361 5468
rect 12065 5414 12111 5466
rect 12111 5414 12121 5466
rect 12145 5414 12175 5466
rect 12175 5414 12187 5466
rect 12187 5414 12201 5466
rect 12225 5414 12239 5466
rect 12239 5414 12251 5466
rect 12251 5414 12281 5466
rect 12305 5414 12315 5466
rect 12315 5414 12361 5466
rect 12065 5412 12121 5414
rect 12145 5412 12201 5414
rect 12225 5412 12281 5414
rect 12305 5412 12361 5414
rect 12806 6840 12862 6896
rect 12990 6568 13046 6624
rect 12990 5072 13046 5128
rect 12898 4936 12954 4992
rect 12065 4378 12121 4380
rect 12145 4378 12201 4380
rect 12225 4378 12281 4380
rect 12305 4378 12361 4380
rect 12065 4326 12111 4378
rect 12111 4326 12121 4378
rect 12145 4326 12175 4378
rect 12175 4326 12187 4378
rect 12187 4326 12201 4378
rect 12225 4326 12239 4378
rect 12239 4326 12251 4378
rect 12251 4326 12281 4378
rect 12305 4326 12315 4378
rect 12315 4326 12361 4378
rect 12065 4324 12121 4326
rect 12145 4324 12201 4326
rect 12225 4324 12281 4326
rect 12305 4324 12361 4326
rect 13634 6704 13690 6760
rect 13542 6296 13598 6352
rect 14922 15952 14978 16008
rect 14738 15408 14794 15464
rect 14738 13232 14794 13288
rect 15658 17720 15714 17776
rect 16486 20848 16542 20904
rect 19154 21428 19156 21448
rect 19156 21428 19208 21448
rect 19208 21428 19210 21448
rect 18510 21256 18566 21312
rect 19154 21392 19210 21428
rect 15952 20154 16008 20156
rect 16032 20154 16088 20156
rect 16112 20154 16168 20156
rect 16192 20154 16248 20156
rect 15952 20102 15998 20154
rect 15998 20102 16008 20154
rect 16032 20102 16062 20154
rect 16062 20102 16074 20154
rect 16074 20102 16088 20154
rect 16112 20102 16126 20154
rect 16126 20102 16138 20154
rect 16138 20102 16168 20154
rect 16192 20102 16202 20154
rect 16202 20102 16248 20154
rect 15952 20100 16008 20102
rect 16032 20100 16088 20102
rect 16112 20100 16168 20102
rect 16192 20100 16248 20102
rect 15952 19066 16008 19068
rect 16032 19066 16088 19068
rect 16112 19066 16168 19068
rect 16192 19066 16248 19068
rect 15952 19014 15998 19066
rect 15998 19014 16008 19066
rect 16032 19014 16062 19066
rect 16062 19014 16074 19066
rect 16074 19014 16088 19066
rect 16112 19014 16126 19066
rect 16126 19014 16138 19066
rect 16138 19014 16168 19066
rect 16192 19014 16202 19066
rect 16202 19014 16248 19066
rect 15952 19012 16008 19014
rect 16032 19012 16088 19014
rect 16112 19012 16168 19014
rect 16192 19012 16248 19014
rect 15952 17978 16008 17980
rect 16032 17978 16088 17980
rect 16112 17978 16168 17980
rect 16192 17978 16248 17980
rect 15952 17926 15998 17978
rect 15998 17926 16008 17978
rect 16032 17926 16062 17978
rect 16062 17926 16074 17978
rect 16074 17926 16088 17978
rect 16112 17926 16126 17978
rect 16126 17926 16138 17978
rect 16138 17926 16168 17978
rect 16192 17926 16202 17978
rect 16202 17926 16248 17978
rect 15952 17924 16008 17926
rect 16032 17924 16088 17926
rect 16112 17924 16168 17926
rect 16192 17924 16248 17926
rect 15750 15544 15806 15600
rect 15014 12008 15070 12064
rect 15014 11872 15070 11928
rect 14922 11092 14924 11112
rect 14924 11092 14976 11112
rect 14976 11092 14978 11112
rect 14922 11056 14978 11092
rect 15198 12416 15254 12472
rect 14922 10240 14978 10296
rect 16578 19352 16634 19408
rect 16394 18264 16450 18320
rect 16946 20340 16948 20360
rect 16948 20340 17000 20360
rect 17000 20340 17002 20360
rect 16946 20304 17002 20340
rect 16762 19080 16818 19136
rect 16670 18944 16726 19000
rect 17222 19488 17278 19544
rect 17222 19252 17224 19272
rect 17224 19252 17276 19272
rect 17276 19252 17278 19272
rect 17222 19216 17278 19252
rect 17222 18964 17278 19000
rect 17222 18944 17224 18964
rect 17224 18944 17276 18964
rect 17276 18944 17278 18964
rect 16854 18536 16910 18592
rect 16670 18400 16726 18456
rect 16578 18028 16580 18048
rect 16580 18028 16632 18048
rect 16632 18028 16634 18048
rect 16578 17992 16634 18028
rect 16578 17876 16634 17912
rect 16578 17856 16580 17876
rect 16580 17856 16632 17876
rect 16632 17856 16634 17876
rect 15952 16890 16008 16892
rect 16032 16890 16088 16892
rect 16112 16890 16168 16892
rect 16192 16890 16248 16892
rect 15952 16838 15998 16890
rect 15998 16838 16008 16890
rect 16032 16838 16062 16890
rect 16062 16838 16074 16890
rect 16074 16838 16088 16890
rect 16112 16838 16126 16890
rect 16126 16838 16138 16890
rect 16138 16838 16168 16890
rect 16192 16838 16202 16890
rect 16202 16838 16248 16890
rect 15952 16836 16008 16838
rect 16032 16836 16088 16838
rect 16112 16836 16168 16838
rect 16192 16836 16248 16838
rect 16486 16768 16542 16824
rect 16762 17720 16818 17776
rect 17130 17312 17186 17368
rect 17222 17176 17278 17232
rect 16578 16668 16580 16688
rect 16580 16668 16632 16688
rect 16632 16668 16634 16688
rect 16578 16632 16634 16668
rect 15952 15802 16008 15804
rect 16032 15802 16088 15804
rect 16112 15802 16168 15804
rect 16192 15802 16248 15804
rect 15952 15750 15998 15802
rect 15998 15750 16008 15802
rect 16032 15750 16062 15802
rect 16062 15750 16074 15802
rect 16074 15750 16088 15802
rect 16112 15750 16126 15802
rect 16126 15750 16138 15802
rect 16138 15750 16168 15802
rect 16192 15750 16202 15802
rect 16202 15750 16248 15802
rect 15952 15748 16008 15750
rect 16032 15748 16088 15750
rect 16112 15748 16168 15750
rect 16192 15748 16248 15750
rect 16670 16360 16726 16416
rect 15952 14714 16008 14716
rect 16032 14714 16088 14716
rect 16112 14714 16168 14716
rect 16192 14714 16248 14716
rect 15952 14662 15998 14714
rect 15998 14662 16008 14714
rect 16032 14662 16062 14714
rect 16062 14662 16074 14714
rect 16074 14662 16088 14714
rect 16112 14662 16126 14714
rect 16126 14662 16138 14714
rect 16138 14662 16168 14714
rect 16192 14662 16202 14714
rect 16202 14662 16248 14714
rect 15952 14660 16008 14662
rect 16032 14660 16088 14662
rect 16112 14660 16168 14662
rect 16192 14660 16248 14662
rect 16486 13776 16542 13832
rect 15952 13626 16008 13628
rect 16032 13626 16088 13628
rect 16112 13626 16168 13628
rect 16192 13626 16248 13628
rect 15952 13574 15998 13626
rect 15998 13574 16008 13626
rect 16032 13574 16062 13626
rect 16062 13574 16074 13626
rect 16074 13574 16088 13626
rect 16112 13574 16126 13626
rect 16126 13574 16138 13626
rect 16138 13574 16168 13626
rect 16192 13574 16202 13626
rect 16202 13574 16248 13626
rect 15952 13572 16008 13574
rect 16032 13572 16088 13574
rect 16112 13572 16168 13574
rect 16192 13572 16248 13574
rect 16946 16496 17002 16552
rect 16946 15272 17002 15328
rect 17130 15680 17186 15736
rect 16946 14864 17002 14920
rect 17866 20168 17922 20224
rect 17774 19624 17830 19680
rect 17866 18164 17868 18184
rect 17868 18164 17920 18184
rect 17920 18164 17922 18184
rect 17866 18128 17922 18164
rect 17774 17720 17830 17776
rect 17498 16768 17554 16824
rect 17406 15816 17462 15872
rect 17406 15680 17462 15736
rect 17222 14456 17278 14512
rect 15750 12416 15806 12472
rect 15952 12538 16008 12540
rect 16032 12538 16088 12540
rect 16112 12538 16168 12540
rect 16192 12538 16248 12540
rect 15952 12486 15998 12538
rect 15998 12486 16008 12538
rect 16032 12486 16062 12538
rect 16062 12486 16074 12538
rect 16074 12486 16088 12538
rect 16112 12486 16126 12538
rect 16126 12486 16138 12538
rect 16138 12486 16168 12538
rect 16192 12486 16202 12538
rect 16202 12486 16248 12538
rect 15952 12484 16008 12486
rect 16032 12484 16088 12486
rect 16112 12484 16168 12486
rect 16192 12484 16248 12486
rect 15750 12144 15806 12200
rect 15750 11464 15806 11520
rect 15474 11192 15530 11248
rect 15658 11192 15714 11248
rect 15382 10784 15438 10840
rect 15952 11450 16008 11452
rect 16032 11450 16088 11452
rect 16112 11450 16168 11452
rect 16192 11450 16248 11452
rect 15952 11398 15998 11450
rect 15998 11398 16008 11450
rect 16032 11398 16062 11450
rect 16062 11398 16074 11450
rect 16074 11398 16088 11450
rect 16112 11398 16126 11450
rect 16126 11398 16138 11450
rect 16138 11398 16168 11450
rect 16192 11398 16202 11450
rect 16202 11398 16248 11450
rect 15952 11396 16008 11398
rect 16032 11396 16088 11398
rect 16112 11396 16168 11398
rect 16192 11396 16248 11398
rect 14738 10004 14740 10024
rect 14740 10004 14792 10024
rect 14792 10004 14794 10024
rect 14738 9968 14794 10004
rect 14554 9560 14610 9616
rect 14186 9288 14242 9344
rect 13450 5888 13506 5944
rect 13358 5244 13360 5264
rect 13360 5244 13412 5264
rect 13412 5244 13414 5264
rect 13358 5208 13414 5244
rect 14278 6604 14280 6624
rect 14280 6604 14332 6624
rect 14332 6604 14334 6624
rect 14278 6568 14334 6604
rect 15382 9152 15438 9208
rect 14738 6704 14794 6760
rect 14462 6024 14518 6080
rect 13910 4700 13912 4720
rect 13912 4700 13964 4720
rect 13964 4700 13966 4720
rect 13910 4664 13966 4700
rect 12065 3290 12121 3292
rect 12145 3290 12201 3292
rect 12225 3290 12281 3292
rect 12305 3290 12361 3292
rect 12065 3238 12111 3290
rect 12111 3238 12121 3290
rect 12145 3238 12175 3290
rect 12175 3238 12187 3290
rect 12187 3238 12201 3290
rect 12225 3238 12239 3290
rect 12239 3238 12251 3290
rect 12251 3238 12281 3290
rect 12305 3238 12315 3290
rect 12315 3238 12361 3290
rect 12065 3236 12121 3238
rect 12145 3236 12201 3238
rect 12225 3236 12281 3238
rect 12305 3236 12361 3238
rect 14186 4936 14242 4992
rect 16118 10648 16174 10704
rect 15952 10362 16008 10364
rect 16032 10362 16088 10364
rect 16112 10362 16168 10364
rect 16192 10362 16248 10364
rect 15952 10310 15998 10362
rect 15998 10310 16008 10362
rect 16032 10310 16062 10362
rect 16062 10310 16074 10362
rect 16074 10310 16088 10362
rect 16112 10310 16126 10362
rect 16126 10310 16138 10362
rect 16138 10310 16168 10362
rect 16192 10310 16202 10362
rect 16202 10310 16248 10362
rect 15952 10308 16008 10310
rect 16032 10308 16088 10310
rect 16112 10308 16168 10310
rect 16192 10308 16248 10310
rect 16486 12552 16542 12608
rect 16394 11328 16450 11384
rect 15842 9580 15898 9616
rect 15842 9560 15844 9580
rect 15844 9560 15896 9580
rect 15896 9560 15898 9580
rect 15952 9274 16008 9276
rect 16032 9274 16088 9276
rect 16112 9274 16168 9276
rect 16192 9274 16248 9276
rect 15952 9222 15998 9274
rect 15998 9222 16008 9274
rect 16032 9222 16062 9274
rect 16062 9222 16074 9274
rect 16074 9222 16088 9274
rect 16112 9222 16126 9274
rect 16126 9222 16138 9274
rect 16138 9222 16168 9274
rect 16192 9222 16202 9274
rect 16202 9222 16248 9274
rect 15952 9220 16008 9222
rect 16032 9220 16088 9222
rect 16112 9220 16168 9222
rect 16192 9220 16248 9222
rect 15952 8186 16008 8188
rect 16032 8186 16088 8188
rect 16112 8186 16168 8188
rect 16192 8186 16248 8188
rect 15952 8134 15998 8186
rect 15998 8134 16008 8186
rect 16032 8134 16062 8186
rect 16062 8134 16074 8186
rect 16074 8134 16088 8186
rect 16112 8134 16126 8186
rect 16126 8134 16138 8186
rect 16138 8134 16168 8186
rect 16192 8134 16202 8186
rect 16202 8134 16248 8186
rect 15952 8132 16008 8134
rect 16032 8132 16088 8134
rect 16112 8132 16168 8134
rect 16192 8132 16248 8134
rect 16394 8608 16450 8664
rect 16946 13232 17002 13288
rect 16854 12960 16910 13016
rect 16670 12008 16726 12064
rect 16670 11056 16726 11112
rect 19246 20984 19302 21040
rect 18418 20712 18474 20768
rect 18694 19896 18750 19952
rect 18602 19624 18658 19680
rect 18142 17312 18198 17368
rect 17866 16360 17922 16416
rect 17774 15680 17830 15736
rect 17774 14184 17830 14240
rect 17774 14068 17830 14104
rect 17774 14048 17776 14068
rect 17776 14048 17828 14068
rect 17828 14048 17830 14068
rect 17774 13640 17830 13696
rect 18510 18808 18566 18864
rect 18510 17584 18566 17640
rect 18418 16904 18474 16960
rect 18878 19624 18934 19680
rect 19246 20032 19302 20088
rect 19522 20712 19578 20768
rect 19154 18264 19210 18320
rect 18970 17992 19026 18048
rect 18970 17856 19026 17912
rect 18878 16904 18934 16960
rect 19839 20698 19895 20700
rect 19919 20698 19975 20700
rect 19999 20698 20055 20700
rect 20079 20698 20135 20700
rect 19839 20646 19885 20698
rect 19885 20646 19895 20698
rect 19919 20646 19949 20698
rect 19949 20646 19961 20698
rect 19961 20646 19975 20698
rect 19999 20646 20013 20698
rect 20013 20646 20025 20698
rect 20025 20646 20055 20698
rect 20079 20646 20089 20698
rect 20089 20646 20135 20698
rect 19839 20644 19895 20646
rect 19919 20644 19975 20646
rect 19999 20644 20055 20646
rect 20079 20644 20135 20646
rect 19706 19896 19762 19952
rect 19839 19610 19895 19612
rect 19919 19610 19975 19612
rect 19999 19610 20055 19612
rect 20079 19610 20135 19612
rect 19839 19558 19885 19610
rect 19885 19558 19895 19610
rect 19919 19558 19949 19610
rect 19949 19558 19961 19610
rect 19961 19558 19975 19610
rect 19999 19558 20013 19610
rect 20013 19558 20025 19610
rect 20025 19558 20055 19610
rect 20079 19558 20089 19610
rect 20089 19558 20135 19610
rect 19839 19556 19895 19558
rect 19919 19556 19975 19558
rect 19999 19556 20055 19558
rect 20079 19556 20135 19558
rect 19430 18828 19486 18864
rect 19430 18808 19432 18828
rect 19432 18808 19484 18828
rect 19484 18808 19486 18828
rect 19338 18400 19394 18456
rect 20258 18944 20314 19000
rect 20718 20848 20774 20904
rect 21546 20712 21602 20768
rect 21362 20168 21418 20224
rect 21086 20032 21142 20088
rect 20810 19080 20866 19136
rect 20626 18944 20682 19000
rect 19839 18522 19895 18524
rect 19919 18522 19975 18524
rect 19999 18522 20055 18524
rect 20079 18522 20135 18524
rect 19839 18470 19885 18522
rect 19885 18470 19895 18522
rect 19919 18470 19949 18522
rect 19949 18470 19961 18522
rect 19961 18470 19975 18522
rect 19999 18470 20013 18522
rect 20013 18470 20025 18522
rect 20025 18470 20055 18522
rect 20079 18470 20089 18522
rect 20089 18470 20135 18522
rect 19839 18468 19895 18470
rect 19919 18468 19975 18470
rect 19999 18468 20055 18470
rect 20079 18468 20135 18470
rect 20258 18400 20314 18456
rect 19430 17992 19486 18048
rect 19430 17856 19486 17912
rect 19338 17604 19394 17640
rect 19338 17584 19340 17604
rect 19340 17584 19392 17604
rect 19392 17584 19394 17604
rect 18694 15000 18750 15056
rect 18418 14356 18420 14376
rect 18420 14356 18472 14376
rect 18472 14356 18474 14376
rect 18418 14320 18474 14356
rect 18234 13912 18290 13968
rect 18970 15272 19026 15328
rect 17406 13096 17462 13152
rect 17958 13096 18014 13152
rect 17314 12552 17370 12608
rect 17130 11736 17186 11792
rect 17590 11736 17646 11792
rect 19614 17176 19670 17232
rect 20166 18264 20222 18320
rect 19839 17434 19895 17436
rect 19919 17434 19975 17436
rect 19999 17434 20055 17436
rect 20079 17434 20135 17436
rect 19839 17382 19885 17434
rect 19885 17382 19895 17434
rect 19919 17382 19949 17434
rect 19949 17382 19961 17434
rect 19961 17382 19975 17434
rect 19999 17382 20013 17434
rect 20013 17382 20025 17434
rect 20025 17382 20055 17434
rect 20079 17382 20089 17434
rect 20089 17382 20135 17434
rect 19839 17380 19895 17382
rect 19919 17380 19975 17382
rect 19999 17380 20055 17382
rect 20079 17380 20135 17382
rect 19890 17176 19946 17232
rect 20258 17312 20314 17368
rect 19062 14592 19118 14648
rect 19614 16224 19670 16280
rect 19522 15564 19578 15600
rect 19522 15544 19524 15564
rect 19524 15544 19576 15564
rect 19576 15544 19578 15564
rect 19839 16346 19895 16348
rect 19919 16346 19975 16348
rect 19999 16346 20055 16348
rect 20079 16346 20135 16348
rect 19839 16294 19885 16346
rect 19885 16294 19895 16346
rect 19919 16294 19949 16346
rect 19949 16294 19961 16346
rect 19961 16294 19975 16346
rect 19999 16294 20013 16346
rect 20013 16294 20025 16346
rect 20025 16294 20055 16346
rect 20079 16294 20089 16346
rect 20089 16294 20135 16346
rect 19839 16292 19895 16294
rect 19919 16292 19975 16294
rect 19999 16292 20055 16294
rect 20079 16292 20135 16294
rect 20074 15680 20130 15736
rect 19522 14612 19578 14648
rect 19522 14592 19524 14612
rect 19524 14592 19576 14612
rect 19576 14592 19578 14612
rect 19839 15258 19895 15260
rect 19919 15258 19975 15260
rect 19999 15258 20055 15260
rect 20079 15258 20135 15260
rect 19839 15206 19885 15258
rect 19885 15206 19895 15258
rect 19919 15206 19949 15258
rect 19949 15206 19961 15258
rect 19961 15206 19975 15258
rect 19999 15206 20013 15258
rect 20013 15206 20025 15258
rect 20025 15206 20055 15258
rect 20079 15206 20089 15258
rect 20089 15206 20135 15258
rect 19839 15204 19895 15206
rect 19919 15204 19975 15206
rect 19999 15204 20055 15206
rect 20079 15204 20135 15206
rect 19890 14764 19892 14784
rect 19892 14764 19944 14784
rect 19944 14764 19946 14784
rect 19890 14728 19946 14764
rect 19522 14456 19578 14512
rect 19706 14456 19762 14512
rect 18418 12980 18474 13016
rect 18418 12960 18420 12980
rect 18420 12960 18472 12980
rect 18472 12960 18474 12980
rect 17958 12144 18014 12200
rect 19246 12824 19302 12880
rect 18878 11872 18934 11928
rect 18970 11600 19026 11656
rect 18326 11076 18382 11112
rect 18326 11056 18328 11076
rect 18328 11056 18380 11076
rect 18380 11056 18382 11076
rect 18510 10920 18566 10976
rect 18970 10412 18972 10432
rect 18972 10412 19024 10432
rect 19024 10412 19026 10432
rect 18970 10376 19026 10412
rect 18878 10124 18934 10160
rect 18878 10104 18880 10124
rect 18880 10104 18932 10124
rect 18932 10104 18934 10124
rect 16946 8880 17002 8936
rect 15952 7098 16008 7100
rect 16032 7098 16088 7100
rect 16112 7098 16168 7100
rect 16192 7098 16248 7100
rect 15952 7046 15998 7098
rect 15998 7046 16008 7098
rect 16032 7046 16062 7098
rect 16062 7046 16074 7098
rect 16074 7046 16088 7098
rect 16112 7046 16126 7098
rect 16126 7046 16138 7098
rect 16138 7046 16168 7098
rect 16192 7046 16202 7098
rect 16202 7046 16248 7098
rect 15952 7044 16008 7046
rect 16032 7044 16088 7046
rect 16112 7044 16168 7046
rect 16192 7044 16248 7046
rect 14186 2932 14188 2952
rect 14188 2932 14240 2952
rect 14240 2932 14242 2952
rect 14186 2896 14242 2932
rect 15952 6010 16008 6012
rect 16032 6010 16088 6012
rect 16112 6010 16168 6012
rect 16192 6010 16248 6012
rect 15952 5958 15998 6010
rect 15998 5958 16008 6010
rect 16032 5958 16062 6010
rect 16062 5958 16074 6010
rect 16074 5958 16088 6010
rect 16112 5958 16126 6010
rect 16126 5958 16138 6010
rect 16138 5958 16168 6010
rect 16192 5958 16202 6010
rect 16202 5958 16248 6010
rect 15952 5956 16008 5958
rect 16032 5956 16088 5958
rect 16112 5956 16168 5958
rect 16192 5956 16248 5958
rect 16210 5344 16266 5400
rect 15566 5072 15622 5128
rect 15750 5108 15752 5128
rect 15752 5108 15804 5128
rect 15804 5108 15806 5128
rect 15750 5072 15806 5108
rect 15474 4936 15530 4992
rect 15750 4820 15806 4856
rect 15750 4800 15752 4820
rect 15752 4800 15804 4820
rect 15804 4800 15806 4820
rect 15952 4922 16008 4924
rect 16032 4922 16088 4924
rect 16112 4922 16168 4924
rect 16192 4922 16248 4924
rect 15952 4870 15998 4922
rect 15998 4870 16008 4922
rect 16032 4870 16062 4922
rect 16062 4870 16074 4922
rect 16074 4870 16088 4922
rect 16112 4870 16126 4922
rect 16126 4870 16138 4922
rect 16138 4870 16168 4922
rect 16192 4870 16202 4922
rect 16202 4870 16248 4922
rect 15952 4868 16008 4870
rect 16032 4868 16088 4870
rect 16112 4868 16168 4870
rect 16192 4868 16248 4870
rect 15952 3834 16008 3836
rect 16032 3834 16088 3836
rect 16112 3834 16168 3836
rect 16192 3834 16248 3836
rect 15952 3782 15998 3834
rect 15998 3782 16008 3834
rect 16032 3782 16062 3834
rect 16062 3782 16074 3834
rect 16074 3782 16088 3834
rect 16112 3782 16126 3834
rect 16126 3782 16138 3834
rect 16138 3782 16168 3834
rect 16192 3782 16202 3834
rect 16202 3782 16248 3834
rect 15952 3780 16008 3782
rect 16032 3780 16088 3782
rect 16112 3780 16168 3782
rect 16192 3780 16248 3782
rect 16578 6840 16634 6896
rect 16578 6568 16634 6624
rect 16578 4800 16634 4856
rect 16946 6432 17002 6488
rect 18234 7520 18290 7576
rect 19706 14184 19762 14240
rect 19839 14170 19895 14172
rect 19919 14170 19975 14172
rect 19999 14170 20055 14172
rect 20079 14170 20135 14172
rect 19839 14118 19885 14170
rect 19885 14118 19895 14170
rect 19919 14118 19949 14170
rect 19949 14118 19961 14170
rect 19961 14118 19975 14170
rect 19999 14118 20013 14170
rect 20013 14118 20025 14170
rect 20025 14118 20055 14170
rect 20079 14118 20089 14170
rect 20089 14118 20135 14170
rect 19839 14116 19895 14118
rect 19919 14116 19975 14118
rect 19999 14116 20055 14118
rect 20079 14116 20135 14118
rect 19706 13368 19762 13424
rect 20534 17448 20590 17504
rect 20626 17040 20682 17096
rect 20442 16224 20498 16280
rect 20350 15680 20406 15736
rect 20994 16904 21050 16960
rect 20718 15952 20774 16008
rect 20626 15272 20682 15328
rect 20534 15136 20590 15192
rect 20718 14864 20774 14920
rect 19839 13082 19895 13084
rect 19919 13082 19975 13084
rect 19999 13082 20055 13084
rect 20079 13082 20135 13084
rect 19839 13030 19885 13082
rect 19885 13030 19895 13082
rect 19919 13030 19949 13082
rect 19949 13030 19961 13082
rect 19961 13030 19975 13082
rect 19999 13030 20013 13082
rect 20013 13030 20025 13082
rect 20025 13030 20055 13082
rect 20079 13030 20089 13082
rect 20089 13030 20135 13082
rect 19839 13028 19895 13030
rect 19919 13028 19975 13030
rect 19999 13028 20055 13030
rect 20079 13028 20135 13030
rect 20258 13096 20314 13152
rect 20074 12860 20076 12880
rect 20076 12860 20128 12880
rect 20128 12860 20130 12880
rect 20074 12824 20130 12860
rect 20442 12688 20498 12744
rect 19338 10376 19394 10432
rect 19154 9016 19210 9072
rect 19154 8472 19210 8528
rect 19338 7948 19394 7984
rect 19338 7928 19340 7948
rect 19340 7928 19392 7948
rect 19392 7928 19394 7948
rect 18326 5344 18382 5400
rect 18326 5072 18382 5128
rect 15952 2746 16008 2748
rect 16032 2746 16088 2748
rect 16112 2746 16168 2748
rect 16192 2746 16248 2748
rect 15952 2694 15998 2746
rect 15998 2694 16008 2746
rect 16032 2694 16062 2746
rect 16062 2694 16074 2746
rect 16074 2694 16088 2746
rect 16112 2694 16126 2746
rect 16126 2694 16138 2746
rect 16138 2694 16168 2746
rect 16192 2694 16202 2746
rect 16202 2694 16248 2746
rect 15952 2692 16008 2694
rect 16032 2692 16088 2694
rect 16112 2692 16168 2694
rect 16192 2692 16248 2694
rect 4291 2202 4347 2204
rect 4371 2202 4427 2204
rect 4451 2202 4507 2204
rect 4531 2202 4587 2204
rect 4291 2150 4337 2202
rect 4337 2150 4347 2202
rect 4371 2150 4401 2202
rect 4401 2150 4413 2202
rect 4413 2150 4427 2202
rect 4451 2150 4465 2202
rect 4465 2150 4477 2202
rect 4477 2150 4507 2202
rect 4531 2150 4541 2202
rect 4541 2150 4587 2202
rect 4291 2148 4347 2150
rect 4371 2148 4427 2150
rect 4451 2148 4507 2150
rect 4531 2148 4587 2150
rect 12065 2202 12121 2204
rect 12145 2202 12201 2204
rect 12225 2202 12281 2204
rect 12305 2202 12361 2204
rect 12065 2150 12111 2202
rect 12111 2150 12121 2202
rect 12145 2150 12175 2202
rect 12175 2150 12187 2202
rect 12187 2150 12201 2202
rect 12225 2150 12239 2202
rect 12239 2150 12251 2202
rect 12251 2150 12281 2202
rect 12305 2150 12315 2202
rect 12315 2150 12361 2202
rect 12065 2148 12121 2150
rect 12145 2148 12201 2150
rect 12225 2148 12281 2150
rect 12305 2148 12361 2150
rect 8178 1658 8234 1660
rect 8258 1658 8314 1660
rect 8338 1658 8394 1660
rect 8418 1658 8474 1660
rect 8178 1606 8224 1658
rect 8224 1606 8234 1658
rect 8258 1606 8288 1658
rect 8288 1606 8300 1658
rect 8300 1606 8314 1658
rect 8338 1606 8352 1658
rect 8352 1606 8364 1658
rect 8364 1606 8394 1658
rect 8418 1606 8428 1658
rect 8428 1606 8474 1658
rect 8178 1604 8234 1606
rect 8258 1604 8314 1606
rect 8338 1604 8394 1606
rect 8418 1604 8474 1606
rect 20166 12300 20222 12336
rect 20166 12280 20168 12300
rect 20168 12280 20220 12300
rect 20220 12280 20222 12300
rect 19839 11994 19895 11996
rect 19919 11994 19975 11996
rect 19999 11994 20055 11996
rect 20079 11994 20135 11996
rect 19839 11942 19885 11994
rect 19885 11942 19895 11994
rect 19919 11942 19949 11994
rect 19949 11942 19961 11994
rect 19961 11942 19975 11994
rect 19999 11942 20013 11994
rect 20013 11942 20025 11994
rect 20025 11942 20055 11994
rect 20079 11942 20089 11994
rect 20089 11942 20135 11994
rect 19839 11940 19895 11942
rect 19919 11940 19975 11942
rect 19999 11940 20055 11942
rect 20079 11940 20135 11942
rect 20350 11872 20406 11928
rect 19798 11600 19854 11656
rect 20442 11328 20498 11384
rect 20810 12280 20866 12336
rect 21362 19896 21418 19952
rect 21546 20168 21602 20224
rect 21362 19624 21418 19680
rect 21270 18400 21326 18456
rect 21454 19488 21510 19544
rect 21914 19488 21970 19544
rect 21454 18944 21510 19000
rect 21362 17584 21418 17640
rect 21270 16496 21326 16552
rect 21178 15816 21234 15872
rect 21638 17584 21694 17640
rect 21546 16360 21602 16416
rect 21546 15816 21602 15872
rect 23386 21256 23442 21312
rect 22282 20168 22338 20224
rect 22834 21004 22890 21040
rect 23726 21242 23782 21244
rect 23806 21242 23862 21244
rect 23886 21242 23942 21244
rect 23966 21242 24022 21244
rect 23726 21190 23772 21242
rect 23772 21190 23782 21242
rect 23806 21190 23836 21242
rect 23836 21190 23848 21242
rect 23848 21190 23862 21242
rect 23886 21190 23900 21242
rect 23900 21190 23912 21242
rect 23912 21190 23942 21242
rect 23966 21190 23976 21242
rect 23976 21190 24022 21242
rect 23726 21188 23782 21190
rect 23806 21188 23862 21190
rect 23886 21188 23942 21190
rect 23966 21188 24022 21190
rect 22834 20984 22836 21004
rect 22836 20984 22888 21004
rect 22888 20984 22890 21004
rect 22742 19760 22798 19816
rect 21914 16496 21970 16552
rect 22282 17076 22284 17096
rect 22284 17076 22336 17096
rect 22336 17076 22338 17096
rect 22282 17040 22338 17076
rect 23294 20440 23350 20496
rect 23110 20304 23166 20360
rect 23018 19796 23020 19816
rect 23020 19796 23072 19816
rect 23072 19796 23074 19816
rect 23018 19760 23074 19796
rect 23754 20440 23810 20496
rect 23726 20154 23782 20156
rect 23806 20154 23862 20156
rect 23886 20154 23942 20156
rect 23966 20154 24022 20156
rect 23726 20102 23772 20154
rect 23772 20102 23782 20154
rect 23806 20102 23836 20154
rect 23836 20102 23848 20154
rect 23848 20102 23862 20154
rect 23886 20102 23900 20154
rect 23900 20102 23912 20154
rect 23912 20102 23942 20154
rect 23966 20102 23976 20154
rect 23976 20102 24022 20154
rect 23726 20100 23782 20102
rect 23806 20100 23862 20102
rect 23886 20100 23942 20102
rect 23966 20100 24022 20102
rect 23478 19488 23534 19544
rect 23202 19080 23258 19136
rect 22926 18264 22982 18320
rect 22650 17992 22706 18048
rect 22558 17040 22614 17096
rect 22282 16768 22338 16824
rect 22006 15000 22062 15056
rect 21822 14320 21878 14376
rect 19706 11092 19708 11112
rect 19708 11092 19760 11112
rect 19760 11092 19762 11112
rect 19706 11056 19762 11092
rect 19839 10906 19895 10908
rect 19919 10906 19975 10908
rect 19999 10906 20055 10908
rect 20079 10906 20135 10908
rect 19839 10854 19885 10906
rect 19885 10854 19895 10906
rect 19919 10854 19949 10906
rect 19949 10854 19961 10906
rect 19961 10854 19975 10906
rect 19999 10854 20013 10906
rect 20013 10854 20025 10906
rect 20025 10854 20055 10906
rect 20079 10854 20089 10906
rect 20089 10854 20135 10906
rect 19839 10852 19895 10854
rect 19919 10852 19975 10854
rect 19999 10852 20055 10854
rect 20079 10852 20135 10854
rect 20442 10512 20498 10568
rect 19839 9818 19895 9820
rect 19919 9818 19975 9820
rect 19999 9818 20055 9820
rect 20079 9818 20135 9820
rect 19839 9766 19885 9818
rect 19885 9766 19895 9818
rect 19919 9766 19949 9818
rect 19949 9766 19961 9818
rect 19961 9766 19975 9818
rect 19999 9766 20013 9818
rect 20013 9766 20025 9818
rect 20025 9766 20055 9818
rect 20079 9766 20089 9818
rect 20089 9766 20135 9818
rect 19839 9764 19895 9766
rect 19919 9764 19975 9766
rect 19999 9764 20055 9766
rect 20079 9764 20135 9766
rect 19839 8730 19895 8732
rect 19919 8730 19975 8732
rect 19999 8730 20055 8732
rect 20079 8730 20135 8732
rect 19839 8678 19885 8730
rect 19885 8678 19895 8730
rect 19919 8678 19949 8730
rect 19949 8678 19961 8730
rect 19961 8678 19975 8730
rect 19999 8678 20013 8730
rect 20013 8678 20025 8730
rect 20025 8678 20055 8730
rect 20079 8678 20089 8730
rect 20089 8678 20135 8730
rect 19839 8676 19895 8678
rect 19919 8676 19975 8678
rect 19999 8676 20055 8678
rect 20079 8676 20135 8678
rect 19798 8492 19854 8528
rect 19798 8472 19800 8492
rect 19800 8472 19852 8492
rect 19852 8472 19854 8492
rect 19246 6024 19302 6080
rect 20902 9968 20958 10024
rect 20626 9560 20682 9616
rect 20534 9016 20590 9072
rect 20258 7792 20314 7848
rect 19839 7642 19895 7644
rect 19919 7642 19975 7644
rect 19999 7642 20055 7644
rect 20079 7642 20135 7644
rect 19839 7590 19885 7642
rect 19885 7590 19895 7642
rect 19919 7590 19949 7642
rect 19949 7590 19961 7642
rect 19961 7590 19975 7642
rect 19999 7590 20013 7642
rect 20013 7590 20025 7642
rect 20025 7590 20055 7642
rect 20079 7590 20089 7642
rect 20089 7590 20135 7642
rect 19839 7588 19895 7590
rect 19919 7588 19975 7590
rect 19999 7588 20055 7590
rect 20079 7588 20135 7590
rect 20166 7112 20222 7168
rect 19839 6554 19895 6556
rect 19919 6554 19975 6556
rect 19999 6554 20055 6556
rect 20079 6554 20135 6556
rect 19839 6502 19885 6554
rect 19885 6502 19895 6554
rect 19919 6502 19949 6554
rect 19949 6502 19961 6554
rect 19961 6502 19975 6554
rect 19999 6502 20013 6554
rect 20013 6502 20025 6554
rect 20025 6502 20055 6554
rect 20079 6502 20089 6554
rect 20089 6502 20135 6554
rect 19839 6500 19895 6502
rect 19919 6500 19975 6502
rect 19999 6500 20055 6502
rect 20079 6500 20135 6502
rect 19338 5752 19394 5808
rect 19839 5466 19895 5468
rect 19919 5466 19975 5468
rect 19999 5466 20055 5468
rect 20079 5466 20135 5468
rect 19839 5414 19885 5466
rect 19885 5414 19895 5466
rect 19919 5414 19949 5466
rect 19949 5414 19961 5466
rect 19961 5414 19975 5466
rect 19999 5414 20013 5466
rect 20013 5414 20025 5466
rect 20025 5414 20055 5466
rect 20079 5414 20089 5466
rect 20089 5414 20135 5466
rect 19839 5412 19895 5414
rect 19919 5412 19975 5414
rect 19999 5412 20055 5414
rect 20079 5412 20135 5414
rect 19839 4378 19895 4380
rect 19919 4378 19975 4380
rect 19999 4378 20055 4380
rect 20079 4378 20135 4380
rect 19839 4326 19885 4378
rect 19885 4326 19895 4378
rect 19919 4326 19949 4378
rect 19949 4326 19961 4378
rect 19961 4326 19975 4378
rect 19999 4326 20013 4378
rect 20013 4326 20025 4378
rect 20025 4326 20055 4378
rect 20079 4326 20089 4378
rect 20089 4326 20135 4378
rect 19839 4324 19895 4326
rect 19919 4324 19975 4326
rect 19999 4324 20055 4326
rect 20079 4324 20135 4326
rect 20534 8064 20590 8120
rect 20442 7112 20498 7168
rect 21178 9832 21234 9888
rect 20718 7692 20720 7712
rect 20720 7692 20772 7712
rect 20772 7692 20774 7712
rect 20718 7656 20774 7692
rect 20534 6976 20590 7032
rect 20442 4120 20498 4176
rect 19839 3290 19895 3292
rect 19919 3290 19975 3292
rect 19999 3290 20055 3292
rect 20079 3290 20135 3292
rect 19839 3238 19885 3290
rect 19885 3238 19895 3290
rect 19919 3238 19949 3290
rect 19949 3238 19961 3290
rect 19961 3238 19975 3290
rect 19999 3238 20013 3290
rect 20013 3238 20025 3290
rect 20025 3238 20055 3290
rect 20079 3238 20089 3290
rect 20089 3238 20135 3290
rect 19839 3236 19895 3238
rect 19919 3236 19975 3238
rect 19999 3236 20055 3238
rect 20079 3236 20135 3238
rect 22006 14048 22062 14104
rect 22006 13932 22062 13968
rect 22006 13912 22008 13932
rect 22008 13912 22060 13932
rect 22060 13912 22062 13932
rect 23294 17584 23350 17640
rect 22834 15408 22890 15464
rect 22834 15000 22890 15056
rect 22282 13776 22338 13832
rect 22742 14456 22798 14512
rect 22558 13368 22614 13424
rect 22006 13096 22062 13152
rect 21730 12280 21786 12336
rect 21730 12044 21732 12064
rect 21732 12044 21784 12064
rect 21784 12044 21786 12064
rect 21730 12008 21786 12044
rect 21362 11464 21418 11520
rect 21914 11212 21970 11248
rect 21914 11192 21916 11212
rect 21916 11192 21968 11212
rect 21968 11192 21970 11212
rect 21362 9560 21418 9616
rect 21362 5208 21418 5264
rect 21270 4020 21272 4040
rect 21272 4020 21324 4040
rect 21324 4020 21326 4040
rect 21270 3984 21326 4020
rect 20994 3596 21050 3632
rect 20994 3576 20996 3596
rect 20996 3576 21048 3596
rect 21048 3576 21050 3596
rect 22742 12688 22798 12744
rect 23726 19066 23782 19068
rect 23806 19066 23862 19068
rect 23886 19066 23942 19068
rect 23966 19066 24022 19068
rect 23726 19014 23772 19066
rect 23772 19014 23782 19066
rect 23806 19014 23836 19066
rect 23836 19014 23848 19066
rect 23848 19014 23862 19066
rect 23886 19014 23900 19066
rect 23900 19014 23912 19066
rect 23912 19014 23942 19066
rect 23966 19014 23976 19066
rect 23976 19014 24022 19066
rect 23726 19012 23782 19014
rect 23806 19012 23862 19014
rect 23886 19012 23942 19014
rect 23966 19012 24022 19014
rect 23726 17978 23782 17980
rect 23806 17978 23862 17980
rect 23886 17978 23942 17980
rect 23966 17978 24022 17980
rect 23726 17926 23772 17978
rect 23772 17926 23782 17978
rect 23806 17926 23836 17978
rect 23836 17926 23848 17978
rect 23848 17926 23862 17978
rect 23886 17926 23900 17978
rect 23900 17926 23912 17978
rect 23912 17926 23942 17978
rect 23966 17926 23976 17978
rect 23976 17926 24022 17978
rect 23726 17924 23782 17926
rect 23806 17924 23862 17926
rect 23886 17924 23942 17926
rect 23966 17924 24022 17926
rect 23570 17856 23626 17912
rect 23386 15700 23442 15736
rect 23386 15680 23388 15700
rect 23388 15680 23440 15700
rect 23440 15680 23442 15700
rect 23386 15544 23442 15600
rect 23294 14456 23350 14512
rect 24306 17856 24362 17912
rect 24214 17448 24270 17504
rect 24030 17176 24086 17232
rect 23726 16890 23782 16892
rect 23806 16890 23862 16892
rect 23886 16890 23942 16892
rect 23966 16890 24022 16892
rect 23726 16838 23772 16890
rect 23772 16838 23782 16890
rect 23806 16838 23836 16890
rect 23836 16838 23848 16890
rect 23848 16838 23862 16890
rect 23886 16838 23900 16890
rect 23900 16838 23912 16890
rect 23912 16838 23942 16890
rect 23966 16838 23976 16890
rect 23976 16838 24022 16890
rect 23726 16836 23782 16838
rect 23806 16836 23862 16838
rect 23886 16836 23942 16838
rect 23966 16836 24022 16838
rect 24122 16768 24178 16824
rect 23938 16496 23994 16552
rect 23570 15816 23626 15872
rect 23726 15802 23782 15804
rect 23806 15802 23862 15804
rect 23886 15802 23942 15804
rect 23966 15802 24022 15804
rect 23726 15750 23772 15802
rect 23772 15750 23782 15802
rect 23806 15750 23836 15802
rect 23836 15750 23848 15802
rect 23848 15750 23862 15802
rect 23886 15750 23900 15802
rect 23900 15750 23912 15802
rect 23912 15750 23942 15802
rect 23966 15750 23976 15802
rect 23976 15750 24022 15802
rect 23726 15748 23782 15750
rect 23806 15748 23862 15750
rect 23886 15748 23942 15750
rect 23966 15748 24022 15750
rect 23726 14714 23782 14716
rect 23806 14714 23862 14716
rect 23886 14714 23942 14716
rect 23966 14714 24022 14716
rect 23726 14662 23772 14714
rect 23772 14662 23782 14714
rect 23806 14662 23836 14714
rect 23836 14662 23848 14714
rect 23848 14662 23862 14714
rect 23886 14662 23900 14714
rect 23900 14662 23912 14714
rect 23912 14662 23942 14714
rect 23966 14662 23976 14714
rect 23976 14662 24022 14714
rect 23726 14660 23782 14662
rect 23806 14660 23862 14662
rect 23886 14660 23942 14662
rect 23966 14660 24022 14662
rect 23938 14048 23994 14104
rect 23726 13626 23782 13628
rect 23806 13626 23862 13628
rect 23886 13626 23942 13628
rect 23966 13626 24022 13628
rect 23726 13574 23772 13626
rect 23772 13574 23782 13626
rect 23806 13574 23836 13626
rect 23836 13574 23848 13626
rect 23848 13574 23862 13626
rect 23886 13574 23900 13626
rect 23900 13574 23912 13626
rect 23912 13574 23942 13626
rect 23966 13574 23976 13626
rect 23976 13574 24022 13626
rect 23726 13572 23782 13574
rect 23806 13572 23862 13574
rect 23886 13572 23942 13574
rect 23966 13572 24022 13574
rect 26054 21936 26110 21992
rect 24674 21800 24730 21856
rect 24674 20712 24730 20768
rect 26606 21800 26662 21856
rect 25410 21004 25466 21040
rect 25410 20984 25412 21004
rect 25412 20984 25464 21004
rect 25464 20984 25466 21004
rect 24766 19488 24822 19544
rect 24950 18708 24952 18728
rect 24952 18708 25004 18728
rect 25004 18708 25006 18728
rect 24950 18672 25006 18708
rect 24674 18148 24730 18184
rect 24674 18128 24676 18148
rect 24676 18128 24728 18148
rect 24728 18128 24730 18148
rect 24858 17740 24914 17776
rect 24858 17720 24860 17740
rect 24860 17720 24912 17740
rect 24912 17720 24914 17740
rect 24858 17312 24914 17368
rect 24214 15272 24270 15328
rect 24214 14728 24270 14784
rect 24490 15272 24546 15328
rect 24858 14864 24914 14920
rect 24398 13796 24454 13832
rect 24398 13776 24400 13796
rect 24400 13776 24452 13796
rect 24452 13776 24454 13796
rect 22650 12144 22706 12200
rect 22834 11600 22890 11656
rect 21730 7792 21786 7848
rect 22374 7948 22430 7984
rect 22374 7928 22376 7948
rect 22376 7928 22428 7948
rect 22428 7928 22430 7948
rect 21822 6568 21878 6624
rect 22006 6432 22062 6488
rect 22098 5072 22154 5128
rect 20074 2896 20130 2952
rect 21454 3304 21510 3360
rect 21914 3984 21970 4040
rect 22834 9560 22890 9616
rect 23110 9560 23166 9616
rect 22742 8064 22798 8120
rect 22466 6060 22468 6080
rect 22468 6060 22520 6080
rect 22520 6060 22522 6080
rect 22466 6024 22522 6060
rect 22650 6840 22706 6896
rect 23726 12538 23782 12540
rect 23806 12538 23862 12540
rect 23886 12538 23942 12540
rect 23966 12538 24022 12540
rect 23726 12486 23772 12538
rect 23772 12486 23782 12538
rect 23806 12486 23836 12538
rect 23836 12486 23848 12538
rect 23848 12486 23862 12538
rect 23886 12486 23900 12538
rect 23900 12486 23912 12538
rect 23912 12486 23942 12538
rect 23966 12486 23976 12538
rect 23976 12486 24022 12538
rect 23726 12484 23782 12486
rect 23806 12484 23862 12486
rect 23886 12484 23942 12486
rect 23966 12484 24022 12486
rect 23754 12300 23810 12336
rect 23754 12280 23756 12300
rect 23756 12280 23808 12300
rect 23808 12280 23810 12300
rect 23754 12008 23810 12064
rect 24306 13232 24362 13288
rect 24490 12688 24546 12744
rect 25318 16940 25320 16960
rect 25320 16940 25372 16960
rect 25372 16940 25374 16960
rect 25318 16904 25374 16940
rect 25226 16768 25282 16824
rect 25502 16088 25558 16144
rect 25318 15408 25374 15464
rect 23726 11450 23782 11452
rect 23806 11450 23862 11452
rect 23886 11450 23942 11452
rect 23966 11450 24022 11452
rect 23726 11398 23772 11450
rect 23772 11398 23782 11450
rect 23806 11398 23836 11450
rect 23836 11398 23848 11450
rect 23848 11398 23862 11450
rect 23886 11398 23900 11450
rect 23900 11398 23912 11450
rect 23912 11398 23942 11450
rect 23966 11398 23976 11450
rect 23976 11398 24022 11450
rect 23726 11396 23782 11398
rect 23806 11396 23862 11398
rect 23886 11396 23942 11398
rect 23966 11396 24022 11398
rect 23726 10362 23782 10364
rect 23806 10362 23862 10364
rect 23886 10362 23942 10364
rect 23966 10362 24022 10364
rect 23726 10310 23772 10362
rect 23772 10310 23782 10362
rect 23806 10310 23836 10362
rect 23836 10310 23848 10362
rect 23848 10310 23862 10362
rect 23886 10310 23900 10362
rect 23900 10310 23912 10362
rect 23912 10310 23942 10362
rect 23966 10310 23976 10362
rect 23976 10310 24022 10362
rect 23726 10308 23782 10310
rect 23806 10308 23862 10310
rect 23886 10308 23942 10310
rect 23966 10308 24022 10310
rect 24766 12416 24822 12472
rect 25226 14320 25282 14376
rect 25318 13776 25374 13832
rect 25686 15036 25688 15056
rect 25688 15036 25740 15056
rect 25740 15036 25742 15056
rect 25686 15000 25742 15036
rect 25870 15136 25926 15192
rect 25686 12416 25742 12472
rect 24858 11736 24914 11792
rect 24582 11056 24638 11112
rect 23662 10004 23664 10024
rect 23664 10004 23716 10024
rect 23716 10004 23718 10024
rect 23662 9968 23718 10004
rect 24214 9968 24270 10024
rect 23202 8492 23258 8528
rect 23202 8472 23204 8492
rect 23204 8472 23256 8492
rect 23256 8472 23258 8492
rect 23726 9274 23782 9276
rect 23806 9274 23862 9276
rect 23886 9274 23942 9276
rect 23966 9274 24022 9276
rect 23726 9222 23772 9274
rect 23772 9222 23782 9274
rect 23806 9222 23836 9274
rect 23836 9222 23848 9274
rect 23848 9222 23862 9274
rect 23886 9222 23900 9274
rect 23900 9222 23912 9274
rect 23912 9222 23942 9274
rect 23966 9222 23976 9274
rect 23976 9222 24022 9274
rect 23726 9220 23782 9222
rect 23806 9220 23862 9222
rect 23886 9220 23942 9222
rect 23966 9220 24022 9222
rect 24398 9832 24454 9888
rect 24950 10648 25006 10704
rect 24214 8880 24270 8936
rect 23726 8186 23782 8188
rect 23806 8186 23862 8188
rect 23886 8186 23942 8188
rect 23966 8186 24022 8188
rect 23726 8134 23772 8186
rect 23772 8134 23782 8186
rect 23806 8134 23836 8186
rect 23836 8134 23848 8186
rect 23848 8134 23862 8186
rect 23886 8134 23900 8186
rect 23900 8134 23912 8186
rect 23912 8134 23942 8186
rect 23966 8134 23976 8186
rect 23976 8134 24022 8186
rect 23726 8132 23782 8134
rect 23806 8132 23862 8134
rect 23886 8132 23942 8134
rect 23966 8132 24022 8134
rect 23386 7656 23442 7712
rect 22834 6704 22890 6760
rect 23726 7098 23782 7100
rect 23806 7098 23862 7100
rect 23886 7098 23942 7100
rect 23966 7098 24022 7100
rect 23726 7046 23772 7098
rect 23772 7046 23782 7098
rect 23806 7046 23836 7098
rect 23836 7046 23848 7098
rect 23848 7046 23862 7098
rect 23886 7046 23900 7098
rect 23900 7046 23912 7098
rect 23912 7046 23942 7098
rect 23966 7046 23976 7098
rect 23976 7046 24022 7098
rect 23726 7044 23782 7046
rect 23806 7044 23862 7046
rect 23886 7044 23942 7046
rect 23966 7044 24022 7046
rect 24858 9052 24860 9072
rect 24860 9052 24912 9072
rect 24912 9052 24914 9072
rect 24858 9016 24914 9052
rect 24122 6704 24178 6760
rect 24030 6296 24086 6352
rect 23726 6010 23782 6012
rect 23806 6010 23862 6012
rect 23886 6010 23942 6012
rect 23966 6010 24022 6012
rect 23726 5958 23772 6010
rect 23772 5958 23782 6010
rect 23806 5958 23836 6010
rect 23836 5958 23848 6010
rect 23848 5958 23862 6010
rect 23886 5958 23900 6010
rect 23900 5958 23912 6010
rect 23912 5958 23942 6010
rect 23966 5958 23976 6010
rect 23976 5958 24022 6010
rect 23726 5956 23782 5958
rect 23806 5956 23862 5958
rect 23886 5956 23942 5958
rect 23966 5956 24022 5958
rect 25594 9832 25650 9888
rect 29734 21936 29790 21992
rect 28078 21800 28134 21856
rect 27613 21786 27669 21788
rect 27693 21786 27749 21788
rect 27773 21786 27829 21788
rect 27853 21786 27909 21788
rect 27613 21734 27659 21786
rect 27659 21734 27669 21786
rect 27693 21734 27723 21786
rect 27723 21734 27735 21786
rect 27735 21734 27749 21786
rect 27773 21734 27787 21786
rect 27787 21734 27799 21786
rect 27799 21734 27829 21786
rect 27853 21734 27863 21786
rect 27863 21734 27909 21786
rect 27613 21732 27669 21734
rect 27693 21732 27749 21734
rect 27773 21732 27829 21734
rect 27853 21732 27909 21734
rect 27434 21664 27490 21720
rect 27710 21528 27766 21584
rect 26330 19624 26386 19680
rect 26238 17040 26294 17096
rect 26054 15272 26110 15328
rect 26698 19352 26754 19408
rect 26606 17584 26662 17640
rect 26330 16360 26386 16416
rect 26422 15680 26478 15736
rect 26422 14184 26478 14240
rect 27066 19488 27122 19544
rect 26974 19352 27030 19408
rect 27342 19760 27398 19816
rect 26974 16904 27030 16960
rect 27066 16224 27122 16280
rect 27158 14728 27214 14784
rect 26974 14048 27030 14104
rect 26514 13912 26570 13968
rect 26330 12280 26386 12336
rect 27066 13268 27068 13288
rect 27068 13268 27120 13288
rect 27120 13268 27122 13288
rect 27066 13232 27122 13268
rect 26606 11872 26662 11928
rect 26514 10512 26570 10568
rect 26054 9832 26110 9888
rect 26238 9424 26294 9480
rect 25962 7928 26018 7984
rect 25870 7792 25926 7848
rect 24398 6024 24454 6080
rect 24214 5888 24270 5944
rect 25226 7248 25282 7304
rect 24950 6196 24952 6216
rect 24952 6196 25004 6216
rect 25004 6196 25006 6216
rect 22374 4800 22430 4856
rect 24306 5652 24308 5672
rect 24308 5652 24360 5672
rect 24360 5652 24362 5672
rect 24306 5616 24362 5652
rect 23938 5072 23994 5128
rect 23726 4922 23782 4924
rect 23806 4922 23862 4924
rect 23886 4922 23942 4924
rect 23966 4922 24022 4924
rect 23726 4870 23772 4922
rect 23772 4870 23782 4922
rect 23806 4870 23836 4922
rect 23836 4870 23848 4922
rect 23848 4870 23862 4922
rect 23886 4870 23900 4922
rect 23900 4870 23912 4922
rect 23912 4870 23942 4922
rect 23966 4870 23976 4922
rect 23976 4870 24022 4922
rect 23726 4868 23782 4870
rect 23806 4868 23862 4870
rect 23886 4868 23942 4870
rect 23966 4868 24022 4870
rect 23478 4664 23534 4720
rect 21730 3052 21786 3088
rect 21730 3032 21732 3052
rect 21732 3032 21784 3052
rect 21784 3032 21786 3052
rect 15952 1658 16008 1660
rect 16032 1658 16088 1660
rect 16112 1658 16168 1660
rect 16192 1658 16248 1660
rect 15952 1606 15998 1658
rect 15998 1606 16008 1658
rect 16032 1606 16062 1658
rect 16062 1606 16074 1658
rect 16074 1606 16088 1658
rect 16112 1606 16126 1658
rect 16126 1606 16138 1658
rect 16138 1606 16168 1658
rect 16192 1606 16202 1658
rect 16202 1606 16248 1658
rect 15952 1604 16008 1606
rect 16032 1604 16088 1606
rect 16112 1604 16168 1606
rect 16192 1604 16248 1606
rect 19839 2202 19895 2204
rect 19919 2202 19975 2204
rect 19999 2202 20055 2204
rect 20079 2202 20135 2204
rect 19839 2150 19885 2202
rect 19885 2150 19895 2202
rect 19919 2150 19949 2202
rect 19949 2150 19961 2202
rect 19961 2150 19975 2202
rect 19999 2150 20013 2202
rect 20013 2150 20025 2202
rect 20025 2150 20055 2202
rect 20079 2150 20089 2202
rect 20089 2150 20135 2202
rect 19839 2148 19895 2150
rect 19919 2148 19975 2150
rect 19999 2148 20055 2150
rect 20079 2148 20135 2150
rect 23018 3984 23074 4040
rect 23294 4020 23296 4040
rect 23296 4020 23348 4040
rect 23348 4020 23350 4040
rect 23294 3984 23350 4020
rect 23726 3834 23782 3836
rect 23806 3834 23862 3836
rect 23886 3834 23942 3836
rect 23966 3834 24022 3836
rect 23726 3782 23772 3834
rect 23772 3782 23782 3834
rect 23806 3782 23836 3834
rect 23836 3782 23848 3834
rect 23848 3782 23862 3834
rect 23886 3782 23900 3834
rect 23900 3782 23912 3834
rect 23912 3782 23942 3834
rect 23966 3782 23976 3834
rect 23976 3782 24022 3834
rect 23726 3780 23782 3782
rect 23806 3780 23862 3782
rect 23886 3780 23942 3782
rect 23966 3780 24022 3782
rect 24030 3440 24086 3496
rect 24398 4120 24454 4176
rect 24950 6160 25006 6196
rect 25594 6704 25650 6760
rect 25410 6568 25466 6624
rect 25502 6296 25558 6352
rect 24858 5772 24914 5808
rect 24858 5752 24860 5772
rect 24860 5752 24912 5772
rect 24912 5752 24914 5772
rect 24766 4528 24822 4584
rect 23726 2746 23782 2748
rect 23806 2746 23862 2748
rect 23886 2746 23942 2748
rect 23966 2746 24022 2748
rect 23726 2694 23772 2746
rect 23772 2694 23782 2746
rect 23806 2694 23836 2746
rect 23836 2694 23848 2746
rect 23848 2694 23862 2746
rect 23886 2694 23900 2746
rect 23900 2694 23912 2746
rect 23912 2694 23942 2746
rect 23966 2694 23976 2746
rect 23976 2694 24022 2746
rect 23726 2692 23782 2694
rect 23806 2692 23862 2694
rect 23886 2692 23942 2694
rect 23966 2692 24022 2694
rect 24674 3052 24730 3088
rect 24674 3032 24676 3052
rect 24676 3032 24728 3052
rect 24728 3032 24730 3052
rect 25226 5208 25282 5264
rect 25042 3984 25098 4040
rect 24858 3304 24914 3360
rect 25134 3712 25190 3768
rect 25686 6432 25742 6488
rect 27613 20698 27669 20700
rect 27693 20698 27749 20700
rect 27773 20698 27829 20700
rect 27853 20698 27909 20700
rect 27613 20646 27659 20698
rect 27659 20646 27669 20698
rect 27693 20646 27723 20698
rect 27723 20646 27735 20698
rect 27735 20646 27749 20698
rect 27773 20646 27787 20698
rect 27787 20646 27799 20698
rect 27799 20646 27829 20698
rect 27853 20646 27863 20698
rect 27863 20646 27909 20698
rect 27613 20644 27669 20646
rect 27693 20644 27749 20646
rect 27773 20644 27829 20646
rect 27853 20644 27909 20646
rect 27613 19610 27669 19612
rect 27693 19610 27749 19612
rect 27773 19610 27829 19612
rect 27853 19610 27909 19612
rect 27613 19558 27659 19610
rect 27659 19558 27669 19610
rect 27693 19558 27723 19610
rect 27723 19558 27735 19610
rect 27735 19558 27749 19610
rect 27773 19558 27787 19610
rect 27787 19558 27799 19610
rect 27799 19558 27829 19610
rect 27853 19558 27863 19610
rect 27863 19558 27909 19610
rect 27613 19556 27669 19558
rect 27693 19556 27749 19558
rect 27773 19556 27829 19558
rect 27853 19556 27909 19558
rect 27613 18522 27669 18524
rect 27693 18522 27749 18524
rect 27773 18522 27829 18524
rect 27853 18522 27909 18524
rect 27613 18470 27659 18522
rect 27659 18470 27669 18522
rect 27693 18470 27723 18522
rect 27723 18470 27735 18522
rect 27735 18470 27749 18522
rect 27773 18470 27787 18522
rect 27787 18470 27799 18522
rect 27799 18470 27829 18522
rect 27853 18470 27863 18522
rect 27863 18470 27909 18522
rect 27613 18468 27669 18470
rect 27693 18468 27749 18470
rect 27773 18468 27829 18470
rect 27853 18468 27909 18470
rect 27802 18264 27858 18320
rect 27613 17434 27669 17436
rect 27693 17434 27749 17436
rect 27773 17434 27829 17436
rect 27853 17434 27909 17436
rect 27613 17382 27659 17434
rect 27659 17382 27669 17434
rect 27693 17382 27723 17434
rect 27723 17382 27735 17434
rect 27735 17382 27749 17434
rect 27773 17382 27787 17434
rect 27787 17382 27799 17434
rect 27799 17382 27829 17434
rect 27853 17382 27863 17434
rect 27863 17382 27909 17434
rect 27613 17380 27669 17382
rect 27693 17380 27749 17382
rect 27773 17380 27829 17382
rect 27853 17380 27909 17382
rect 30010 21800 30066 21856
rect 30286 21800 30342 21856
rect 27613 16346 27669 16348
rect 27693 16346 27749 16348
rect 27773 16346 27829 16348
rect 27853 16346 27909 16348
rect 27613 16294 27659 16346
rect 27659 16294 27669 16346
rect 27693 16294 27723 16346
rect 27723 16294 27735 16346
rect 27735 16294 27749 16346
rect 27773 16294 27787 16346
rect 27787 16294 27799 16346
rect 27799 16294 27829 16346
rect 27853 16294 27863 16346
rect 27863 16294 27909 16346
rect 27613 16292 27669 16294
rect 27693 16292 27749 16294
rect 27773 16292 27829 16294
rect 27853 16292 27909 16294
rect 27710 15680 27766 15736
rect 28354 18128 28410 18184
rect 27613 15258 27669 15260
rect 27693 15258 27749 15260
rect 27773 15258 27829 15260
rect 27853 15258 27909 15260
rect 27613 15206 27659 15258
rect 27659 15206 27669 15258
rect 27693 15206 27723 15258
rect 27723 15206 27735 15258
rect 27735 15206 27749 15258
rect 27773 15206 27787 15258
rect 27787 15206 27799 15258
rect 27799 15206 27829 15258
rect 27853 15206 27863 15258
rect 27863 15206 27909 15258
rect 27613 15204 27669 15206
rect 27693 15204 27749 15206
rect 27773 15204 27829 15206
rect 27853 15204 27909 15206
rect 27613 14170 27669 14172
rect 27693 14170 27749 14172
rect 27773 14170 27829 14172
rect 27853 14170 27909 14172
rect 27613 14118 27659 14170
rect 27659 14118 27669 14170
rect 27693 14118 27723 14170
rect 27723 14118 27735 14170
rect 27735 14118 27749 14170
rect 27773 14118 27787 14170
rect 27787 14118 27799 14170
rect 27799 14118 27829 14170
rect 27853 14118 27863 14170
rect 27863 14118 27909 14170
rect 27613 14116 27669 14118
rect 27693 14116 27749 14118
rect 27773 14116 27829 14118
rect 27853 14116 27909 14118
rect 27434 13388 27490 13424
rect 27434 13368 27436 13388
rect 27436 13368 27488 13388
rect 27488 13368 27490 13388
rect 27613 13082 27669 13084
rect 27693 13082 27749 13084
rect 27773 13082 27829 13084
rect 27853 13082 27909 13084
rect 27613 13030 27659 13082
rect 27659 13030 27669 13082
rect 27693 13030 27723 13082
rect 27723 13030 27735 13082
rect 27735 13030 27749 13082
rect 27773 13030 27787 13082
rect 27787 13030 27799 13082
rect 27799 13030 27829 13082
rect 27853 13030 27863 13082
rect 27863 13030 27909 13082
rect 27613 13028 27669 13030
rect 27693 13028 27749 13030
rect 27773 13028 27829 13030
rect 27853 13028 27909 13030
rect 27526 12844 27582 12880
rect 27526 12824 27528 12844
rect 27528 12824 27580 12844
rect 27580 12824 27582 12844
rect 28722 16632 28778 16688
rect 28906 19216 28962 19272
rect 28446 14320 28502 14376
rect 28630 13776 28686 13832
rect 29182 18808 29238 18864
rect 30286 20712 30342 20768
rect 29734 20440 29790 20496
rect 29734 15564 29790 15600
rect 29734 15544 29736 15564
rect 29736 15544 29788 15564
rect 29788 15544 29790 15564
rect 31500 21242 31556 21244
rect 31580 21242 31636 21244
rect 31660 21242 31716 21244
rect 31740 21242 31796 21244
rect 31500 21190 31546 21242
rect 31546 21190 31556 21242
rect 31580 21190 31610 21242
rect 31610 21190 31622 21242
rect 31622 21190 31636 21242
rect 31660 21190 31674 21242
rect 31674 21190 31686 21242
rect 31686 21190 31716 21242
rect 31740 21190 31750 21242
rect 31750 21190 31796 21242
rect 31500 21188 31556 21190
rect 31580 21188 31636 21190
rect 31660 21188 31716 21190
rect 31740 21188 31796 21190
rect 30194 17856 30250 17912
rect 30102 14456 30158 14512
rect 31500 20154 31556 20156
rect 31580 20154 31636 20156
rect 31660 20154 31716 20156
rect 31740 20154 31796 20156
rect 31500 20102 31546 20154
rect 31546 20102 31556 20154
rect 31580 20102 31610 20154
rect 31610 20102 31622 20154
rect 31622 20102 31636 20154
rect 31660 20102 31674 20154
rect 31674 20102 31686 20154
rect 31686 20102 31716 20154
rect 31740 20102 31750 20154
rect 31750 20102 31796 20154
rect 31500 20100 31556 20102
rect 31580 20100 31636 20102
rect 31660 20100 31716 20102
rect 31740 20100 31796 20102
rect 31500 19066 31556 19068
rect 31580 19066 31636 19068
rect 31660 19066 31716 19068
rect 31740 19066 31796 19068
rect 31500 19014 31546 19066
rect 31546 19014 31556 19066
rect 31580 19014 31610 19066
rect 31610 19014 31622 19066
rect 31622 19014 31636 19066
rect 31660 19014 31674 19066
rect 31674 19014 31686 19066
rect 31686 19014 31716 19066
rect 31740 19014 31750 19066
rect 31750 19014 31796 19066
rect 31500 19012 31556 19014
rect 31580 19012 31636 19014
rect 31660 19012 31716 19014
rect 31740 19012 31796 19014
rect 31500 17978 31556 17980
rect 31580 17978 31636 17980
rect 31660 17978 31716 17980
rect 31740 17978 31796 17980
rect 31500 17926 31546 17978
rect 31546 17926 31556 17978
rect 31580 17926 31610 17978
rect 31610 17926 31622 17978
rect 31622 17926 31636 17978
rect 31660 17926 31674 17978
rect 31674 17926 31686 17978
rect 31686 17926 31716 17978
rect 31740 17926 31750 17978
rect 31750 17926 31796 17978
rect 31500 17924 31556 17926
rect 31580 17924 31636 17926
rect 31660 17924 31716 17926
rect 31740 17924 31796 17926
rect 31500 16890 31556 16892
rect 31580 16890 31636 16892
rect 31660 16890 31716 16892
rect 31740 16890 31796 16892
rect 31500 16838 31546 16890
rect 31546 16838 31556 16890
rect 31580 16838 31610 16890
rect 31610 16838 31622 16890
rect 31622 16838 31636 16890
rect 31660 16838 31674 16890
rect 31674 16838 31686 16890
rect 31686 16838 31716 16890
rect 31740 16838 31750 16890
rect 31750 16838 31796 16890
rect 31500 16836 31556 16838
rect 31580 16836 31636 16838
rect 31660 16836 31716 16838
rect 31740 16836 31796 16838
rect 31500 15802 31556 15804
rect 31580 15802 31636 15804
rect 31660 15802 31716 15804
rect 31740 15802 31796 15804
rect 31500 15750 31546 15802
rect 31546 15750 31556 15802
rect 31580 15750 31610 15802
rect 31610 15750 31622 15802
rect 31622 15750 31636 15802
rect 31660 15750 31674 15802
rect 31674 15750 31686 15802
rect 31686 15750 31716 15802
rect 31740 15750 31750 15802
rect 31750 15750 31796 15802
rect 31500 15748 31556 15750
rect 31580 15748 31636 15750
rect 31660 15748 31716 15750
rect 31740 15748 31796 15750
rect 31500 14714 31556 14716
rect 31580 14714 31636 14716
rect 31660 14714 31716 14716
rect 31740 14714 31796 14716
rect 31500 14662 31546 14714
rect 31546 14662 31556 14714
rect 31580 14662 31610 14714
rect 31610 14662 31622 14714
rect 31622 14662 31636 14714
rect 31660 14662 31674 14714
rect 31674 14662 31686 14714
rect 31686 14662 31716 14714
rect 31740 14662 31750 14714
rect 31750 14662 31796 14714
rect 31500 14660 31556 14662
rect 31580 14660 31636 14662
rect 31660 14660 31716 14662
rect 31740 14660 31796 14662
rect 31500 13626 31556 13628
rect 31580 13626 31636 13628
rect 31660 13626 31716 13628
rect 31740 13626 31796 13628
rect 31500 13574 31546 13626
rect 31546 13574 31556 13626
rect 31580 13574 31610 13626
rect 31610 13574 31622 13626
rect 31622 13574 31636 13626
rect 31660 13574 31674 13626
rect 31674 13574 31686 13626
rect 31686 13574 31716 13626
rect 31740 13574 31750 13626
rect 31750 13574 31796 13626
rect 31500 13572 31556 13574
rect 31580 13572 31636 13574
rect 31660 13572 31716 13574
rect 31740 13572 31796 13574
rect 31500 12538 31556 12540
rect 31580 12538 31636 12540
rect 31660 12538 31716 12540
rect 31740 12538 31796 12540
rect 31500 12486 31546 12538
rect 31546 12486 31556 12538
rect 31580 12486 31610 12538
rect 31610 12486 31622 12538
rect 31622 12486 31636 12538
rect 31660 12486 31674 12538
rect 31674 12486 31686 12538
rect 31686 12486 31716 12538
rect 31740 12486 31750 12538
rect 31750 12486 31796 12538
rect 31500 12484 31556 12486
rect 31580 12484 31636 12486
rect 31660 12484 31716 12486
rect 31740 12484 31796 12486
rect 27613 11994 27669 11996
rect 27693 11994 27749 11996
rect 27773 11994 27829 11996
rect 27853 11994 27909 11996
rect 27613 11942 27659 11994
rect 27659 11942 27669 11994
rect 27693 11942 27723 11994
rect 27723 11942 27735 11994
rect 27735 11942 27749 11994
rect 27773 11942 27787 11994
rect 27787 11942 27799 11994
rect 27799 11942 27829 11994
rect 27853 11942 27863 11994
rect 27863 11942 27909 11994
rect 27613 11940 27669 11942
rect 27693 11940 27749 11942
rect 27773 11940 27829 11942
rect 27853 11940 27909 11942
rect 27613 10906 27669 10908
rect 27693 10906 27749 10908
rect 27773 10906 27829 10908
rect 27853 10906 27909 10908
rect 27613 10854 27659 10906
rect 27659 10854 27669 10906
rect 27693 10854 27723 10906
rect 27723 10854 27735 10906
rect 27735 10854 27749 10906
rect 27773 10854 27787 10906
rect 27787 10854 27799 10906
rect 27799 10854 27829 10906
rect 27853 10854 27863 10906
rect 27863 10854 27909 10906
rect 27613 10852 27669 10854
rect 27693 10852 27749 10854
rect 27773 10852 27829 10854
rect 27853 10852 27909 10854
rect 27618 10104 27674 10160
rect 27613 9818 27669 9820
rect 27693 9818 27749 9820
rect 27773 9818 27829 9820
rect 27853 9818 27909 9820
rect 27613 9766 27659 9818
rect 27659 9766 27669 9818
rect 27693 9766 27723 9818
rect 27723 9766 27735 9818
rect 27735 9766 27749 9818
rect 27773 9766 27787 9818
rect 27787 9766 27799 9818
rect 27799 9766 27829 9818
rect 27853 9766 27863 9818
rect 27863 9766 27909 9818
rect 27613 9764 27669 9766
rect 27693 9764 27749 9766
rect 27773 9764 27829 9766
rect 27853 9764 27909 9766
rect 27802 9560 27858 9616
rect 29734 12144 29790 12200
rect 29918 11736 29974 11792
rect 31500 11450 31556 11452
rect 31580 11450 31636 11452
rect 31660 11450 31716 11452
rect 31740 11450 31796 11452
rect 31500 11398 31546 11450
rect 31546 11398 31556 11450
rect 31580 11398 31610 11450
rect 31610 11398 31622 11450
rect 31622 11398 31636 11450
rect 31660 11398 31674 11450
rect 31674 11398 31686 11450
rect 31686 11398 31716 11450
rect 31740 11398 31750 11450
rect 31750 11398 31796 11450
rect 31500 11396 31556 11398
rect 31580 11396 31636 11398
rect 31660 11396 31716 11398
rect 31740 11396 31796 11398
rect 31500 10362 31556 10364
rect 31580 10362 31636 10364
rect 31660 10362 31716 10364
rect 31740 10362 31796 10364
rect 31500 10310 31546 10362
rect 31546 10310 31556 10362
rect 31580 10310 31610 10362
rect 31610 10310 31622 10362
rect 31622 10310 31636 10362
rect 31660 10310 31674 10362
rect 31674 10310 31686 10362
rect 31686 10310 31716 10362
rect 31740 10310 31750 10362
rect 31750 10310 31796 10362
rect 31500 10308 31556 10310
rect 31580 10308 31636 10310
rect 31660 10308 31716 10310
rect 31740 10308 31796 10310
rect 31500 9274 31556 9276
rect 31580 9274 31636 9276
rect 31660 9274 31716 9276
rect 31740 9274 31796 9276
rect 31500 9222 31546 9274
rect 31546 9222 31556 9274
rect 31580 9222 31610 9274
rect 31610 9222 31622 9274
rect 31622 9222 31636 9274
rect 31660 9222 31674 9274
rect 31674 9222 31686 9274
rect 31686 9222 31716 9274
rect 31740 9222 31750 9274
rect 31750 9222 31796 9274
rect 31500 9220 31556 9222
rect 31580 9220 31636 9222
rect 31660 9220 31716 9222
rect 31740 9220 31796 9222
rect 27613 8730 27669 8732
rect 27693 8730 27749 8732
rect 27773 8730 27829 8732
rect 27853 8730 27909 8732
rect 27613 8678 27659 8730
rect 27659 8678 27669 8730
rect 27693 8678 27723 8730
rect 27723 8678 27735 8730
rect 27735 8678 27749 8730
rect 27773 8678 27787 8730
rect 27787 8678 27799 8730
rect 27799 8678 27829 8730
rect 27853 8678 27863 8730
rect 27863 8678 27909 8730
rect 27613 8676 27669 8678
rect 27693 8676 27749 8678
rect 27773 8676 27829 8678
rect 27853 8676 27909 8678
rect 25686 6024 25742 6080
rect 25502 5516 25504 5536
rect 25504 5516 25556 5536
rect 25556 5516 25558 5536
rect 25502 5480 25558 5516
rect 25778 4664 25834 4720
rect 25226 3440 25282 3496
rect 25594 4004 25650 4040
rect 25594 3984 25596 4004
rect 25596 3984 25648 4004
rect 25648 3984 25650 4004
rect 26238 5908 26294 5944
rect 26238 5888 26240 5908
rect 26240 5888 26292 5908
rect 26292 5888 26294 5908
rect 25962 5092 26018 5128
rect 25962 5072 25964 5092
rect 25964 5072 26016 5092
rect 26016 5072 26018 5092
rect 26698 6432 26754 6488
rect 26422 5752 26478 5808
rect 26514 5652 26516 5672
rect 26516 5652 26568 5672
rect 26568 5652 26570 5672
rect 26514 5616 26570 5652
rect 27066 5480 27122 5536
rect 26882 4700 26884 4720
rect 26884 4700 26936 4720
rect 26936 4700 26938 4720
rect 26882 4664 26938 4700
rect 26882 4528 26938 4584
rect 27158 5208 27214 5264
rect 27158 4020 27160 4040
rect 27160 4020 27212 4040
rect 27212 4020 27214 4040
rect 27158 3984 27214 4020
rect 27613 7642 27669 7644
rect 27693 7642 27749 7644
rect 27773 7642 27829 7644
rect 27853 7642 27909 7644
rect 27613 7590 27659 7642
rect 27659 7590 27669 7642
rect 27693 7590 27723 7642
rect 27723 7590 27735 7642
rect 27735 7590 27749 7642
rect 27773 7590 27787 7642
rect 27787 7590 27799 7642
rect 27799 7590 27829 7642
rect 27853 7590 27863 7642
rect 27863 7590 27909 7642
rect 27613 7588 27669 7590
rect 27693 7588 27749 7590
rect 27773 7588 27829 7590
rect 27853 7588 27909 7590
rect 27613 6554 27669 6556
rect 27693 6554 27749 6556
rect 27773 6554 27829 6556
rect 27853 6554 27909 6556
rect 27613 6502 27659 6554
rect 27659 6502 27669 6554
rect 27693 6502 27723 6554
rect 27723 6502 27735 6554
rect 27735 6502 27749 6554
rect 27773 6502 27787 6554
rect 27787 6502 27799 6554
rect 27799 6502 27829 6554
rect 27853 6502 27863 6554
rect 27863 6502 27909 6554
rect 27613 6500 27669 6502
rect 27693 6500 27749 6502
rect 27773 6500 27829 6502
rect 27853 6500 27909 6502
rect 31500 8186 31556 8188
rect 31580 8186 31636 8188
rect 31660 8186 31716 8188
rect 31740 8186 31796 8188
rect 31500 8134 31546 8186
rect 31546 8134 31556 8186
rect 31580 8134 31610 8186
rect 31610 8134 31622 8186
rect 31622 8134 31636 8186
rect 31660 8134 31674 8186
rect 31674 8134 31686 8186
rect 31686 8134 31716 8186
rect 31740 8134 31750 8186
rect 31750 8134 31796 8186
rect 31500 8132 31556 8134
rect 31580 8132 31636 8134
rect 31660 8132 31716 8134
rect 31740 8132 31796 8134
rect 28354 7812 28410 7848
rect 28354 7792 28356 7812
rect 28356 7792 28408 7812
rect 28408 7792 28410 7812
rect 27618 6180 27674 6216
rect 27618 6160 27620 6180
rect 27620 6160 27672 6180
rect 27672 6160 27674 6180
rect 27613 5466 27669 5468
rect 27693 5466 27749 5468
rect 27773 5466 27829 5468
rect 27853 5466 27909 5468
rect 27613 5414 27659 5466
rect 27659 5414 27669 5466
rect 27693 5414 27723 5466
rect 27723 5414 27735 5466
rect 27735 5414 27749 5466
rect 27773 5414 27787 5466
rect 27787 5414 27799 5466
rect 27799 5414 27829 5466
rect 27853 5414 27863 5466
rect 27863 5414 27909 5466
rect 27613 5412 27669 5414
rect 27693 5412 27749 5414
rect 27773 5412 27829 5414
rect 27853 5412 27909 5414
rect 27618 4528 27674 4584
rect 27613 4378 27669 4380
rect 27693 4378 27749 4380
rect 27773 4378 27829 4380
rect 27853 4378 27909 4380
rect 27613 4326 27659 4378
rect 27659 4326 27669 4378
rect 27693 4326 27723 4378
rect 27723 4326 27735 4378
rect 27735 4326 27749 4378
rect 27773 4326 27787 4378
rect 27787 4326 27799 4378
rect 27799 4326 27829 4378
rect 27853 4326 27863 4378
rect 27863 4326 27909 4378
rect 27613 4324 27669 4326
rect 27693 4324 27749 4326
rect 27773 4324 27829 4326
rect 27853 4324 27909 4326
rect 31500 7098 31556 7100
rect 31580 7098 31636 7100
rect 31660 7098 31716 7100
rect 31740 7098 31796 7100
rect 31500 7046 31546 7098
rect 31546 7046 31556 7098
rect 31580 7046 31610 7098
rect 31610 7046 31622 7098
rect 31622 7046 31636 7098
rect 31660 7046 31674 7098
rect 31674 7046 31686 7098
rect 31686 7046 31716 7098
rect 31740 7046 31750 7098
rect 31750 7046 31796 7098
rect 31500 7044 31556 7046
rect 31580 7044 31636 7046
rect 31660 7044 31716 7046
rect 31740 7044 31796 7046
rect 31500 6010 31556 6012
rect 31580 6010 31636 6012
rect 31660 6010 31716 6012
rect 31740 6010 31796 6012
rect 31500 5958 31546 6010
rect 31546 5958 31556 6010
rect 31580 5958 31610 6010
rect 31610 5958 31622 6010
rect 31622 5958 31636 6010
rect 31660 5958 31674 6010
rect 31674 5958 31686 6010
rect 31686 5958 31716 6010
rect 31740 5958 31750 6010
rect 31750 5958 31796 6010
rect 31500 5956 31556 5958
rect 31580 5956 31636 5958
rect 31660 5956 31716 5958
rect 31740 5956 31796 5958
rect 27613 3290 27669 3292
rect 27693 3290 27749 3292
rect 27773 3290 27829 3292
rect 27853 3290 27909 3292
rect 27613 3238 27659 3290
rect 27659 3238 27669 3290
rect 27693 3238 27723 3290
rect 27723 3238 27735 3290
rect 27735 3238 27749 3290
rect 27773 3238 27787 3290
rect 27787 3238 27799 3290
rect 27799 3238 27829 3290
rect 27853 3238 27863 3290
rect 27863 3238 27909 3290
rect 27613 3236 27669 3238
rect 27693 3236 27749 3238
rect 27773 3236 27829 3238
rect 27853 3236 27909 3238
rect 23726 1658 23782 1660
rect 23806 1658 23862 1660
rect 23886 1658 23942 1660
rect 23966 1658 24022 1660
rect 23726 1606 23772 1658
rect 23772 1606 23782 1658
rect 23806 1606 23836 1658
rect 23836 1606 23848 1658
rect 23848 1606 23862 1658
rect 23886 1606 23900 1658
rect 23900 1606 23912 1658
rect 23912 1606 23942 1658
rect 23966 1606 23976 1658
rect 23976 1606 24022 1658
rect 23726 1604 23782 1606
rect 23806 1604 23862 1606
rect 23886 1604 23942 1606
rect 23966 1604 24022 1606
rect 27613 2202 27669 2204
rect 27693 2202 27749 2204
rect 27773 2202 27829 2204
rect 27853 2202 27909 2204
rect 27613 2150 27659 2202
rect 27659 2150 27669 2202
rect 27693 2150 27723 2202
rect 27723 2150 27735 2202
rect 27735 2150 27749 2202
rect 27773 2150 27787 2202
rect 27787 2150 27799 2202
rect 27799 2150 27829 2202
rect 27853 2150 27863 2202
rect 27863 2150 27909 2202
rect 27613 2148 27669 2150
rect 27693 2148 27749 2150
rect 27773 2148 27829 2150
rect 27853 2148 27909 2150
rect 28262 3712 28318 3768
rect 31500 4922 31556 4924
rect 31580 4922 31636 4924
rect 31660 4922 31716 4924
rect 31740 4922 31796 4924
rect 31500 4870 31546 4922
rect 31546 4870 31556 4922
rect 31580 4870 31610 4922
rect 31610 4870 31622 4922
rect 31622 4870 31636 4922
rect 31660 4870 31674 4922
rect 31674 4870 31686 4922
rect 31686 4870 31716 4922
rect 31740 4870 31750 4922
rect 31750 4870 31796 4922
rect 31500 4868 31556 4870
rect 31580 4868 31636 4870
rect 31660 4868 31716 4870
rect 31740 4868 31796 4870
rect 31500 3834 31556 3836
rect 31580 3834 31636 3836
rect 31660 3834 31716 3836
rect 31740 3834 31796 3836
rect 31500 3782 31546 3834
rect 31546 3782 31556 3834
rect 31580 3782 31610 3834
rect 31610 3782 31622 3834
rect 31622 3782 31636 3834
rect 31660 3782 31674 3834
rect 31674 3782 31686 3834
rect 31686 3782 31716 3834
rect 31740 3782 31750 3834
rect 31750 3782 31796 3834
rect 31500 3780 31556 3782
rect 31580 3780 31636 3782
rect 31660 3780 31716 3782
rect 31740 3780 31796 3782
rect 28630 3032 28686 3088
rect 31500 2746 31556 2748
rect 31580 2746 31636 2748
rect 31660 2746 31716 2748
rect 31740 2746 31796 2748
rect 31500 2694 31546 2746
rect 31546 2694 31556 2746
rect 31580 2694 31610 2746
rect 31610 2694 31622 2746
rect 31622 2694 31636 2746
rect 31660 2694 31674 2746
rect 31674 2694 31686 2746
rect 31686 2694 31716 2746
rect 31740 2694 31750 2746
rect 31750 2694 31796 2746
rect 31500 2692 31556 2694
rect 31580 2692 31636 2694
rect 31660 2692 31716 2694
rect 31740 2692 31796 2694
rect 31500 1658 31556 1660
rect 31580 1658 31636 1660
rect 31660 1658 31716 1660
rect 31740 1658 31796 1660
rect 31500 1606 31546 1658
rect 31546 1606 31556 1658
rect 31580 1606 31610 1658
rect 31610 1606 31622 1658
rect 31622 1606 31636 1658
rect 31660 1606 31674 1658
rect 31674 1606 31686 1658
rect 31686 1606 31716 1658
rect 31740 1606 31750 1658
rect 31750 1606 31796 1658
rect 31500 1604 31556 1606
rect 31580 1604 31636 1606
rect 31660 1604 31716 1606
rect 31740 1604 31796 1606
rect 4291 1114 4347 1116
rect 4371 1114 4427 1116
rect 4451 1114 4507 1116
rect 4531 1114 4587 1116
rect 4291 1062 4337 1114
rect 4337 1062 4347 1114
rect 4371 1062 4401 1114
rect 4401 1062 4413 1114
rect 4413 1062 4427 1114
rect 4451 1062 4465 1114
rect 4465 1062 4477 1114
rect 4477 1062 4507 1114
rect 4531 1062 4541 1114
rect 4541 1062 4587 1114
rect 4291 1060 4347 1062
rect 4371 1060 4427 1062
rect 4451 1060 4507 1062
rect 4531 1060 4587 1062
rect 12065 1114 12121 1116
rect 12145 1114 12201 1116
rect 12225 1114 12281 1116
rect 12305 1114 12361 1116
rect 12065 1062 12111 1114
rect 12111 1062 12121 1114
rect 12145 1062 12175 1114
rect 12175 1062 12187 1114
rect 12187 1062 12201 1114
rect 12225 1062 12239 1114
rect 12239 1062 12251 1114
rect 12251 1062 12281 1114
rect 12305 1062 12315 1114
rect 12315 1062 12361 1114
rect 12065 1060 12121 1062
rect 12145 1060 12201 1062
rect 12225 1060 12281 1062
rect 12305 1060 12361 1062
rect 19839 1114 19895 1116
rect 19919 1114 19975 1116
rect 19999 1114 20055 1116
rect 20079 1114 20135 1116
rect 19839 1062 19885 1114
rect 19885 1062 19895 1114
rect 19919 1062 19949 1114
rect 19949 1062 19961 1114
rect 19961 1062 19975 1114
rect 19999 1062 20013 1114
rect 20013 1062 20025 1114
rect 20025 1062 20055 1114
rect 20079 1062 20089 1114
rect 20089 1062 20135 1114
rect 19839 1060 19895 1062
rect 19919 1060 19975 1062
rect 19999 1060 20055 1062
rect 20079 1060 20135 1062
rect 27613 1114 27669 1116
rect 27693 1114 27749 1116
rect 27773 1114 27829 1116
rect 27853 1114 27909 1116
rect 27613 1062 27659 1114
rect 27659 1062 27669 1114
rect 27693 1062 27723 1114
rect 27723 1062 27735 1114
rect 27735 1062 27749 1114
rect 27773 1062 27787 1114
rect 27787 1062 27799 1114
rect 27799 1062 27829 1114
rect 27853 1062 27863 1114
rect 27863 1062 27909 1114
rect 27613 1060 27669 1062
rect 27693 1060 27749 1062
rect 27773 1060 27829 1062
rect 27853 1060 27909 1062
rect 8178 570 8234 572
rect 8258 570 8314 572
rect 8338 570 8394 572
rect 8418 570 8474 572
rect 8178 518 8224 570
rect 8224 518 8234 570
rect 8258 518 8288 570
rect 8288 518 8300 570
rect 8300 518 8314 570
rect 8338 518 8352 570
rect 8352 518 8364 570
rect 8364 518 8394 570
rect 8418 518 8428 570
rect 8428 518 8474 570
rect 8178 516 8234 518
rect 8258 516 8314 518
rect 8338 516 8394 518
rect 8418 516 8474 518
rect 15952 570 16008 572
rect 16032 570 16088 572
rect 16112 570 16168 572
rect 16192 570 16248 572
rect 15952 518 15998 570
rect 15998 518 16008 570
rect 16032 518 16062 570
rect 16062 518 16074 570
rect 16074 518 16088 570
rect 16112 518 16126 570
rect 16126 518 16138 570
rect 16138 518 16168 570
rect 16192 518 16202 570
rect 16202 518 16248 570
rect 15952 516 16008 518
rect 16032 516 16088 518
rect 16112 516 16168 518
rect 16192 516 16248 518
rect 23726 570 23782 572
rect 23806 570 23862 572
rect 23886 570 23942 572
rect 23966 570 24022 572
rect 23726 518 23772 570
rect 23772 518 23782 570
rect 23806 518 23836 570
rect 23836 518 23848 570
rect 23848 518 23862 570
rect 23886 518 23900 570
rect 23900 518 23912 570
rect 23912 518 23942 570
rect 23966 518 23976 570
rect 23976 518 24022 570
rect 23726 516 23782 518
rect 23806 516 23862 518
rect 23886 516 23942 518
rect 23966 516 24022 518
rect 31500 570 31556 572
rect 31580 570 31636 572
rect 31660 570 31716 572
rect 31740 570 31796 572
rect 31500 518 31546 570
rect 31546 518 31556 570
rect 31580 518 31610 570
rect 31610 518 31622 570
rect 31622 518 31636 570
rect 31660 518 31674 570
rect 31674 518 31686 570
rect 31686 518 31716 570
rect 31740 518 31750 570
rect 31750 518 31796 570
rect 31500 516 31556 518
rect 31580 516 31636 518
rect 31660 516 31716 518
rect 31740 516 31796 518
<< metal3 >>
rect 13721 22130 13787 22133
rect 14774 22130 14780 22132
rect 13721 22128 14780 22130
rect 13721 22072 13726 22128
rect 13782 22072 14780 22128
rect 13721 22070 14780 22072
rect 13721 22067 13787 22070
rect 14774 22068 14780 22070
rect 14844 22068 14850 22132
rect 4521 21996 4587 21997
rect 4470 21932 4476 21996
rect 4540 21994 4587 21996
rect 4540 21992 4632 21994
rect 4582 21936 4632 21992
rect 4540 21934 4632 21936
rect 4540 21932 4587 21934
rect 9622 21932 9628 21996
rect 9692 21994 9698 21996
rect 12525 21994 12591 21997
rect 9692 21992 12591 21994
rect 9692 21936 12530 21992
rect 12586 21936 12591 21992
rect 9692 21934 12591 21936
rect 9692 21932 9698 21934
rect 4521 21931 4587 21932
rect 12525 21931 12591 21934
rect 13721 21994 13787 21997
rect 16246 21994 16252 21996
rect 13721 21992 16252 21994
rect 13721 21936 13726 21992
rect 13782 21936 16252 21992
rect 13721 21934 16252 21936
rect 13721 21931 13787 21934
rect 16246 21932 16252 21934
rect 16316 21932 16322 21996
rect 25078 21932 25084 21996
rect 25148 21994 25154 21996
rect 26049 21994 26115 21997
rect 25148 21992 26115 21994
rect 25148 21936 26054 21992
rect 26110 21936 26115 21992
rect 25148 21934 26115 21936
rect 25148 21932 25154 21934
rect 26049 21931 26115 21934
rect 28758 21932 28764 21996
rect 28828 21994 28834 21996
rect 29729 21994 29795 21997
rect 28828 21992 29795 21994
rect 28828 21936 29734 21992
rect 29790 21936 29795 21992
rect 28828 21934 29795 21936
rect 28828 21932 28834 21934
rect 29729 21931 29795 21934
rect 6678 21796 6684 21860
rect 6748 21858 6754 21860
rect 7005 21858 7071 21861
rect 6748 21856 7071 21858
rect 6748 21800 7010 21856
rect 7066 21800 7071 21856
rect 6748 21798 7071 21800
rect 6748 21796 6754 21798
rect 7005 21795 7071 21798
rect 7414 21796 7420 21860
rect 7484 21858 7490 21860
rect 8845 21858 8911 21861
rect 7484 21856 8911 21858
rect 7484 21800 8850 21856
rect 8906 21800 8911 21856
rect 7484 21798 8911 21800
rect 7484 21796 7490 21798
rect 8845 21795 8911 21798
rect 12566 21796 12572 21860
rect 12636 21858 12642 21860
rect 13813 21858 13879 21861
rect 12636 21856 13879 21858
rect 12636 21800 13818 21856
rect 13874 21800 13879 21856
rect 12636 21798 13879 21800
rect 12636 21796 12642 21798
rect 13813 21795 13879 21798
rect 24342 21796 24348 21860
rect 24412 21858 24418 21860
rect 24669 21858 24735 21861
rect 24412 21856 24735 21858
rect 24412 21800 24674 21856
rect 24730 21800 24735 21856
rect 24412 21798 24735 21800
rect 24412 21796 24418 21798
rect 24669 21795 24735 21798
rect 25814 21796 25820 21860
rect 25884 21858 25890 21860
rect 26601 21858 26667 21861
rect 28073 21860 28139 21861
rect 25884 21856 26667 21858
rect 25884 21800 26606 21856
rect 26662 21800 26667 21856
rect 25884 21798 26667 21800
rect 25884 21796 25890 21798
rect 26601 21795 26667 21798
rect 28022 21796 28028 21860
rect 28092 21858 28139 21860
rect 28092 21856 28184 21858
rect 28134 21800 28184 21856
rect 28092 21798 28184 21800
rect 28092 21796 28139 21798
rect 29494 21796 29500 21860
rect 29564 21858 29570 21860
rect 30005 21858 30071 21861
rect 30281 21860 30347 21861
rect 30230 21858 30236 21860
rect 29564 21856 30071 21858
rect 29564 21800 30010 21856
rect 30066 21800 30071 21856
rect 29564 21798 30071 21800
rect 30190 21798 30236 21858
rect 30300 21856 30347 21860
rect 30342 21800 30347 21856
rect 29564 21796 29570 21798
rect 28073 21795 28139 21796
rect 30005 21795 30071 21798
rect 30230 21796 30236 21798
rect 30300 21796 30347 21800
rect 30281 21795 30347 21796
rect 4281 21792 4597 21793
rect 4281 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4597 21792
rect 4281 21727 4597 21728
rect 12055 21792 12371 21793
rect 12055 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12371 21792
rect 12055 21727 12371 21728
rect 19829 21792 20145 21793
rect 19829 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20145 21792
rect 19829 21727 20145 21728
rect 27603 21792 27919 21793
rect 27603 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27919 21792
rect 27603 21727 27919 21728
rect 13353 21724 13419 21725
rect 13302 21722 13308 21724
rect 13262 21662 13308 21722
rect 13372 21720 13419 21724
rect 13414 21664 13419 21720
rect 13302 21660 13308 21662
rect 13372 21660 13419 21664
rect 26550 21660 26556 21724
rect 26620 21722 26626 21724
rect 27429 21722 27495 21725
rect 26620 21720 27495 21722
rect 26620 21664 27434 21720
rect 27490 21664 27495 21720
rect 26620 21662 27495 21664
rect 26620 21660 26626 21662
rect 13353 21659 13419 21660
rect 27429 21659 27495 21662
rect 3734 21524 3740 21588
rect 3804 21586 3810 21588
rect 4981 21586 5047 21589
rect 3804 21584 5047 21586
rect 3804 21528 4986 21584
rect 5042 21528 5047 21584
rect 3804 21526 5047 21528
rect 3804 21524 3810 21526
rect 4981 21523 5047 21526
rect 13537 21586 13603 21589
rect 14038 21586 14044 21588
rect 13537 21584 14044 21586
rect 13537 21528 13542 21584
rect 13598 21528 14044 21584
rect 13537 21526 14044 21528
rect 13537 21523 13603 21526
rect 14038 21524 14044 21526
rect 14108 21524 14114 21588
rect 14733 21586 14799 21589
rect 17718 21586 17724 21588
rect 14733 21584 17724 21586
rect 14733 21528 14738 21584
rect 14794 21528 17724 21584
rect 14733 21526 17724 21528
rect 14733 21523 14799 21526
rect 17718 21524 17724 21526
rect 17788 21524 17794 21588
rect 27286 21524 27292 21588
rect 27356 21586 27362 21588
rect 27705 21586 27771 21589
rect 27356 21584 27771 21586
rect 27356 21528 27710 21584
rect 27766 21528 27771 21584
rect 27356 21526 27771 21528
rect 27356 21524 27362 21526
rect 27705 21523 27771 21526
rect 15101 21450 15167 21453
rect 15510 21450 15516 21452
rect 15101 21448 15516 21450
rect 15101 21392 15106 21448
rect 15162 21392 15516 21448
rect 15101 21390 15516 21392
rect 15101 21387 15167 21390
rect 15510 21388 15516 21390
rect 15580 21388 15586 21452
rect 15745 21450 15811 21453
rect 19149 21450 19215 21453
rect 15745 21448 19215 21450
rect 15745 21392 15750 21448
rect 15806 21392 19154 21448
rect 19210 21392 19215 21448
rect 15745 21390 19215 21392
rect 15745 21387 15811 21390
rect 19149 21387 19215 21390
rect 790 21252 796 21316
rect 860 21314 866 21316
rect 1301 21314 1367 21317
rect 6177 21314 6243 21317
rect 860 21312 6243 21314
rect 860 21256 1306 21312
rect 1362 21256 6182 21312
rect 6238 21256 6243 21312
rect 860 21254 6243 21256
rect 860 21252 866 21254
rect 1301 21251 1367 21254
rect 6177 21251 6243 21254
rect 13261 21314 13327 21317
rect 14181 21314 14247 21317
rect 13261 21312 14247 21314
rect 13261 21256 13266 21312
rect 13322 21256 14186 21312
rect 14242 21256 14247 21312
rect 13261 21254 14247 21256
rect 13261 21251 13327 21254
rect 14181 21251 14247 21254
rect 18505 21314 18571 21317
rect 23381 21314 23447 21317
rect 18505 21312 23447 21314
rect 18505 21256 18510 21312
rect 18566 21256 23386 21312
rect 23442 21256 23447 21312
rect 18505 21254 23447 21256
rect 18505 21251 18571 21254
rect 23381 21251 23447 21254
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 15942 21248 16258 21249
rect 15942 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16258 21248
rect 15942 21183 16258 21184
rect 23716 21248 24032 21249
rect 23716 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24032 21248
rect 23716 21183 24032 21184
rect 31490 21248 31806 21249
rect 31490 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31806 21248
rect 31490 21183 31806 21184
rect 1526 21116 1532 21180
rect 1596 21178 1602 21180
rect 2129 21178 2195 21181
rect 1596 21176 2195 21178
rect 1596 21120 2134 21176
rect 2190 21120 2195 21176
rect 1596 21118 2195 21120
rect 1596 21116 1602 21118
rect 2129 21115 2195 21118
rect 2998 21116 3004 21180
rect 3068 21178 3074 21180
rect 3969 21178 4035 21181
rect 3068 21176 4035 21178
rect 3068 21120 3974 21176
rect 4030 21120 4035 21176
rect 3068 21118 4035 21120
rect 3068 21116 3074 21118
rect 3969 21115 4035 21118
rect 5942 21116 5948 21180
rect 6012 21178 6018 21180
rect 6453 21178 6519 21181
rect 6012 21176 6519 21178
rect 6012 21120 6458 21176
rect 6514 21120 6519 21176
rect 6012 21118 6519 21120
rect 6012 21116 6018 21118
rect 6453 21115 6519 21118
rect 10409 21044 10475 21045
rect 10358 21042 10364 21044
rect 10318 20982 10364 21042
rect 10428 21040 10475 21044
rect 10470 20984 10475 21040
rect 10358 20980 10364 20982
rect 10428 20980 10475 20984
rect 10409 20979 10475 20980
rect 12341 21042 12407 21045
rect 12750 21042 12756 21044
rect 12341 21040 12756 21042
rect 12341 20984 12346 21040
rect 12402 20984 12756 21040
rect 12341 20982 12756 20984
rect 12341 20979 12407 20982
rect 12750 20980 12756 20982
rect 12820 20980 12826 21044
rect 19241 21042 19307 21045
rect 19374 21042 19380 21044
rect 19241 21040 19380 21042
rect 19241 20984 19246 21040
rect 19302 20984 19380 21040
rect 19241 20982 19380 20984
rect 19241 20979 19307 20982
rect 19374 20980 19380 20982
rect 19444 20980 19450 21044
rect 22829 21042 22895 21045
rect 25405 21042 25471 21045
rect 22829 21040 25471 21042
rect 22829 20984 22834 21040
rect 22890 20984 25410 21040
rect 25466 20984 25471 21040
rect 22829 20982 25471 20984
rect 22829 20979 22895 20982
rect 25405 20979 25471 20982
rect 11421 20906 11487 20909
rect 15101 20906 15167 20909
rect 11421 20904 15167 20906
rect 11421 20848 11426 20904
rect 11482 20848 15106 20904
rect 15162 20848 15167 20904
rect 11421 20846 15167 20848
rect 11421 20843 11487 20846
rect 15101 20843 15167 20846
rect 16481 20906 16547 20909
rect 20713 20906 20779 20909
rect 16481 20904 20779 20906
rect 16481 20848 16486 20904
rect 16542 20848 20718 20904
rect 20774 20848 20779 20904
rect 16481 20846 20779 20848
rect 16481 20843 16547 20846
rect 20713 20843 20779 20846
rect 1577 20770 1643 20773
rect 2262 20770 2268 20772
rect 1577 20768 2268 20770
rect 1577 20712 1582 20768
rect 1638 20712 2268 20768
rect 1577 20710 2268 20712
rect 1577 20707 1643 20710
rect 2262 20708 2268 20710
rect 2332 20770 2338 20772
rect 3325 20770 3391 20773
rect 6361 20772 6427 20773
rect 2332 20768 3391 20770
rect 2332 20712 3330 20768
rect 3386 20712 3391 20768
rect 2332 20710 3391 20712
rect 2332 20708 2338 20710
rect 3325 20707 3391 20710
rect 6310 20708 6316 20772
rect 6380 20770 6427 20772
rect 10317 20770 10383 20773
rect 10910 20770 10916 20772
rect 6380 20768 6472 20770
rect 6422 20712 6472 20768
rect 6380 20710 6472 20712
rect 10317 20768 10916 20770
rect 10317 20712 10322 20768
rect 10378 20712 10916 20768
rect 10317 20710 10916 20712
rect 6380 20708 6427 20710
rect 6361 20707 6427 20708
rect 10317 20707 10383 20710
rect 10910 20708 10916 20710
rect 10980 20708 10986 20772
rect 18413 20770 18479 20773
rect 19517 20770 19583 20773
rect 18413 20768 19583 20770
rect 18413 20712 18418 20768
rect 18474 20712 19522 20768
rect 19578 20712 19583 20768
rect 18413 20710 19583 20712
rect 18413 20707 18479 20710
rect 19517 20707 19583 20710
rect 21541 20770 21607 20773
rect 24669 20770 24735 20773
rect 21541 20768 24735 20770
rect 21541 20712 21546 20768
rect 21602 20712 24674 20768
rect 24730 20712 24735 20768
rect 21541 20710 24735 20712
rect 21541 20707 21607 20710
rect 24669 20707 24735 20710
rect 30046 20708 30052 20772
rect 30116 20770 30122 20772
rect 30281 20770 30347 20773
rect 30116 20768 30347 20770
rect 30116 20712 30286 20768
rect 30342 20712 30347 20768
rect 30116 20710 30347 20712
rect 30116 20708 30122 20710
rect 30281 20707 30347 20710
rect 4281 20704 4597 20705
rect 4281 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4597 20704
rect 4281 20639 4597 20640
rect 12055 20704 12371 20705
rect 12055 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12371 20704
rect 12055 20639 12371 20640
rect 19829 20704 20145 20705
rect 19829 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20145 20704
rect 19829 20639 20145 20640
rect 27603 20704 27919 20705
rect 27603 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27919 20704
rect 27603 20639 27919 20640
rect 7925 20636 7991 20637
rect 7925 20632 7972 20636
rect 8036 20634 8042 20636
rect 8661 20634 8727 20637
rect 11789 20636 11855 20637
rect 9622 20634 9628 20636
rect 7925 20576 7930 20632
rect 7925 20572 7972 20576
rect 8036 20574 8082 20634
rect 8661 20632 9628 20634
rect 8661 20576 8666 20632
rect 8722 20576 9628 20632
rect 8661 20574 9628 20576
rect 8036 20572 8042 20574
rect 7925 20571 7991 20572
rect 8661 20571 8727 20574
rect 9622 20572 9628 20574
rect 9692 20572 9698 20636
rect 11789 20632 11836 20636
rect 11900 20634 11906 20636
rect 13721 20634 13787 20637
rect 16982 20634 16988 20636
rect 11789 20576 11794 20632
rect 11789 20572 11836 20576
rect 11900 20574 11946 20634
rect 13678 20632 16988 20634
rect 13678 20576 13726 20632
rect 13782 20576 16988 20632
rect 13678 20574 16988 20576
rect 11900 20572 11906 20574
rect 11789 20571 11855 20572
rect 13678 20571 13787 20574
rect 16982 20572 16988 20574
rect 17052 20572 17058 20636
rect 7833 20498 7899 20501
rect 13678 20498 13738 20571
rect 7833 20496 13738 20498
rect 7833 20440 7838 20496
rect 7894 20440 13738 20496
rect 7833 20438 13738 20440
rect 15929 20498 15995 20501
rect 23289 20498 23355 20501
rect 15929 20496 23355 20498
rect 15929 20440 15934 20496
rect 15990 20440 23294 20496
rect 23350 20440 23355 20496
rect 15929 20438 23355 20440
rect 7833 20435 7899 20438
rect 15929 20435 15995 20438
rect 23289 20435 23355 20438
rect 23749 20498 23815 20501
rect 29729 20498 29795 20501
rect 23749 20496 29795 20498
rect 23749 20440 23754 20496
rect 23810 20440 29734 20496
rect 29790 20440 29795 20496
rect 23749 20438 29795 20440
rect 23749 20435 23815 20438
rect 29729 20435 29795 20438
rect 16941 20362 17007 20365
rect 17718 20362 17724 20364
rect 16941 20360 17724 20362
rect 16941 20304 16946 20360
rect 17002 20304 17724 20360
rect 16941 20302 17724 20304
rect 16941 20299 17007 20302
rect 17718 20300 17724 20302
rect 17788 20362 17794 20364
rect 23105 20362 23171 20365
rect 17788 20360 23171 20362
rect 17788 20304 23110 20360
rect 23166 20304 23171 20360
rect 17788 20302 23171 20304
rect 17788 20300 17794 20302
rect 23105 20299 23171 20302
rect 17861 20226 17927 20229
rect 21357 20226 21423 20229
rect 17861 20224 21423 20226
rect 17861 20168 17866 20224
rect 17922 20168 21362 20224
rect 21418 20168 21423 20224
rect 17861 20166 21423 20168
rect 17861 20163 17927 20166
rect 21357 20163 21423 20166
rect 21541 20226 21607 20229
rect 22277 20226 22343 20229
rect 21541 20224 22343 20226
rect 21541 20168 21546 20224
rect 21602 20168 22282 20224
rect 22338 20168 22343 20224
rect 21541 20166 22343 20168
rect 21541 20163 21607 20166
rect 22277 20163 22343 20166
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 15942 20160 16258 20161
rect 15942 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16258 20160
rect 15942 20095 16258 20096
rect 23716 20160 24032 20161
rect 23716 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24032 20160
rect 23716 20095 24032 20096
rect 31490 20160 31806 20161
rect 31490 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31806 20160
rect 31490 20095 31806 20096
rect 19241 20090 19307 20093
rect 21081 20090 21147 20093
rect 19241 20088 21147 20090
rect 19241 20032 19246 20088
rect 19302 20032 21086 20088
rect 21142 20032 21147 20088
rect 19241 20030 21147 20032
rect 19241 20027 19307 20030
rect 21081 20027 21147 20030
rect 10777 19954 10843 19957
rect 18689 19954 18755 19957
rect 10777 19952 18755 19954
rect 10777 19896 10782 19952
rect 10838 19896 18694 19952
rect 18750 19896 18755 19952
rect 10777 19894 18755 19896
rect 10777 19891 10843 19894
rect 18689 19891 18755 19894
rect 19701 19954 19767 19957
rect 21357 19954 21423 19957
rect 19701 19952 21423 19954
rect 19701 19896 19706 19952
rect 19762 19896 21362 19952
rect 21418 19896 21423 19952
rect 19701 19894 21423 19896
rect 19701 19891 19767 19894
rect 21357 19891 21423 19894
rect 15101 19818 15167 19821
rect 22737 19818 22803 19821
rect 15101 19816 22803 19818
rect 15101 19760 15106 19816
rect 15162 19760 22742 19816
rect 22798 19760 22803 19816
rect 15101 19758 22803 19760
rect 15101 19755 15167 19758
rect 22737 19755 22803 19758
rect 23013 19818 23079 19821
rect 27337 19818 27403 19821
rect 23013 19816 27403 19818
rect 23013 19760 23018 19816
rect 23074 19760 27342 19816
rect 27398 19760 27403 19816
rect 23013 19758 27403 19760
rect 23013 19755 23079 19758
rect 27337 19755 27403 19758
rect 10133 19684 10199 19685
rect 10133 19682 10180 19684
rect 10088 19680 10180 19682
rect 10088 19624 10138 19680
rect 10088 19622 10180 19624
rect 10133 19620 10180 19622
rect 10244 19620 10250 19684
rect 17769 19682 17835 19685
rect 15150 19680 17835 19682
rect 15150 19624 17774 19680
rect 17830 19624 17835 19680
rect 15150 19622 17835 19624
rect 10133 19619 10199 19620
rect 4281 19616 4597 19617
rect 4281 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4597 19616
rect 4281 19551 4597 19552
rect 12055 19616 12371 19617
rect 12055 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12371 19616
rect 12055 19551 12371 19552
rect 6545 19546 6611 19549
rect 11145 19546 11211 19549
rect 6545 19544 11211 19546
rect 6545 19488 6550 19544
rect 6606 19488 11150 19544
rect 11206 19488 11211 19544
rect 6545 19486 11211 19488
rect 6545 19483 6611 19486
rect 11145 19483 11211 19486
rect 4245 19410 4311 19413
rect 5390 19410 5396 19412
rect 4245 19408 5396 19410
rect 4245 19352 4250 19408
rect 4306 19352 5396 19408
rect 4245 19350 5396 19352
rect 4245 19347 4311 19350
rect 5390 19348 5396 19350
rect 5460 19348 5466 19412
rect 9489 19410 9555 19413
rect 10041 19410 10107 19413
rect 13261 19410 13327 19413
rect 13486 19410 13492 19412
rect 9489 19408 13492 19410
rect 9489 19352 9494 19408
rect 9550 19352 10046 19408
rect 10102 19352 13266 19408
rect 13322 19352 13492 19408
rect 9489 19350 13492 19352
rect 9489 19347 9555 19350
rect 10041 19347 10107 19350
rect 13261 19347 13327 19350
rect 13486 19348 13492 19350
rect 13556 19348 13562 19412
rect 15150 19410 15210 19622
rect 17769 19619 17835 19622
rect 18597 19682 18663 19685
rect 18873 19682 18939 19685
rect 18597 19680 18939 19682
rect 18597 19624 18602 19680
rect 18658 19624 18878 19680
rect 18934 19624 18939 19680
rect 18597 19622 18939 19624
rect 18597 19619 18663 19622
rect 18873 19619 18939 19622
rect 21357 19682 21423 19685
rect 26325 19682 26391 19685
rect 21357 19680 26391 19682
rect 21357 19624 21362 19680
rect 21418 19624 26330 19680
rect 26386 19624 26391 19680
rect 21357 19622 26391 19624
rect 21357 19619 21423 19622
rect 26325 19619 26391 19622
rect 19829 19616 20145 19617
rect 19829 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20145 19616
rect 19829 19551 20145 19552
rect 27603 19616 27919 19617
rect 27603 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27919 19616
rect 27603 19551 27919 19552
rect 17217 19546 17283 19549
rect 21449 19548 21515 19549
rect 17217 19544 18154 19546
rect 17217 19488 17222 19544
rect 17278 19488 18154 19544
rect 17217 19486 18154 19488
rect 17217 19483 17283 19486
rect 13678 19350 15210 19410
rect 16573 19410 16639 19413
rect 18094 19410 18154 19486
rect 21398 19484 21404 19548
rect 21468 19546 21515 19548
rect 21909 19548 21975 19549
rect 23473 19548 23539 19549
rect 21468 19544 21560 19546
rect 21510 19488 21560 19544
rect 21468 19486 21560 19488
rect 21909 19544 21956 19548
rect 22020 19546 22026 19548
rect 23422 19546 23428 19548
rect 21909 19488 21914 19544
rect 21468 19484 21515 19486
rect 21449 19483 21515 19484
rect 21909 19484 21956 19488
rect 22020 19486 22066 19546
rect 23382 19486 23428 19546
rect 23492 19544 23539 19548
rect 23534 19488 23539 19544
rect 22020 19484 22026 19486
rect 23422 19484 23428 19486
rect 23492 19484 23539 19488
rect 21909 19483 21975 19484
rect 23473 19483 23539 19484
rect 24761 19546 24827 19549
rect 27061 19546 27127 19549
rect 24761 19544 27127 19546
rect 24761 19488 24766 19544
rect 24822 19488 27066 19544
rect 27122 19488 27127 19544
rect 24761 19486 27127 19488
rect 24761 19483 24827 19486
rect 27061 19483 27127 19486
rect 26693 19410 26759 19413
rect 16573 19408 17970 19410
rect 16573 19352 16578 19408
rect 16634 19352 17970 19408
rect 16573 19350 17970 19352
rect 18094 19408 26759 19410
rect 18094 19352 26698 19408
rect 26754 19352 26759 19408
rect 18094 19350 26759 19352
rect 5206 19212 5212 19276
rect 5276 19274 5282 19276
rect 6637 19274 6703 19277
rect 5276 19272 6703 19274
rect 5276 19216 6642 19272
rect 6698 19216 6703 19272
rect 5276 19214 6703 19216
rect 5276 19212 5282 19214
rect 6637 19211 6703 19214
rect 10685 19274 10751 19277
rect 11094 19274 11100 19276
rect 10685 19272 11100 19274
rect 10685 19216 10690 19272
rect 10746 19216 11100 19272
rect 10685 19214 11100 19216
rect 10685 19211 10751 19214
rect 11094 19212 11100 19214
rect 11164 19212 11170 19276
rect 11421 19274 11487 19277
rect 13678 19274 13738 19350
rect 16573 19347 16639 19350
rect 11421 19272 13738 19274
rect 11421 19216 11426 19272
rect 11482 19216 13738 19272
rect 11421 19214 13738 19216
rect 13905 19274 13971 19277
rect 17217 19274 17283 19277
rect 13905 19272 17283 19274
rect 13905 19216 13910 19272
rect 13966 19216 17222 19272
rect 17278 19216 17283 19272
rect 13905 19214 17283 19216
rect 17910 19274 17970 19350
rect 26693 19347 26759 19350
rect 26969 19410 27035 19413
rect 27102 19410 27108 19412
rect 26969 19408 27108 19410
rect 26969 19352 26974 19408
rect 27030 19352 27108 19408
rect 26969 19350 27108 19352
rect 26969 19347 27035 19350
rect 27102 19348 27108 19350
rect 27172 19348 27178 19412
rect 28901 19274 28967 19277
rect 17910 19272 28967 19274
rect 17910 19216 28906 19272
rect 28962 19216 28967 19272
rect 17910 19214 28967 19216
rect 11421 19211 11487 19214
rect 13905 19211 13971 19214
rect 17217 19211 17283 19214
rect 28901 19211 28967 19214
rect 11605 19138 11671 19141
rect 15285 19138 15351 19141
rect 11605 19136 15351 19138
rect 11605 19080 11610 19136
rect 11666 19080 15290 19136
rect 15346 19080 15351 19136
rect 11605 19078 15351 19080
rect 11605 19075 11671 19078
rect 15285 19075 15351 19078
rect 16757 19138 16823 19141
rect 20805 19138 20871 19141
rect 23197 19138 23263 19141
rect 16757 19136 23263 19138
rect 16757 19080 16762 19136
rect 16818 19080 20810 19136
rect 20866 19080 23202 19136
rect 23258 19080 23263 19136
rect 16757 19078 23263 19080
rect 16757 19075 16823 19078
rect 20805 19075 20871 19078
rect 23197 19075 23263 19078
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 15942 19072 16258 19073
rect 15942 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16258 19072
rect 15942 19007 16258 19008
rect 23716 19072 24032 19073
rect 23716 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24032 19072
rect 23716 19007 24032 19008
rect 31490 19072 31806 19073
rect 31490 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31806 19072
rect 31490 19007 31806 19008
rect 11145 19002 11211 19005
rect 13721 19002 13787 19005
rect 15193 19002 15259 19005
rect 11145 19000 11898 19002
rect 11145 18944 11150 19000
rect 11206 18944 11898 19000
rect 11145 18942 11898 18944
rect 11145 18939 11211 18942
rect 2497 18866 2563 18869
rect 4337 18866 4403 18869
rect 11513 18866 11579 18869
rect 11838 18868 11898 18942
rect 13721 19000 15259 19002
rect 13721 18944 13726 19000
rect 13782 18944 15198 19000
rect 15254 18944 15259 19000
rect 13721 18942 15259 18944
rect 13721 18939 13787 18942
rect 15193 18939 15259 18942
rect 16665 19002 16731 19005
rect 16798 19002 16804 19004
rect 16665 19000 16804 19002
rect 16665 18944 16670 19000
rect 16726 18944 16804 19000
rect 16665 18942 16804 18944
rect 16665 18939 16731 18942
rect 16798 18940 16804 18942
rect 16868 18940 16874 19004
rect 17217 19002 17283 19005
rect 20253 19002 20319 19005
rect 20478 19002 20484 19004
rect 17217 19000 19810 19002
rect 17217 18944 17222 19000
rect 17278 18944 19810 19000
rect 17217 18942 19810 18944
rect 17217 18939 17283 18942
rect 2497 18864 11579 18866
rect 2497 18808 2502 18864
rect 2558 18808 4342 18864
rect 4398 18808 11518 18864
rect 11574 18808 11579 18864
rect 2497 18806 11579 18808
rect 2497 18803 2563 18806
rect 4337 18803 4403 18806
rect 11513 18803 11579 18806
rect 11830 18804 11836 18868
rect 11900 18804 11906 18868
rect 18505 18866 18571 18869
rect 19425 18866 19491 18869
rect 18505 18864 19491 18866
rect 18505 18808 18510 18864
rect 18566 18808 19430 18864
rect 19486 18808 19491 18864
rect 18505 18806 19491 18808
rect 19750 18866 19810 18942
rect 20253 19000 20484 19002
rect 20253 18944 20258 19000
rect 20314 18944 20484 19000
rect 20253 18942 20484 18944
rect 20253 18939 20319 18942
rect 20478 18940 20484 18942
rect 20548 18940 20554 19004
rect 20621 19002 20687 19005
rect 21449 19002 21515 19005
rect 20621 19000 21515 19002
rect 20621 18944 20626 19000
rect 20682 18944 21454 19000
rect 21510 18944 21515 19000
rect 20621 18942 21515 18944
rect 20621 18939 20687 18942
rect 21449 18939 21515 18942
rect 29177 18866 29243 18869
rect 19750 18864 29243 18866
rect 19750 18808 29182 18864
rect 29238 18808 29243 18864
rect 19750 18806 29243 18808
rect 18505 18803 18571 18806
rect 19425 18803 19491 18806
rect 29177 18803 29243 18806
rect 4245 18730 4311 18733
rect 5901 18730 5967 18733
rect 9121 18730 9187 18733
rect 4245 18728 9187 18730
rect 4245 18672 4250 18728
rect 4306 18672 5906 18728
rect 5962 18672 9126 18728
rect 9182 18672 9187 18728
rect 4245 18670 9187 18672
rect 4245 18667 4311 18670
rect 5901 18667 5967 18670
rect 9121 18667 9187 18670
rect 11053 18730 11119 18733
rect 24945 18730 25011 18733
rect 11053 18728 25011 18730
rect 11053 18672 11058 18728
rect 11114 18672 24950 18728
rect 25006 18672 25011 18728
rect 11053 18670 25011 18672
rect 11053 18667 11119 18670
rect 24945 18667 25011 18670
rect 14273 18594 14339 18597
rect 16849 18594 16915 18597
rect 14273 18592 16915 18594
rect 14273 18536 14278 18592
rect 14334 18536 16854 18592
rect 16910 18536 16915 18592
rect 14273 18534 16915 18536
rect 14273 18531 14339 18534
rect 16849 18531 16915 18534
rect 4281 18528 4597 18529
rect 4281 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4597 18528
rect 4281 18463 4597 18464
rect 12055 18528 12371 18529
rect 12055 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12371 18528
rect 12055 18463 12371 18464
rect 19829 18528 20145 18529
rect 19829 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20145 18528
rect 19829 18463 20145 18464
rect 27603 18528 27919 18529
rect 27603 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27919 18528
rect 27603 18463 27919 18464
rect 12985 18458 13051 18461
rect 14641 18458 14707 18461
rect 12985 18456 14707 18458
rect 12985 18400 12990 18456
rect 13046 18400 14646 18456
rect 14702 18400 14707 18456
rect 12985 18398 14707 18400
rect 12985 18395 13051 18398
rect 14641 18395 14707 18398
rect 16665 18458 16731 18461
rect 19333 18458 19399 18461
rect 16665 18456 19399 18458
rect 16665 18400 16670 18456
rect 16726 18400 19338 18456
rect 19394 18400 19399 18456
rect 16665 18398 19399 18400
rect 16665 18395 16731 18398
rect 19333 18395 19399 18398
rect 20253 18458 20319 18461
rect 21265 18458 21331 18461
rect 20253 18456 21331 18458
rect 20253 18400 20258 18456
rect 20314 18400 21270 18456
rect 21326 18400 21331 18456
rect 20253 18398 21331 18400
rect 20253 18395 20319 18398
rect 21265 18395 21331 18398
rect 5441 18322 5507 18325
rect 7649 18322 7715 18325
rect 9029 18322 9095 18325
rect 5441 18320 9095 18322
rect 5441 18264 5446 18320
rect 5502 18264 7654 18320
rect 7710 18264 9034 18320
rect 9090 18264 9095 18320
rect 5441 18262 9095 18264
rect 5441 18259 5507 18262
rect 7649 18259 7715 18262
rect 9029 18259 9095 18262
rect 9806 18260 9812 18324
rect 9876 18322 9882 18324
rect 9949 18322 10015 18325
rect 9876 18320 10015 18322
rect 9876 18264 9954 18320
rect 10010 18264 10015 18320
rect 9876 18262 10015 18264
rect 9876 18260 9882 18262
rect 9949 18259 10015 18262
rect 13353 18322 13419 18325
rect 16389 18322 16455 18325
rect 13353 18320 16455 18322
rect 13353 18264 13358 18320
rect 13414 18264 16394 18320
rect 16450 18264 16455 18320
rect 13353 18262 16455 18264
rect 13353 18259 13419 18262
rect 16389 18259 16455 18262
rect 19149 18322 19215 18325
rect 20161 18322 20227 18325
rect 19149 18320 20227 18322
rect 19149 18264 19154 18320
rect 19210 18264 20166 18320
rect 20222 18264 20227 18320
rect 19149 18262 20227 18264
rect 19149 18259 19215 18262
rect 20161 18259 20227 18262
rect 22921 18322 22987 18325
rect 27797 18322 27863 18325
rect 22921 18320 27863 18322
rect 22921 18264 22926 18320
rect 22982 18264 27802 18320
rect 27858 18264 27863 18320
rect 22921 18262 27863 18264
rect 22921 18259 22987 18262
rect 27797 18259 27863 18262
rect 3785 18186 3851 18189
rect 4429 18186 4495 18189
rect 3785 18184 4495 18186
rect 3785 18128 3790 18184
rect 3846 18128 4434 18184
rect 4490 18128 4495 18184
rect 3785 18126 4495 18128
rect 3785 18123 3851 18126
rect 4429 18123 4495 18126
rect 6453 18186 6519 18189
rect 13353 18186 13419 18189
rect 6453 18184 13419 18186
rect 6453 18128 6458 18184
rect 6514 18128 13358 18184
rect 13414 18128 13419 18184
rect 6453 18126 13419 18128
rect 6453 18123 6519 18126
rect 13353 18123 13419 18126
rect 17861 18186 17927 18189
rect 18270 18186 18276 18188
rect 17861 18184 18276 18186
rect 17861 18128 17866 18184
rect 17922 18128 18276 18184
rect 17861 18126 18276 18128
rect 17861 18123 17927 18126
rect 18270 18124 18276 18126
rect 18340 18186 18346 18188
rect 24669 18186 24735 18189
rect 28349 18186 28415 18189
rect 18340 18184 28415 18186
rect 18340 18128 24674 18184
rect 24730 18128 28354 18184
rect 28410 18128 28415 18184
rect 18340 18126 28415 18128
rect 18340 18124 18346 18126
rect 24669 18123 24735 18126
rect 28349 18123 28415 18126
rect 2681 18050 2747 18053
rect 3969 18050 4035 18053
rect 2681 18048 4035 18050
rect 2681 17992 2686 18048
rect 2742 17992 3974 18048
rect 4030 17992 4035 18048
rect 2681 17990 4035 17992
rect 2681 17987 2747 17990
rect 3969 17987 4035 17990
rect 8569 18050 8635 18053
rect 10869 18050 10935 18053
rect 8569 18048 10935 18050
rect 8569 17992 8574 18048
rect 8630 17992 10874 18048
rect 10930 17992 10935 18048
rect 8569 17990 10935 17992
rect 8569 17987 8635 17990
rect 10869 17987 10935 17990
rect 11789 18050 11855 18053
rect 14641 18050 14707 18053
rect 11789 18048 14707 18050
rect 11789 17992 11794 18048
rect 11850 17992 14646 18048
rect 14702 17992 14707 18048
rect 11789 17990 14707 17992
rect 11789 17987 11855 17990
rect 14641 17987 14707 17990
rect 16573 18050 16639 18053
rect 18638 18050 18644 18052
rect 16573 18048 18644 18050
rect 16573 17992 16578 18048
rect 16634 17992 18644 18048
rect 16573 17990 18644 17992
rect 16573 17987 16639 17990
rect 18638 17988 18644 17990
rect 18708 18050 18714 18052
rect 18965 18050 19031 18053
rect 18708 18048 19031 18050
rect 18708 17992 18970 18048
rect 19026 17992 19031 18048
rect 18708 17990 19031 17992
rect 18708 17988 18714 17990
rect 18965 17987 19031 17990
rect 19425 18050 19491 18053
rect 22645 18050 22711 18053
rect 19425 18048 22711 18050
rect 19425 17992 19430 18048
rect 19486 17992 22650 18048
rect 22706 17992 22711 18048
rect 19425 17990 22711 17992
rect 19425 17987 19491 17990
rect 22645 17987 22711 17990
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 15942 17984 16258 17985
rect 15942 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16258 17984
rect 15942 17919 16258 17920
rect 23716 17984 24032 17985
rect 23716 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24032 17984
rect 23716 17919 24032 17920
rect 31490 17984 31806 17985
rect 31490 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31806 17984
rect 31490 17919 31806 17920
rect 10133 17914 10199 17917
rect 8710 17912 10199 17914
rect 8710 17856 10138 17912
rect 10194 17856 10199 17912
rect 8710 17854 10199 17856
rect 8109 17778 8175 17781
rect 8710 17778 8770 17854
rect 10133 17851 10199 17854
rect 11145 17914 11211 17917
rect 11973 17914 12039 17917
rect 11145 17912 12039 17914
rect 11145 17856 11150 17912
rect 11206 17856 11978 17912
rect 12034 17856 12039 17912
rect 11145 17854 12039 17856
rect 11145 17851 11211 17854
rect 11973 17851 12039 17854
rect 16573 17914 16639 17917
rect 18965 17914 19031 17917
rect 16573 17912 19031 17914
rect 16573 17856 16578 17912
rect 16634 17856 18970 17912
rect 19026 17856 19031 17912
rect 16573 17854 19031 17856
rect 16573 17851 16639 17854
rect 18965 17851 19031 17854
rect 19425 17914 19491 17917
rect 23565 17914 23631 17917
rect 19425 17912 23631 17914
rect 19425 17856 19430 17912
rect 19486 17856 23570 17912
rect 23626 17856 23631 17912
rect 19425 17854 23631 17856
rect 19425 17851 19491 17854
rect 23565 17851 23631 17854
rect 24301 17914 24367 17917
rect 30189 17914 30255 17917
rect 24301 17912 30255 17914
rect 24301 17856 24306 17912
rect 24362 17856 30194 17912
rect 30250 17856 30255 17912
rect 24301 17854 30255 17856
rect 24301 17851 24367 17854
rect 30189 17851 30255 17854
rect 8109 17776 8770 17778
rect 8109 17720 8114 17776
rect 8170 17720 8770 17776
rect 8109 17718 8770 17720
rect 10133 17778 10199 17781
rect 11237 17778 11303 17781
rect 10133 17776 11303 17778
rect 10133 17720 10138 17776
rect 10194 17720 11242 17776
rect 11298 17720 11303 17776
rect 10133 17718 11303 17720
rect 8109 17715 8175 17718
rect 10133 17715 10199 17718
rect 11237 17715 11303 17718
rect 13537 17778 13603 17781
rect 15653 17778 15719 17781
rect 13537 17776 15719 17778
rect 13537 17720 13542 17776
rect 13598 17720 15658 17776
rect 15714 17720 15719 17776
rect 13537 17718 15719 17720
rect 13537 17715 13603 17718
rect 15653 17715 15719 17718
rect 16757 17778 16823 17781
rect 17769 17778 17835 17781
rect 24853 17778 24919 17781
rect 16757 17776 24919 17778
rect 16757 17720 16762 17776
rect 16818 17720 17774 17776
rect 17830 17720 24858 17776
rect 24914 17720 24919 17776
rect 16757 17718 24919 17720
rect 16757 17715 16823 17718
rect 17769 17715 17835 17718
rect 24853 17715 24919 17718
rect 5441 17642 5507 17645
rect 14089 17642 14155 17645
rect 18505 17642 18571 17645
rect 19333 17642 19399 17645
rect 21357 17642 21423 17645
rect 21633 17642 21699 17645
rect 5441 17640 17786 17642
rect 5441 17584 5446 17640
rect 5502 17584 14094 17640
rect 14150 17584 17786 17640
rect 5441 17582 17786 17584
rect 5441 17579 5507 17582
rect 14089 17579 14155 17582
rect 7833 17506 7899 17509
rect 10961 17506 11027 17509
rect 7833 17504 11027 17506
rect 7833 17448 7838 17504
rect 7894 17448 10966 17504
rect 11022 17448 11027 17504
rect 7833 17446 11027 17448
rect 17726 17506 17786 17582
rect 18505 17640 19399 17642
rect 18505 17584 18510 17640
rect 18566 17584 19338 17640
rect 19394 17584 19399 17640
rect 18505 17582 19399 17584
rect 18505 17579 18571 17582
rect 19333 17579 19399 17582
rect 19566 17640 21699 17642
rect 19566 17584 21362 17640
rect 21418 17584 21638 17640
rect 21694 17584 21699 17640
rect 19566 17582 21699 17584
rect 19566 17506 19626 17582
rect 21357 17579 21423 17582
rect 21633 17579 21699 17582
rect 23289 17642 23355 17645
rect 26601 17642 26667 17645
rect 23289 17640 26667 17642
rect 23289 17584 23294 17640
rect 23350 17584 26606 17640
rect 26662 17584 26667 17640
rect 23289 17582 26667 17584
rect 23289 17579 23355 17582
rect 26601 17579 26667 17582
rect 17726 17446 19626 17506
rect 20529 17506 20595 17509
rect 24209 17506 24275 17509
rect 20529 17504 24275 17506
rect 20529 17448 20534 17504
rect 20590 17448 24214 17504
rect 24270 17448 24275 17504
rect 20529 17446 24275 17448
rect 7833 17443 7899 17446
rect 10961 17443 11027 17446
rect 20529 17443 20595 17446
rect 24209 17443 24275 17446
rect 4281 17440 4597 17441
rect 4281 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4597 17440
rect 4281 17375 4597 17376
rect 12055 17440 12371 17441
rect 12055 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12371 17440
rect 12055 17375 12371 17376
rect 19829 17440 20145 17441
rect 19829 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20145 17440
rect 19829 17375 20145 17376
rect 27603 17440 27919 17441
rect 27603 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27919 17440
rect 27603 17375 27919 17376
rect 9213 17370 9279 17373
rect 10501 17370 10567 17373
rect 9213 17368 10567 17370
rect 9213 17312 9218 17368
rect 9274 17312 10506 17368
rect 10562 17312 10567 17368
rect 9213 17310 10567 17312
rect 9213 17307 9279 17310
rect 10501 17307 10567 17310
rect 14641 17370 14707 17373
rect 15285 17370 15351 17373
rect 17125 17372 17191 17373
rect 17125 17370 17172 17372
rect 14641 17368 17172 17370
rect 14641 17312 14646 17368
rect 14702 17312 15290 17368
rect 15346 17312 17130 17368
rect 14641 17310 17172 17312
rect 14641 17307 14707 17310
rect 15285 17307 15351 17310
rect 17125 17308 17172 17310
rect 17236 17308 17242 17372
rect 18137 17368 18203 17373
rect 18137 17312 18142 17368
rect 18198 17312 18203 17368
rect 17125 17307 17191 17308
rect 18137 17307 18203 17312
rect 20253 17370 20319 17373
rect 24853 17370 24919 17373
rect 20253 17368 24919 17370
rect 20253 17312 20258 17368
rect 20314 17312 24858 17368
rect 24914 17312 24919 17368
rect 20253 17310 24919 17312
rect 20253 17307 20319 17310
rect 24853 17307 24919 17310
rect 5073 17234 5139 17237
rect 10726 17234 10732 17236
rect 5073 17232 10732 17234
rect 5073 17176 5078 17232
rect 5134 17176 10732 17232
rect 5073 17174 10732 17176
rect 5073 17171 5139 17174
rect 10726 17172 10732 17174
rect 10796 17234 10802 17236
rect 10869 17234 10935 17237
rect 10796 17232 10935 17234
rect 10796 17176 10874 17232
rect 10930 17176 10935 17232
rect 10796 17174 10935 17176
rect 10796 17172 10802 17174
rect 10869 17171 10935 17174
rect 17217 17234 17283 17237
rect 18140 17234 18200 17307
rect 19609 17236 19675 17237
rect 19558 17234 19564 17236
rect 17217 17232 18200 17234
rect 17217 17176 17222 17232
rect 17278 17176 18200 17232
rect 17217 17174 18200 17176
rect 19518 17174 19564 17234
rect 19628 17232 19675 17236
rect 19670 17176 19675 17232
rect 17217 17171 17283 17174
rect 19558 17172 19564 17174
rect 19628 17172 19675 17176
rect 19609 17171 19675 17172
rect 19885 17234 19951 17237
rect 24025 17234 24091 17237
rect 19885 17232 24091 17234
rect 19885 17176 19890 17232
rect 19946 17176 24030 17232
rect 24086 17176 24091 17232
rect 19885 17174 24091 17176
rect 19885 17171 19951 17174
rect 24025 17171 24091 17174
rect 8477 17098 8543 17101
rect 11973 17098 12039 17101
rect 20621 17098 20687 17101
rect 22277 17098 22343 17101
rect 22553 17098 22619 17101
rect 26233 17098 26299 17101
rect 8477 17096 11898 17098
rect 8477 17040 8482 17096
rect 8538 17040 11898 17096
rect 8477 17038 11898 17040
rect 8477 17035 8543 17038
rect 9305 16962 9371 16965
rect 10961 16962 11027 16965
rect 9305 16960 11027 16962
rect 9305 16904 9310 16960
rect 9366 16904 10966 16960
rect 11022 16904 11027 16960
rect 9305 16902 11027 16904
rect 11838 16962 11898 17038
rect 11973 17096 20687 17098
rect 11973 17040 11978 17096
rect 12034 17040 20626 17096
rect 20682 17040 20687 17096
rect 11973 17038 20687 17040
rect 11973 17035 12039 17038
rect 20621 17035 20687 17038
rect 20808 17096 22343 17098
rect 20808 17040 22282 17096
rect 22338 17040 22343 17096
rect 20808 17038 22343 17040
rect 11973 16962 12039 16965
rect 11838 16960 12039 16962
rect 11838 16904 11978 16960
rect 12034 16904 12039 16960
rect 11838 16902 12039 16904
rect 9305 16899 9371 16902
rect 10961 16899 11027 16902
rect 11973 16899 12039 16902
rect 18413 16962 18479 16965
rect 18873 16962 18939 16965
rect 20808 16962 20868 17038
rect 22277 17035 22343 17038
rect 22510 17096 26299 17098
rect 22510 17040 22558 17096
rect 22614 17040 26238 17096
rect 26294 17040 26299 17096
rect 22510 17038 26299 17040
rect 22510 17035 22619 17038
rect 26233 17035 26299 17038
rect 18413 16960 20868 16962
rect 18413 16904 18418 16960
rect 18474 16904 18878 16960
rect 18934 16904 20868 16960
rect 18413 16902 20868 16904
rect 20989 16962 21055 16965
rect 22510 16962 22570 17035
rect 20989 16960 22570 16962
rect 20989 16904 20994 16960
rect 21050 16904 22570 16960
rect 20989 16902 22570 16904
rect 25313 16962 25379 16965
rect 26969 16962 27035 16965
rect 25313 16960 27035 16962
rect 25313 16904 25318 16960
rect 25374 16904 26974 16960
rect 27030 16904 27035 16960
rect 25313 16902 27035 16904
rect 18413 16899 18479 16902
rect 18873 16899 18939 16902
rect 20989 16899 21055 16902
rect 25313 16899 25379 16902
rect 26969 16899 27035 16902
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 15942 16896 16258 16897
rect 15942 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16258 16896
rect 15942 16831 16258 16832
rect 23716 16896 24032 16897
rect 23716 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24032 16896
rect 23716 16831 24032 16832
rect 31490 16896 31806 16897
rect 31490 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31806 16896
rect 31490 16831 31806 16832
rect 9397 16826 9463 16829
rect 9622 16826 9628 16828
rect 9397 16824 9628 16826
rect 9397 16768 9402 16824
rect 9458 16768 9628 16824
rect 9397 16766 9628 16768
rect 9397 16763 9463 16766
rect 9622 16764 9628 16766
rect 9692 16764 9698 16828
rect 16481 16826 16547 16829
rect 17493 16826 17559 16829
rect 22277 16826 22343 16829
rect 16481 16824 22343 16826
rect 16481 16768 16486 16824
rect 16542 16768 17498 16824
rect 17554 16768 22282 16824
rect 22338 16768 22343 16824
rect 16481 16766 22343 16768
rect 16481 16763 16547 16766
rect 17493 16763 17559 16766
rect 22277 16763 22343 16766
rect 24117 16826 24183 16829
rect 25221 16826 25287 16829
rect 24117 16824 25287 16826
rect 24117 16768 24122 16824
rect 24178 16768 25226 16824
rect 25282 16768 25287 16824
rect 24117 16766 25287 16768
rect 24117 16763 24183 16766
rect 25221 16763 25287 16766
rect 6637 16690 6703 16693
rect 10593 16690 10659 16693
rect 6637 16688 10659 16690
rect 6637 16632 6642 16688
rect 6698 16632 10598 16688
rect 10654 16632 10659 16688
rect 6637 16630 10659 16632
rect 6637 16627 6703 16630
rect 10593 16627 10659 16630
rect 11789 16690 11855 16693
rect 13537 16690 13603 16693
rect 11789 16688 13603 16690
rect 11789 16632 11794 16688
rect 11850 16632 13542 16688
rect 13598 16632 13603 16688
rect 11789 16630 13603 16632
rect 11789 16627 11855 16630
rect 13537 16627 13603 16630
rect 16573 16690 16639 16693
rect 28717 16690 28783 16693
rect 16573 16688 28783 16690
rect 16573 16632 16578 16688
rect 16634 16632 28722 16688
rect 28778 16632 28783 16688
rect 16573 16630 28783 16632
rect 16573 16627 16639 16630
rect 28717 16627 28783 16630
rect 12065 16554 12131 16557
rect 16941 16554 17007 16557
rect 12065 16552 17007 16554
rect 12065 16496 12070 16552
rect 12126 16496 16946 16552
rect 17002 16496 17007 16552
rect 12065 16494 17007 16496
rect 12065 16491 12131 16494
rect 16941 16491 17007 16494
rect 21265 16554 21331 16557
rect 21398 16554 21404 16556
rect 21265 16552 21404 16554
rect 21265 16496 21270 16552
rect 21326 16496 21404 16552
rect 21265 16494 21404 16496
rect 21265 16491 21331 16494
rect 21398 16492 21404 16494
rect 21468 16492 21474 16556
rect 21909 16554 21975 16557
rect 23933 16554 23999 16557
rect 21909 16552 23999 16554
rect 21909 16496 21914 16552
rect 21970 16496 23938 16552
rect 23994 16496 23999 16552
rect 21909 16494 23999 16496
rect 21909 16491 21975 16494
rect 23933 16491 23999 16494
rect 8477 16418 8543 16421
rect 10685 16418 10751 16421
rect 8477 16416 10751 16418
rect 8477 16360 8482 16416
rect 8538 16360 10690 16416
rect 10746 16360 10751 16416
rect 8477 16358 10751 16360
rect 8477 16355 8543 16358
rect 10685 16355 10751 16358
rect 13486 16356 13492 16420
rect 13556 16418 13562 16420
rect 14457 16418 14523 16421
rect 13556 16416 14523 16418
rect 13556 16360 14462 16416
rect 14518 16360 14523 16416
rect 13556 16358 14523 16360
rect 13556 16356 13562 16358
rect 14457 16355 14523 16358
rect 16665 16418 16731 16421
rect 17861 16418 17927 16421
rect 16665 16416 17927 16418
rect 16665 16360 16670 16416
rect 16726 16360 17866 16416
rect 17922 16360 17927 16416
rect 16665 16358 17927 16360
rect 16665 16355 16731 16358
rect 17861 16355 17927 16358
rect 21541 16418 21607 16421
rect 26325 16418 26391 16421
rect 21541 16416 26391 16418
rect 21541 16360 21546 16416
rect 21602 16360 26330 16416
rect 26386 16360 26391 16416
rect 21541 16358 26391 16360
rect 21541 16355 21607 16358
rect 26325 16355 26391 16358
rect 4281 16352 4597 16353
rect 4281 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4597 16352
rect 4281 16287 4597 16288
rect 12055 16352 12371 16353
rect 12055 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12371 16352
rect 12055 16287 12371 16288
rect 19829 16352 20145 16353
rect 19829 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20145 16352
rect 19829 16287 20145 16288
rect 27603 16352 27919 16353
rect 27603 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27919 16352
rect 27603 16287 27919 16288
rect 18822 16282 18828 16284
rect 14598 16222 18828 16282
rect 5349 16146 5415 16149
rect 10409 16146 10475 16149
rect 5349 16144 10475 16146
rect 5349 16088 5354 16144
rect 5410 16088 10414 16144
rect 10470 16088 10475 16144
rect 5349 16086 10475 16088
rect 5349 16083 5415 16086
rect 10409 16083 10475 16086
rect 11605 16146 11671 16149
rect 14598 16146 14658 16222
rect 18822 16220 18828 16222
rect 18892 16282 18898 16284
rect 19609 16282 19675 16285
rect 18892 16280 19675 16282
rect 18892 16224 19614 16280
rect 19670 16224 19675 16280
rect 18892 16222 19675 16224
rect 18892 16220 18898 16222
rect 19609 16219 19675 16222
rect 20437 16282 20503 16285
rect 27061 16282 27127 16285
rect 20437 16280 27127 16282
rect 20437 16224 20442 16280
rect 20498 16224 27066 16280
rect 27122 16224 27127 16280
rect 20437 16222 27127 16224
rect 20437 16219 20503 16222
rect 27061 16219 27127 16222
rect 11605 16144 14658 16146
rect 11605 16088 11610 16144
rect 11666 16088 14658 16144
rect 11605 16086 14658 16088
rect 14733 16146 14799 16149
rect 25497 16146 25563 16149
rect 14733 16144 25563 16146
rect 14733 16088 14738 16144
rect 14794 16088 25502 16144
rect 25558 16088 25563 16144
rect 14733 16086 25563 16088
rect 11605 16083 11671 16086
rect 14733 16083 14799 16086
rect 25497 16083 25563 16086
rect 14917 16010 14983 16013
rect 20713 16010 20779 16013
rect 30966 16010 30972 16012
rect 14917 16008 17464 16010
rect 14917 15952 14922 16008
rect 14978 15952 17464 16008
rect 14917 15950 17464 15952
rect 14917 15947 14983 15950
rect 17404 15877 17464 15950
rect 20713 16008 30972 16010
rect 20713 15952 20718 16008
rect 20774 15952 30972 16008
rect 20713 15950 30972 15952
rect 20713 15947 20779 15950
rect 30966 15948 30972 15950
rect 31036 15948 31042 16012
rect 17401 15874 17467 15877
rect 21173 15874 21239 15877
rect 17401 15872 21239 15874
rect 17401 15816 17406 15872
rect 17462 15816 21178 15872
rect 21234 15816 21239 15872
rect 17401 15814 21239 15816
rect 17401 15811 17467 15814
rect 21173 15811 21239 15814
rect 21541 15874 21607 15877
rect 23565 15874 23631 15877
rect 21541 15872 23631 15874
rect 21541 15816 21546 15872
rect 21602 15816 23570 15872
rect 23626 15816 23631 15872
rect 21541 15814 23631 15816
rect 21541 15811 21607 15814
rect 23565 15811 23631 15814
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 15942 15808 16258 15809
rect 15942 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16258 15808
rect 15942 15743 16258 15744
rect 23716 15808 24032 15809
rect 23716 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24032 15808
rect 23716 15743 24032 15744
rect 31490 15808 31806 15809
rect 31490 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31806 15808
rect 31490 15743 31806 15744
rect 17125 15738 17191 15741
rect 17401 15738 17467 15741
rect 17125 15736 17467 15738
rect 17125 15680 17130 15736
rect 17186 15680 17406 15736
rect 17462 15680 17467 15736
rect 17125 15678 17467 15680
rect 17125 15675 17191 15678
rect 17401 15675 17467 15678
rect 17769 15738 17835 15741
rect 20069 15738 20135 15741
rect 17769 15736 20135 15738
rect 17769 15680 17774 15736
rect 17830 15680 20074 15736
rect 20130 15680 20135 15736
rect 17769 15678 20135 15680
rect 17769 15675 17835 15678
rect 20069 15675 20135 15678
rect 20345 15738 20411 15741
rect 23381 15738 23447 15741
rect 20345 15736 23447 15738
rect 20345 15680 20350 15736
rect 20406 15680 23386 15736
rect 23442 15680 23447 15736
rect 20345 15678 23447 15680
rect 20345 15675 20411 15678
rect 23381 15675 23447 15678
rect 26417 15738 26483 15741
rect 27705 15738 27771 15741
rect 26417 15736 27771 15738
rect 26417 15680 26422 15736
rect 26478 15680 27710 15736
rect 27766 15680 27771 15736
rect 26417 15678 27771 15680
rect 26417 15675 26483 15678
rect 27705 15675 27771 15678
rect 9673 15602 9739 15605
rect 15745 15602 15811 15605
rect 19517 15602 19583 15605
rect 23381 15604 23447 15605
rect 23381 15602 23428 15604
rect 9673 15600 10012 15602
rect 9673 15544 9678 15600
rect 9734 15544 10012 15600
rect 9673 15542 10012 15544
rect 9673 15539 9739 15542
rect 9952 15469 10012 15542
rect 15745 15600 23076 15602
rect 15745 15544 15750 15600
rect 15806 15544 19522 15600
rect 19578 15544 23076 15600
rect 15745 15542 23076 15544
rect 23340 15600 23428 15602
rect 23492 15602 23498 15604
rect 29729 15602 29795 15605
rect 23492 15600 29795 15602
rect 23340 15544 23386 15600
rect 23492 15544 29734 15600
rect 29790 15544 29795 15600
rect 23340 15542 23428 15544
rect 15745 15539 15811 15542
rect 19517 15539 19583 15542
rect 9949 15464 10015 15469
rect 9949 15408 9954 15464
rect 10010 15408 10015 15464
rect 9949 15403 10015 15408
rect 14733 15466 14799 15469
rect 22829 15466 22895 15469
rect 14733 15464 22895 15466
rect 14733 15408 14738 15464
rect 14794 15408 22834 15464
rect 22890 15408 22895 15464
rect 14733 15406 22895 15408
rect 23016 15466 23076 15542
rect 23381 15540 23428 15542
rect 23492 15542 29795 15544
rect 23492 15540 23498 15542
rect 23381 15539 23447 15540
rect 29729 15539 29795 15542
rect 25313 15466 25379 15469
rect 23016 15464 25379 15466
rect 23016 15408 25318 15464
rect 25374 15408 25379 15464
rect 23016 15406 25379 15408
rect 14733 15403 14799 15406
rect 22829 15403 22895 15406
rect 25313 15403 25379 15406
rect 16798 15268 16804 15332
rect 16868 15330 16874 15332
rect 16941 15330 17007 15333
rect 16868 15328 17970 15330
rect 16868 15272 16946 15328
rect 17002 15272 17970 15328
rect 16868 15270 17970 15272
rect 16868 15268 16874 15270
rect 16941 15267 17007 15270
rect 4281 15264 4597 15265
rect 4281 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4597 15264
rect 4281 15199 4597 15200
rect 12055 15264 12371 15265
rect 12055 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12371 15264
rect 12055 15199 12371 15200
rect 7966 15132 7972 15196
rect 8036 15194 8042 15196
rect 8385 15194 8451 15197
rect 8036 15192 8451 15194
rect 8036 15136 8390 15192
rect 8446 15136 8451 15192
rect 8036 15134 8451 15136
rect 8036 15132 8042 15134
rect 8385 15131 8451 15134
rect 8569 15194 8635 15197
rect 9305 15194 9371 15197
rect 11053 15194 11119 15197
rect 8569 15192 11119 15194
rect 8569 15136 8574 15192
rect 8630 15136 9310 15192
rect 9366 15136 11058 15192
rect 11114 15136 11119 15192
rect 8569 15134 11119 15136
rect 17910 15194 17970 15270
rect 18822 15268 18828 15332
rect 18892 15330 18898 15332
rect 18965 15330 19031 15333
rect 18892 15328 19031 15330
rect 18892 15272 18970 15328
rect 19026 15272 19031 15328
rect 18892 15270 19031 15272
rect 18892 15268 18898 15270
rect 18965 15267 19031 15270
rect 20621 15330 20687 15333
rect 24209 15330 24275 15333
rect 20621 15328 24275 15330
rect 20621 15272 20626 15328
rect 20682 15272 24214 15328
rect 24270 15272 24275 15328
rect 20621 15270 24275 15272
rect 20621 15267 20687 15270
rect 24209 15267 24275 15270
rect 24485 15330 24551 15333
rect 26049 15330 26115 15333
rect 24485 15328 26115 15330
rect 24485 15272 24490 15328
rect 24546 15272 26054 15328
rect 26110 15272 26115 15328
rect 24485 15270 26115 15272
rect 24485 15267 24551 15270
rect 26049 15267 26115 15270
rect 19829 15264 20145 15265
rect 19829 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20145 15264
rect 19829 15199 20145 15200
rect 27603 15264 27919 15265
rect 27603 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27919 15264
rect 27603 15199 27919 15200
rect 20529 15194 20595 15197
rect 25865 15194 25931 15197
rect 17910 15134 19626 15194
rect 8569 15131 8635 15134
rect 9305 15131 9371 15134
rect 11053 15131 11119 15134
rect 10961 15058 11027 15061
rect 18689 15058 18755 15061
rect 19566 15060 19626 15134
rect 20302 15192 25931 15194
rect 20302 15136 20534 15192
rect 20590 15136 25870 15192
rect 25926 15136 25931 15192
rect 20302 15134 25931 15136
rect 10961 15056 18755 15058
rect 10961 15000 10966 15056
rect 11022 15000 18694 15056
rect 18750 15000 18755 15056
rect 10961 14998 18755 15000
rect 10961 14995 11027 14998
rect 18689 14995 18755 14998
rect 19558 14996 19564 15060
rect 19628 15058 19634 15060
rect 20302 15058 20362 15134
rect 20529 15131 20595 15134
rect 25865 15131 25931 15134
rect 22001 15060 22067 15061
rect 19628 14998 20362 15058
rect 19628 14996 19634 14998
rect 21950 14996 21956 15060
rect 22020 15058 22067 15060
rect 22829 15058 22895 15061
rect 25681 15058 25747 15061
rect 22020 15056 22112 15058
rect 22062 15000 22112 15056
rect 22020 14998 22112 15000
rect 22829 15056 25747 15058
rect 22829 15000 22834 15056
rect 22890 15000 25686 15056
rect 25742 15000 25747 15056
rect 22829 14998 25747 15000
rect 22020 14996 22067 14998
rect 22001 14995 22067 14996
rect 22829 14995 22895 14998
rect 25681 14995 25747 14998
rect 8937 14922 9003 14925
rect 9806 14922 9812 14924
rect 8937 14920 9812 14922
rect 8937 14864 8942 14920
rect 8998 14864 9812 14920
rect 8937 14862 9812 14864
rect 8937 14859 9003 14862
rect 9806 14860 9812 14862
rect 9876 14922 9882 14924
rect 10777 14922 10843 14925
rect 9876 14920 10843 14922
rect 9876 14864 10782 14920
rect 10838 14864 10843 14920
rect 9876 14862 10843 14864
rect 9876 14860 9882 14862
rect 10777 14859 10843 14862
rect 11881 14922 11947 14925
rect 12525 14922 12591 14925
rect 11881 14920 12591 14922
rect 11881 14864 11886 14920
rect 11942 14864 12530 14920
rect 12586 14864 12591 14920
rect 11881 14862 12591 14864
rect 11881 14859 11947 14862
rect 12525 14859 12591 14862
rect 16941 14922 17007 14925
rect 20713 14922 20779 14925
rect 24853 14922 24919 14925
rect 16941 14920 20779 14922
rect 16941 14864 16946 14920
rect 17002 14864 20718 14920
rect 20774 14864 20779 14920
rect 16941 14862 20779 14864
rect 16941 14859 17007 14862
rect 20713 14859 20779 14862
rect 20854 14920 24919 14922
rect 20854 14864 24858 14920
rect 24914 14864 24919 14920
rect 20854 14862 24919 14864
rect 9765 14786 9831 14789
rect 11513 14786 11579 14789
rect 9765 14784 11579 14786
rect 9765 14728 9770 14784
rect 9826 14728 11518 14784
rect 11574 14728 11579 14784
rect 9765 14726 11579 14728
rect 9765 14723 9831 14726
rect 11513 14723 11579 14726
rect 18638 14724 18644 14788
rect 18708 14786 18714 14788
rect 19885 14786 19951 14789
rect 20854 14786 20914 14862
rect 24853 14859 24919 14862
rect 18708 14784 20914 14786
rect 18708 14728 19890 14784
rect 19946 14728 20914 14784
rect 18708 14726 20914 14728
rect 24209 14786 24275 14789
rect 27153 14786 27219 14789
rect 24209 14784 27219 14786
rect 24209 14728 24214 14784
rect 24270 14728 27158 14784
rect 27214 14728 27219 14784
rect 24209 14726 27219 14728
rect 18708 14724 18714 14726
rect 19885 14723 19951 14726
rect 24209 14723 24275 14726
rect 27153 14723 27219 14726
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 15942 14720 16258 14721
rect 15942 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16258 14720
rect 15942 14655 16258 14656
rect 23716 14720 24032 14721
rect 23716 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24032 14720
rect 23716 14655 24032 14656
rect 31490 14720 31806 14721
rect 31490 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31806 14720
rect 31490 14655 31806 14656
rect 18270 14588 18276 14652
rect 18340 14650 18346 14652
rect 19057 14650 19123 14653
rect 18340 14648 19123 14650
rect 18340 14592 19062 14648
rect 19118 14592 19123 14648
rect 18340 14590 19123 14592
rect 18340 14588 18346 14590
rect 19057 14587 19123 14590
rect 19517 14650 19583 14653
rect 19517 14648 23306 14650
rect 19517 14592 19522 14648
rect 19578 14592 23306 14648
rect 19517 14590 23306 14592
rect 19517 14587 19583 14590
rect 23246 14517 23306 14590
rect 17217 14514 17283 14517
rect 19517 14514 19583 14517
rect 17217 14512 19583 14514
rect 17217 14456 17222 14512
rect 17278 14456 19522 14512
rect 19578 14456 19583 14512
rect 17217 14454 19583 14456
rect 17217 14451 17283 14454
rect 19517 14451 19583 14454
rect 19701 14514 19767 14517
rect 22737 14514 22803 14517
rect 19701 14512 22803 14514
rect 19701 14456 19706 14512
rect 19762 14456 22742 14512
rect 22798 14456 22803 14512
rect 19701 14454 22803 14456
rect 23246 14514 23355 14517
rect 30097 14514 30163 14517
rect 23246 14512 30163 14514
rect 23246 14456 23294 14512
rect 23350 14456 30102 14512
rect 30158 14456 30163 14512
rect 23246 14454 30163 14456
rect 19701 14451 19767 14454
rect 22737 14451 22803 14454
rect 23289 14451 23355 14454
rect 30097 14451 30163 14454
rect 9949 14378 10015 14381
rect 12709 14378 12775 14381
rect 9949 14376 12775 14378
rect 9949 14320 9954 14376
rect 10010 14320 12714 14376
rect 12770 14320 12775 14376
rect 9949 14318 12775 14320
rect 9949 14315 10015 14318
rect 12709 14315 12775 14318
rect 18413 14378 18479 14381
rect 21817 14378 21883 14381
rect 18413 14376 21883 14378
rect 18413 14320 18418 14376
rect 18474 14320 21822 14376
rect 21878 14320 21883 14376
rect 18413 14318 21883 14320
rect 18413 14315 18479 14318
rect 21817 14315 21883 14318
rect 25221 14378 25287 14381
rect 28441 14378 28507 14381
rect 25221 14376 28507 14378
rect 25221 14320 25226 14376
rect 25282 14320 28446 14376
rect 28502 14320 28507 14376
rect 25221 14318 28507 14320
rect 25221 14315 25287 14318
rect 28441 14315 28507 14318
rect 14089 14242 14155 14245
rect 17769 14242 17835 14245
rect 19701 14242 19767 14245
rect 14089 14240 19767 14242
rect 14089 14184 14094 14240
rect 14150 14184 17774 14240
rect 17830 14184 19706 14240
rect 19762 14184 19767 14240
rect 14089 14182 19767 14184
rect 21820 14242 21880 14315
rect 26417 14242 26483 14245
rect 21820 14240 26483 14242
rect 21820 14184 26422 14240
rect 26478 14184 26483 14240
rect 21820 14182 26483 14184
rect 14089 14179 14155 14182
rect 17769 14179 17835 14182
rect 19701 14179 19767 14182
rect 26417 14179 26483 14182
rect 4281 14176 4597 14177
rect 4281 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4597 14176
rect 4281 14111 4597 14112
rect 12055 14176 12371 14177
rect 12055 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12371 14176
rect 12055 14111 12371 14112
rect 19829 14176 20145 14177
rect 19829 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20145 14176
rect 19829 14111 20145 14112
rect 27603 14176 27919 14177
rect 27603 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27919 14176
rect 27603 14111 27919 14112
rect 17166 14044 17172 14108
rect 17236 14106 17242 14108
rect 17769 14106 17835 14109
rect 22001 14106 22067 14109
rect 17236 14104 17835 14106
rect 17236 14048 17774 14104
rect 17830 14048 17835 14104
rect 17236 14046 17835 14048
rect 17236 14044 17242 14046
rect 17769 14043 17835 14046
rect 21176 14104 22067 14106
rect 21176 14048 22006 14104
rect 22062 14048 22067 14104
rect 21176 14046 22067 14048
rect 8569 13970 8635 13973
rect 8886 13970 8892 13972
rect 8569 13968 8892 13970
rect 8569 13912 8574 13968
rect 8630 13912 8892 13968
rect 8569 13910 8892 13912
rect 8569 13907 8635 13910
rect 8886 13908 8892 13910
rect 8956 13970 8962 13972
rect 10133 13970 10199 13973
rect 8956 13968 10199 13970
rect 8956 13912 10138 13968
rect 10194 13912 10199 13968
rect 8956 13910 10199 13912
rect 8956 13908 8962 13910
rect 10133 13907 10199 13910
rect 11237 13970 11303 13973
rect 18229 13970 18295 13973
rect 11237 13968 18295 13970
rect 11237 13912 11242 13968
rect 11298 13912 18234 13968
rect 18290 13912 18295 13968
rect 11237 13910 18295 13912
rect 11237 13907 11303 13910
rect 18229 13907 18295 13910
rect 7649 13834 7715 13837
rect 9949 13834 10015 13837
rect 10501 13834 10567 13837
rect 7649 13832 9690 13834
rect 7649 13776 7654 13832
rect 7710 13776 9690 13832
rect 7649 13774 9690 13776
rect 7649 13771 7715 13774
rect 9630 13698 9690 13774
rect 9949 13832 10567 13834
rect 9949 13776 9954 13832
rect 10010 13776 10506 13832
rect 10562 13776 10567 13832
rect 9949 13774 10567 13776
rect 9949 13771 10015 13774
rect 10501 13771 10567 13774
rect 10777 13834 10843 13837
rect 11881 13834 11947 13837
rect 10777 13832 11947 13834
rect 10777 13776 10782 13832
rect 10838 13776 11886 13832
rect 11942 13776 11947 13832
rect 10777 13774 11947 13776
rect 10777 13771 10843 13774
rect 11881 13771 11947 13774
rect 16481 13834 16547 13837
rect 21176 13834 21236 14046
rect 22001 14043 22067 14046
rect 23933 14106 23999 14109
rect 26969 14106 27035 14109
rect 23933 14104 27035 14106
rect 23933 14048 23938 14104
rect 23994 14048 26974 14104
rect 27030 14048 27035 14104
rect 23933 14046 27035 14048
rect 23933 14043 23999 14046
rect 26969 14043 27035 14046
rect 22001 13970 22067 13973
rect 26509 13970 26575 13973
rect 22001 13968 26575 13970
rect 22001 13912 22006 13968
rect 22062 13912 26514 13968
rect 26570 13912 26575 13968
rect 22001 13910 26575 13912
rect 22001 13907 22067 13910
rect 26509 13907 26575 13910
rect 16481 13832 21236 13834
rect 16481 13776 16486 13832
rect 16542 13776 21236 13832
rect 16481 13774 21236 13776
rect 22277 13834 22343 13837
rect 24393 13834 24459 13837
rect 22277 13832 24459 13834
rect 22277 13776 22282 13832
rect 22338 13776 24398 13832
rect 24454 13776 24459 13832
rect 22277 13774 24459 13776
rect 16481 13771 16547 13774
rect 22277 13771 22343 13774
rect 24393 13771 24459 13774
rect 25313 13834 25379 13837
rect 28625 13834 28691 13837
rect 25313 13832 28691 13834
rect 25313 13776 25318 13832
rect 25374 13776 28630 13832
rect 28686 13776 28691 13832
rect 25313 13774 28691 13776
rect 25313 13771 25379 13774
rect 28625 13771 28691 13774
rect 9949 13698 10015 13701
rect 9630 13696 10015 13698
rect 9630 13640 9954 13696
rect 10010 13640 10015 13696
rect 9630 13638 10015 13640
rect 9949 13635 10015 13638
rect 11329 13698 11395 13701
rect 11789 13698 11855 13701
rect 17769 13700 17835 13701
rect 11329 13696 11855 13698
rect 11329 13640 11334 13696
rect 11390 13640 11794 13696
rect 11850 13640 11855 13696
rect 11329 13638 11855 13640
rect 11329 13635 11395 13638
rect 11789 13635 11855 13638
rect 17718 13636 17724 13700
rect 17788 13698 17835 13700
rect 17788 13696 22110 13698
rect 17830 13640 22110 13696
rect 17788 13638 22110 13640
rect 17788 13636 17835 13638
rect 17769 13635 17835 13636
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 15942 13632 16258 13633
rect 15942 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16258 13632
rect 15942 13567 16258 13568
rect 9622 13364 9628 13428
rect 9692 13426 9698 13428
rect 19701 13426 19767 13429
rect 9692 13424 19767 13426
rect 9692 13368 19706 13424
rect 19762 13368 19767 13424
rect 9692 13366 19767 13368
rect 22050 13426 22110 13638
rect 23716 13632 24032 13633
rect 23716 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24032 13632
rect 23716 13567 24032 13568
rect 31490 13632 31806 13633
rect 31490 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31806 13632
rect 31490 13567 31806 13568
rect 22553 13426 22619 13429
rect 27429 13426 27495 13429
rect 22050 13424 27495 13426
rect 22050 13368 22558 13424
rect 22614 13368 27434 13424
rect 27490 13368 27495 13424
rect 22050 13366 27495 13368
rect 9692 13364 9698 13366
rect 19701 13363 19767 13366
rect 22553 13363 22619 13366
rect 27429 13363 27495 13366
rect 8385 13290 8451 13293
rect 10133 13290 10199 13293
rect 8385 13288 10199 13290
rect 8385 13232 8390 13288
rect 8446 13232 10138 13288
rect 10194 13232 10199 13288
rect 8385 13230 10199 13232
rect 8385 13227 8451 13230
rect 10133 13227 10199 13230
rect 11789 13290 11855 13293
rect 14733 13290 14799 13293
rect 11789 13288 14799 13290
rect 11789 13232 11794 13288
rect 11850 13232 14738 13288
rect 14794 13232 14799 13288
rect 11789 13230 14799 13232
rect 11789 13227 11855 13230
rect 14733 13227 14799 13230
rect 16941 13290 17007 13293
rect 24301 13290 24367 13293
rect 27061 13290 27127 13293
rect 16941 13288 27127 13290
rect 16941 13232 16946 13288
rect 17002 13232 24306 13288
rect 24362 13232 27066 13288
rect 27122 13232 27127 13288
rect 16941 13230 27127 13232
rect 16941 13227 17007 13230
rect 24301 13227 24367 13230
rect 27061 13227 27127 13230
rect 8109 13154 8175 13157
rect 10501 13154 10567 13157
rect 8109 13152 10567 13154
rect 8109 13096 8114 13152
rect 8170 13096 10506 13152
rect 10562 13096 10567 13152
rect 8109 13094 10567 13096
rect 8109 13091 8175 13094
rect 10501 13091 10567 13094
rect 17401 13154 17467 13157
rect 17953 13154 18019 13157
rect 17401 13152 18019 13154
rect 17401 13096 17406 13152
rect 17462 13096 17958 13152
rect 18014 13096 18019 13152
rect 17401 13094 18019 13096
rect 17401 13091 17467 13094
rect 17953 13091 18019 13094
rect 20253 13154 20319 13157
rect 22001 13154 22067 13157
rect 20253 13152 22067 13154
rect 20253 13096 20258 13152
rect 20314 13096 22006 13152
rect 22062 13096 22067 13152
rect 20253 13094 22067 13096
rect 20253 13091 20319 13094
rect 22001 13091 22067 13094
rect 4281 13088 4597 13089
rect 4281 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4597 13088
rect 4281 13023 4597 13024
rect 12055 13088 12371 13089
rect 12055 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12371 13088
rect 12055 13023 12371 13024
rect 19829 13088 20145 13089
rect 19829 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20145 13088
rect 19829 13023 20145 13024
rect 27603 13088 27919 13089
rect 27603 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27919 13088
rect 27603 13023 27919 13024
rect 16849 13018 16915 13021
rect 18413 13018 18479 13021
rect 16849 13016 18479 13018
rect 16849 12960 16854 13016
rect 16910 12960 18418 13016
rect 18474 12960 18479 13016
rect 16849 12958 18479 12960
rect 16849 12955 16915 12958
rect 18413 12955 18479 12958
rect 5165 12882 5231 12885
rect 10869 12882 10935 12885
rect 19241 12882 19307 12885
rect 5165 12880 10935 12882
rect 5165 12824 5170 12880
rect 5226 12824 10874 12880
rect 10930 12824 10935 12880
rect 5165 12822 10935 12824
rect 5165 12819 5231 12822
rect 10869 12819 10935 12822
rect 12390 12880 19307 12882
rect 12390 12824 19246 12880
rect 19302 12824 19307 12880
rect 12390 12822 19307 12824
rect 7925 12746 7991 12749
rect 9949 12746 10015 12749
rect 10777 12746 10843 12749
rect 12390 12746 12450 12822
rect 19241 12819 19307 12822
rect 20069 12882 20135 12885
rect 27521 12882 27587 12885
rect 20069 12880 27587 12882
rect 20069 12824 20074 12880
rect 20130 12824 27526 12880
rect 27582 12824 27587 12880
rect 20069 12822 27587 12824
rect 20069 12819 20135 12822
rect 27521 12819 27587 12822
rect 7925 12744 9690 12746
rect 7925 12688 7930 12744
rect 7986 12688 9690 12744
rect 7925 12686 9690 12688
rect 7925 12683 7991 12686
rect 9630 12612 9690 12686
rect 9949 12744 12450 12746
rect 9949 12688 9954 12744
rect 10010 12688 10782 12744
rect 10838 12688 12450 12744
rect 9949 12686 12450 12688
rect 20437 12746 20503 12749
rect 22737 12746 22803 12749
rect 24485 12746 24551 12749
rect 20437 12744 24551 12746
rect 20437 12688 20442 12744
rect 20498 12688 22742 12744
rect 22798 12688 24490 12744
rect 24546 12688 24551 12744
rect 20437 12686 24551 12688
rect 9949 12683 10015 12686
rect 10777 12683 10843 12686
rect 20437 12683 20503 12686
rect 22737 12683 22803 12686
rect 24485 12683 24551 12686
rect 9622 12548 9628 12612
rect 9692 12548 9698 12612
rect 11145 12610 11211 12613
rect 13077 12610 13143 12613
rect 11145 12608 13143 12610
rect 11145 12552 11150 12608
rect 11206 12552 13082 12608
rect 13138 12552 13143 12608
rect 11145 12550 13143 12552
rect 11145 12547 11211 12550
rect 13077 12547 13143 12550
rect 16481 12610 16547 12613
rect 17309 12610 17375 12613
rect 16481 12608 23490 12610
rect 16481 12552 16486 12608
rect 16542 12552 17314 12608
rect 17370 12552 23490 12608
rect 16481 12550 23490 12552
rect 16481 12547 16547 12550
rect 17309 12547 17375 12550
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 15942 12544 16258 12545
rect 15942 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16258 12544
rect 15942 12479 16258 12480
rect 15193 12474 15259 12477
rect 15745 12474 15811 12477
rect 15193 12472 15811 12474
rect 15193 12416 15198 12472
rect 15254 12416 15750 12472
rect 15806 12416 15811 12472
rect 15193 12414 15811 12416
rect 15193 12411 15259 12414
rect 15745 12411 15811 12414
rect 5349 12338 5415 12341
rect 10685 12338 10751 12341
rect 5349 12336 10751 12338
rect 5349 12280 5354 12336
rect 5410 12280 10690 12336
rect 10746 12280 10751 12336
rect 5349 12278 10751 12280
rect 5349 12275 5415 12278
rect 10685 12275 10751 12278
rect 14457 12338 14523 12341
rect 20161 12338 20227 12341
rect 20805 12338 20871 12341
rect 21725 12338 21791 12341
rect 14457 12336 21791 12338
rect 14457 12280 14462 12336
rect 14518 12280 20166 12336
rect 20222 12280 20810 12336
rect 20866 12280 21730 12336
rect 21786 12280 21791 12336
rect 14457 12278 21791 12280
rect 14457 12275 14523 12278
rect 20161 12275 20227 12278
rect 20805 12275 20871 12278
rect 21725 12275 21791 12278
rect 9121 12202 9187 12205
rect 13629 12202 13695 12205
rect 9121 12200 13695 12202
rect 9121 12144 9126 12200
rect 9182 12144 13634 12200
rect 13690 12144 13695 12200
rect 9121 12142 13695 12144
rect 9121 12139 9187 12142
rect 13629 12139 13695 12142
rect 15745 12202 15811 12205
rect 17953 12202 18019 12205
rect 22645 12202 22711 12205
rect 15745 12200 18019 12202
rect 15745 12144 15750 12200
rect 15806 12144 17958 12200
rect 18014 12144 18019 12200
rect 15745 12142 18019 12144
rect 15745 12139 15811 12142
rect 17953 12139 18019 12142
rect 19290 12200 22711 12202
rect 19290 12144 22650 12200
rect 22706 12144 22711 12200
rect 19290 12142 22711 12144
rect 23430 12202 23490 12550
rect 23716 12544 24032 12545
rect 23716 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24032 12544
rect 23716 12479 24032 12480
rect 31490 12544 31806 12545
rect 31490 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31806 12544
rect 31490 12479 31806 12480
rect 24761 12474 24827 12477
rect 25681 12474 25747 12477
rect 24761 12472 25747 12474
rect 24761 12416 24766 12472
rect 24822 12416 25686 12472
rect 25742 12416 25747 12472
rect 24761 12414 25747 12416
rect 24761 12411 24827 12414
rect 25681 12411 25747 12414
rect 23749 12338 23815 12341
rect 26325 12338 26391 12341
rect 23749 12336 26391 12338
rect 23749 12280 23754 12336
rect 23810 12280 26330 12336
rect 26386 12280 26391 12336
rect 23749 12278 26391 12280
rect 23749 12275 23815 12278
rect 26325 12275 26391 12278
rect 29729 12202 29795 12205
rect 23430 12200 29795 12202
rect 23430 12144 29734 12200
rect 29790 12144 29795 12200
rect 23430 12142 29795 12144
rect 9949 12066 10015 12069
rect 11053 12066 11119 12069
rect 9949 12064 11119 12066
rect 9949 12008 9954 12064
rect 10010 12008 11058 12064
rect 11114 12008 11119 12064
rect 9949 12006 11119 12008
rect 9949 12003 10015 12006
rect 11053 12003 11119 12006
rect 15009 12066 15075 12069
rect 16665 12066 16731 12069
rect 15009 12064 16731 12066
rect 15009 12008 15014 12064
rect 15070 12008 16670 12064
rect 16726 12008 16731 12064
rect 15009 12006 16731 12008
rect 15009 12003 15075 12006
rect 16665 12003 16731 12006
rect 4281 12000 4597 12001
rect 4281 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4597 12000
rect 4281 11935 4597 11936
rect 12055 12000 12371 12001
rect 12055 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12371 12000
rect 12055 11935 12371 11936
rect 15009 11930 15075 11933
rect 18873 11930 18939 11933
rect 19290 11930 19350 12142
rect 22645 12139 22711 12142
rect 29729 12139 29795 12142
rect 21725 12066 21791 12069
rect 23749 12066 23815 12069
rect 21725 12064 23815 12066
rect 21725 12008 21730 12064
rect 21786 12008 23754 12064
rect 23810 12008 23815 12064
rect 21725 12006 23815 12008
rect 21725 12003 21791 12006
rect 23749 12003 23815 12006
rect 19829 12000 20145 12001
rect 19829 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20145 12000
rect 19829 11935 20145 11936
rect 27603 12000 27919 12001
rect 27603 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27919 12000
rect 27603 11935 27919 11936
rect 15009 11928 19350 11930
rect 15009 11872 15014 11928
rect 15070 11872 18878 11928
rect 18934 11872 19350 11928
rect 15009 11870 19350 11872
rect 20345 11930 20411 11933
rect 26601 11930 26667 11933
rect 20345 11928 26667 11930
rect 20345 11872 20350 11928
rect 20406 11872 26606 11928
rect 26662 11872 26667 11928
rect 20345 11870 26667 11872
rect 15009 11867 15075 11870
rect 18873 11867 18939 11870
rect 20345 11867 20411 11870
rect 26601 11867 26667 11870
rect 10041 11794 10107 11797
rect 12065 11794 12131 11797
rect 10041 11792 12131 11794
rect 10041 11736 10046 11792
rect 10102 11736 12070 11792
rect 12126 11736 12131 11792
rect 10041 11734 12131 11736
rect 10041 11731 10107 11734
rect 12065 11731 12131 11734
rect 12985 11794 13051 11797
rect 17125 11794 17191 11797
rect 12985 11792 17191 11794
rect 12985 11736 12990 11792
rect 13046 11736 17130 11792
rect 17186 11736 17191 11792
rect 12985 11734 17191 11736
rect 12985 11731 13051 11734
rect 17125 11731 17191 11734
rect 17585 11794 17651 11797
rect 24853 11794 24919 11797
rect 17585 11792 24919 11794
rect 17585 11736 17590 11792
rect 17646 11736 24858 11792
rect 24914 11736 24919 11792
rect 17585 11734 24919 11736
rect 17585 11731 17651 11734
rect 24853 11731 24919 11734
rect 29913 11794 29979 11797
rect 30046 11794 30052 11796
rect 29913 11792 30052 11794
rect 29913 11736 29918 11792
rect 29974 11736 30052 11792
rect 29913 11734 30052 11736
rect 29913 11731 29979 11734
rect 30046 11732 30052 11734
rect 30116 11732 30122 11796
rect 7097 11658 7163 11661
rect 9029 11658 9095 11661
rect 11697 11658 11763 11661
rect 18965 11658 19031 11661
rect 7097 11656 8632 11658
rect 7097 11600 7102 11656
rect 7158 11600 8632 11656
rect 7097 11598 8632 11600
rect 7097 11595 7163 11598
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 8572 11386 8632 11598
rect 9029 11656 9690 11658
rect 9029 11600 9034 11656
rect 9090 11600 9690 11656
rect 9029 11598 9690 11600
rect 9029 11595 9095 11598
rect 9630 11522 9690 11598
rect 11697 11656 19031 11658
rect 11697 11600 11702 11656
rect 11758 11600 18970 11656
rect 19026 11600 19031 11656
rect 11697 11598 19031 11600
rect 11697 11595 11763 11598
rect 18965 11595 19031 11598
rect 19793 11658 19859 11661
rect 22829 11658 22895 11661
rect 19793 11656 22895 11658
rect 19793 11600 19798 11656
rect 19854 11600 22834 11656
rect 22890 11600 22895 11656
rect 19793 11598 22895 11600
rect 19793 11595 19859 11598
rect 22829 11595 22895 11598
rect 12433 11522 12499 11525
rect 9630 11520 12499 11522
rect 9630 11464 12438 11520
rect 12494 11464 12499 11520
rect 9630 11462 12499 11464
rect 12433 11459 12499 11462
rect 13721 11522 13787 11525
rect 15745 11522 15811 11525
rect 21357 11522 21423 11525
rect 13721 11520 15811 11522
rect 13721 11464 13726 11520
rect 13782 11464 15750 11520
rect 15806 11464 15811 11520
rect 13721 11462 15811 11464
rect 13721 11459 13787 11462
rect 15745 11459 15811 11462
rect 20440 11520 21423 11522
rect 20440 11464 21362 11520
rect 21418 11464 21423 11520
rect 20440 11462 21423 11464
rect 15942 11456 16258 11457
rect 15942 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16258 11456
rect 15942 11391 16258 11392
rect 20440 11389 20500 11462
rect 21357 11459 21423 11462
rect 23716 11456 24032 11457
rect 23716 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24032 11456
rect 23716 11391 24032 11392
rect 31490 11456 31806 11457
rect 31490 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31806 11456
rect 31490 11391 31806 11392
rect 12709 11386 12775 11389
rect 13721 11386 13787 11389
rect 8572 11384 13787 11386
rect 8572 11328 12714 11384
rect 12770 11328 13726 11384
rect 13782 11328 13787 11384
rect 8572 11326 13787 11328
rect 12709 11323 12775 11326
rect 13721 11323 13787 11326
rect 16389 11386 16455 11389
rect 20437 11386 20503 11389
rect 16389 11384 20503 11386
rect 16389 11328 16394 11384
rect 16450 11328 20442 11384
rect 20498 11328 20503 11384
rect 16389 11326 20503 11328
rect 16389 11323 16455 11326
rect 20437 11323 20503 11326
rect 11513 11250 11579 11253
rect 15469 11250 15535 11253
rect 11513 11248 15535 11250
rect 11513 11192 11518 11248
rect 11574 11192 15474 11248
rect 15530 11192 15535 11248
rect 11513 11190 15535 11192
rect 11513 11187 11579 11190
rect 15469 11187 15535 11190
rect 15653 11250 15719 11253
rect 21909 11250 21975 11253
rect 15653 11248 21975 11250
rect 15653 11192 15658 11248
rect 15714 11192 21914 11248
rect 21970 11192 21975 11248
rect 15653 11190 21975 11192
rect 15653 11187 15719 11190
rect 21909 11187 21975 11190
rect 5257 11114 5323 11117
rect 9673 11114 9739 11117
rect 5257 11112 9739 11114
rect 5257 11056 5262 11112
rect 5318 11056 9678 11112
rect 9734 11056 9739 11112
rect 5257 11054 9739 11056
rect 5257 11051 5323 11054
rect 9673 11051 9739 11054
rect 11329 11114 11395 11117
rect 14917 11114 14983 11117
rect 11329 11112 14983 11114
rect 11329 11056 11334 11112
rect 11390 11056 14922 11112
rect 14978 11056 14983 11112
rect 11329 11054 14983 11056
rect 11329 11051 11395 11054
rect 14917 11051 14983 11054
rect 16665 11114 16731 11117
rect 18321 11114 18387 11117
rect 16665 11112 18387 11114
rect 16665 11056 16670 11112
rect 16726 11056 18326 11112
rect 18382 11056 18387 11112
rect 16665 11054 18387 11056
rect 16665 11051 16731 11054
rect 18321 11051 18387 11054
rect 19701 11114 19767 11117
rect 24577 11114 24643 11117
rect 19701 11112 24643 11114
rect 19701 11056 19706 11112
rect 19762 11056 24582 11112
rect 24638 11056 24643 11112
rect 19701 11054 24643 11056
rect 19701 11051 19767 11054
rect 24577 11051 24643 11054
rect 8937 10980 9003 10981
rect 8886 10916 8892 10980
rect 8956 10978 9003 10980
rect 10317 10978 10383 10981
rect 8956 10976 10383 10978
rect 8998 10920 10322 10976
rect 10378 10920 10383 10976
rect 8956 10918 10383 10920
rect 8956 10916 9003 10918
rect 8937 10915 9003 10916
rect 10317 10915 10383 10918
rect 10501 10978 10567 10981
rect 11789 10978 11855 10981
rect 10501 10976 11855 10978
rect 10501 10920 10506 10976
rect 10562 10920 11794 10976
rect 11850 10920 11855 10976
rect 10501 10918 11855 10920
rect 10501 10915 10567 10918
rect 11789 10915 11855 10918
rect 13445 10978 13511 10981
rect 18505 10978 18571 10981
rect 13445 10976 18571 10978
rect 13445 10920 13450 10976
rect 13506 10920 18510 10976
rect 18566 10920 18571 10976
rect 13445 10918 18571 10920
rect 13445 10915 13511 10918
rect 18505 10915 18571 10918
rect 4281 10912 4597 10913
rect 4281 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4597 10912
rect 4281 10847 4597 10848
rect 12055 10912 12371 10913
rect 12055 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12371 10912
rect 12055 10847 12371 10848
rect 19829 10912 20145 10913
rect 19829 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20145 10912
rect 19829 10847 20145 10848
rect 27603 10912 27919 10913
rect 27603 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27919 10912
rect 27603 10847 27919 10848
rect 10726 10780 10732 10844
rect 10796 10842 10802 10844
rect 10869 10842 10935 10845
rect 10796 10840 10935 10842
rect 10796 10784 10874 10840
rect 10930 10784 10935 10840
rect 10796 10782 10935 10784
rect 10796 10780 10802 10782
rect 10869 10779 10935 10782
rect 15377 10840 15443 10845
rect 15377 10784 15382 10840
rect 15438 10784 15443 10840
rect 15377 10779 15443 10784
rect 4061 10706 4127 10709
rect 7741 10706 7807 10709
rect 4061 10704 7807 10706
rect 4061 10648 4066 10704
rect 4122 10648 7746 10704
rect 7802 10648 7807 10704
rect 4061 10646 7807 10648
rect 4061 10643 4127 10646
rect 7741 10643 7807 10646
rect 8661 10706 8727 10709
rect 11329 10706 11395 10709
rect 13353 10706 13419 10709
rect 8661 10704 13419 10706
rect 8661 10648 8666 10704
rect 8722 10648 11334 10704
rect 11390 10648 13358 10704
rect 13414 10648 13419 10704
rect 8661 10646 13419 10648
rect 8661 10643 8727 10646
rect 11329 10643 11395 10646
rect 13353 10643 13419 10646
rect 6545 10570 6611 10573
rect 15380 10570 15440 10779
rect 16113 10706 16179 10709
rect 24945 10706 25011 10709
rect 16113 10704 25011 10706
rect 16113 10648 16118 10704
rect 16174 10648 24950 10704
rect 25006 10648 25011 10704
rect 16113 10646 25011 10648
rect 16113 10643 16179 10646
rect 24945 10643 25011 10646
rect 20437 10570 20503 10573
rect 26509 10570 26575 10573
rect 6545 10568 15440 10570
rect 6545 10512 6550 10568
rect 6606 10512 15440 10568
rect 6545 10510 15440 10512
rect 15702 10568 20503 10570
rect 15702 10512 20442 10568
rect 20498 10512 20503 10568
rect 15702 10510 20503 10512
rect 6545 10507 6611 10510
rect 10133 10434 10199 10437
rect 10501 10434 10567 10437
rect 10133 10432 10567 10434
rect 10133 10376 10138 10432
rect 10194 10376 10506 10432
rect 10562 10376 10567 10432
rect 10133 10374 10567 10376
rect 10133 10371 10199 10374
rect 10501 10371 10567 10374
rect 10961 10434 11027 10437
rect 13169 10434 13235 10437
rect 10961 10432 13235 10434
rect 10961 10376 10966 10432
rect 11022 10376 13174 10432
rect 13230 10376 13235 10432
rect 10961 10374 13235 10376
rect 10961 10371 11027 10374
rect 13169 10371 13235 10374
rect 13629 10434 13695 10437
rect 15702 10434 15762 10510
rect 20437 10507 20503 10510
rect 22050 10568 26575 10570
rect 22050 10512 26514 10568
rect 26570 10512 26575 10568
rect 22050 10510 26575 10512
rect 13629 10432 15762 10434
rect 13629 10376 13634 10432
rect 13690 10376 15762 10432
rect 13629 10374 15762 10376
rect 18965 10434 19031 10437
rect 19333 10434 19399 10437
rect 22050 10434 22110 10510
rect 26509 10507 26575 10510
rect 18965 10432 22110 10434
rect 18965 10376 18970 10432
rect 19026 10376 19338 10432
rect 19394 10376 22110 10432
rect 18965 10374 22110 10376
rect 13629 10371 13695 10374
rect 18965 10371 19031 10374
rect 19333 10371 19399 10374
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 15942 10368 16258 10369
rect 15942 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16258 10368
rect 15942 10303 16258 10304
rect 23716 10368 24032 10369
rect 23716 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24032 10368
rect 23716 10303 24032 10304
rect 31490 10368 31806 10369
rect 31490 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31806 10368
rect 31490 10303 31806 10304
rect 12157 10298 12223 10301
rect 14917 10298 14983 10301
rect 12157 10296 14983 10298
rect 12157 10240 12162 10296
rect 12218 10240 14922 10296
rect 14978 10240 14983 10296
rect 12157 10238 14983 10240
rect 12157 10235 12223 10238
rect 14917 10235 14983 10238
rect 8201 10162 8267 10165
rect 13537 10162 13603 10165
rect 8201 10160 13603 10162
rect 8201 10104 8206 10160
rect 8262 10104 13542 10160
rect 13598 10104 13603 10160
rect 8201 10102 13603 10104
rect 8201 10099 8267 10102
rect 13537 10099 13603 10102
rect 18873 10162 18939 10165
rect 27613 10162 27679 10165
rect 18873 10160 27679 10162
rect 18873 10104 18878 10160
rect 18934 10104 27618 10160
rect 27674 10104 27679 10160
rect 18873 10102 27679 10104
rect 18873 10099 18939 10102
rect 27613 10099 27679 10102
rect 6913 10026 6979 10029
rect 7046 10026 7052 10028
rect 6913 10024 7052 10026
rect 6913 9968 6918 10024
rect 6974 9968 7052 10024
rect 6913 9966 7052 9968
rect 6913 9963 6979 9966
rect 7046 9964 7052 9966
rect 7116 9964 7122 10028
rect 8293 10026 8359 10029
rect 12157 10026 12223 10029
rect 8293 10024 12223 10026
rect 8293 9968 8298 10024
rect 8354 9968 12162 10024
rect 12218 9968 12223 10024
rect 8293 9966 12223 9968
rect 8293 9963 8359 9966
rect 12157 9963 12223 9966
rect 12341 10026 12407 10029
rect 14733 10026 14799 10029
rect 20897 10026 20963 10029
rect 12341 10024 14799 10026
rect 12341 9968 12346 10024
rect 12402 9968 14738 10024
rect 14794 9968 14799 10024
rect 12341 9966 14799 9968
rect 12341 9963 12407 9966
rect 14733 9963 14799 9966
rect 19566 10024 20963 10026
rect 19566 9968 20902 10024
rect 20958 9968 20963 10024
rect 19566 9966 20963 9968
rect 10869 9890 10935 9893
rect 11881 9890 11947 9893
rect 10869 9888 11947 9890
rect 10869 9832 10874 9888
rect 10930 9832 11886 9888
rect 11942 9832 11947 9888
rect 10869 9830 11947 9832
rect 10869 9827 10935 9830
rect 11881 9827 11947 9830
rect 12801 9890 12867 9893
rect 19566 9890 19626 9966
rect 20897 9963 20963 9966
rect 23657 10026 23723 10029
rect 24209 10026 24275 10029
rect 27102 10026 27108 10028
rect 23657 10024 27108 10026
rect 23657 9968 23662 10024
rect 23718 9968 24214 10024
rect 24270 9968 27108 10024
rect 23657 9966 27108 9968
rect 23657 9963 23723 9966
rect 24209 9963 24275 9966
rect 27102 9964 27108 9966
rect 27172 9964 27178 10028
rect 12801 9888 19626 9890
rect 12801 9832 12806 9888
rect 12862 9832 19626 9888
rect 12801 9830 19626 9832
rect 21173 9890 21239 9893
rect 24393 9890 24459 9893
rect 25589 9890 25655 9893
rect 26049 9890 26115 9893
rect 21173 9888 26115 9890
rect 21173 9832 21178 9888
rect 21234 9832 24398 9888
rect 24454 9832 25594 9888
rect 25650 9832 26054 9888
rect 26110 9832 26115 9888
rect 21173 9830 26115 9832
rect 12801 9827 12867 9830
rect 21173 9827 21239 9830
rect 24393 9827 24459 9830
rect 25589 9827 25655 9830
rect 26049 9827 26115 9830
rect 4281 9824 4597 9825
rect 4281 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4597 9824
rect 4281 9759 4597 9760
rect 12055 9824 12371 9825
rect 12055 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12371 9824
rect 12055 9759 12371 9760
rect 19829 9824 20145 9825
rect 19829 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20145 9824
rect 19829 9759 20145 9760
rect 27603 9824 27919 9825
rect 27603 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27919 9824
rect 27603 9759 27919 9760
rect 20302 9694 20914 9754
rect 5165 9618 5231 9621
rect 6177 9618 6243 9621
rect 7373 9618 7439 9621
rect 12249 9618 12315 9621
rect 5165 9616 7439 9618
rect 5165 9560 5170 9616
rect 5226 9560 6182 9616
rect 6238 9560 7378 9616
rect 7434 9560 7439 9616
rect 5165 9558 7439 9560
rect 5165 9555 5231 9558
rect 6177 9555 6243 9558
rect 7373 9555 7439 9558
rect 9630 9616 12315 9618
rect 9630 9560 12254 9616
rect 12310 9560 12315 9616
rect 9630 9558 12315 9560
rect 6085 9482 6151 9485
rect 8845 9482 8911 9485
rect 9630 9482 9690 9558
rect 12249 9555 12315 9558
rect 14549 9618 14615 9621
rect 15837 9618 15903 9621
rect 20302 9618 20362 9694
rect 14549 9616 20362 9618
rect 14549 9560 14554 9616
rect 14610 9560 15842 9616
rect 15898 9560 20362 9616
rect 14549 9558 20362 9560
rect 14549 9555 14615 9558
rect 15837 9555 15903 9558
rect 20478 9556 20484 9620
rect 20548 9618 20554 9620
rect 20621 9618 20687 9621
rect 20548 9616 20687 9618
rect 20548 9560 20626 9616
rect 20682 9560 20687 9616
rect 20548 9558 20687 9560
rect 20854 9618 20914 9694
rect 21357 9618 21423 9621
rect 20854 9616 21423 9618
rect 20854 9560 21362 9616
rect 21418 9560 21423 9616
rect 20854 9558 21423 9560
rect 20548 9556 20554 9558
rect 20621 9555 20687 9558
rect 21357 9555 21423 9558
rect 22829 9618 22895 9621
rect 23105 9618 23171 9621
rect 27797 9618 27863 9621
rect 22829 9616 27863 9618
rect 22829 9560 22834 9616
rect 22890 9560 23110 9616
rect 23166 9560 27802 9616
rect 27858 9560 27863 9616
rect 22829 9558 27863 9560
rect 22829 9555 22895 9558
rect 23105 9555 23171 9558
rect 27797 9555 27863 9558
rect 6085 9480 9690 9482
rect 6085 9424 6090 9480
rect 6146 9424 8850 9480
rect 8906 9424 9690 9480
rect 6085 9422 9690 9424
rect 6085 9419 6151 9422
rect 8845 9419 8911 9422
rect 11830 9420 11836 9484
rect 11900 9482 11906 9484
rect 26233 9482 26299 9485
rect 11900 9480 26299 9482
rect 11900 9424 26238 9480
rect 26294 9424 26299 9480
rect 11900 9422 26299 9424
rect 11900 9420 11906 9422
rect 26233 9419 26299 9422
rect 9622 9284 9628 9348
rect 9692 9346 9698 9348
rect 10133 9346 10199 9349
rect 9692 9344 10199 9346
rect 9692 9288 10138 9344
rect 10194 9288 10199 9344
rect 9692 9286 10199 9288
rect 9692 9284 9698 9286
rect 10133 9283 10199 9286
rect 11053 9346 11119 9349
rect 14181 9346 14247 9349
rect 11053 9344 14247 9346
rect 11053 9288 11058 9344
rect 11114 9288 14186 9344
rect 14242 9288 14247 9344
rect 11053 9286 14247 9288
rect 11053 9283 11119 9286
rect 14181 9283 14247 9286
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 15942 9280 16258 9281
rect 15942 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16258 9280
rect 15942 9215 16258 9216
rect 23716 9280 24032 9281
rect 23716 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24032 9280
rect 23716 9215 24032 9216
rect 31490 9280 31806 9281
rect 31490 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31806 9280
rect 31490 9215 31806 9216
rect 4705 9210 4771 9213
rect 7189 9210 7255 9213
rect 8017 9210 8083 9213
rect 4705 9208 8083 9210
rect 4705 9152 4710 9208
rect 4766 9152 7194 9208
rect 7250 9152 8022 9208
rect 8078 9152 8083 9208
rect 4705 9150 8083 9152
rect 4705 9147 4771 9150
rect 7189 9147 7255 9150
rect 8017 9147 8083 9150
rect 10685 9212 10751 9213
rect 10685 9208 10732 9212
rect 10796 9210 10802 9212
rect 12709 9210 12775 9213
rect 15377 9210 15443 9213
rect 10685 9152 10690 9208
rect 10685 9148 10732 9152
rect 10796 9150 10842 9210
rect 12709 9208 15443 9210
rect 12709 9152 12714 9208
rect 12770 9152 15382 9208
rect 15438 9152 15443 9208
rect 12709 9150 15443 9152
rect 10796 9148 10802 9150
rect 10685 9147 10751 9148
rect 12709 9147 12775 9150
rect 15377 9147 15443 9150
rect 5717 9074 5783 9077
rect 19149 9074 19215 9077
rect 5717 9072 19215 9074
rect 5717 9016 5722 9072
rect 5778 9016 19154 9072
rect 19210 9016 19215 9072
rect 5717 9014 19215 9016
rect 5717 9011 5783 9014
rect 19149 9011 19215 9014
rect 20529 9074 20595 9077
rect 24853 9074 24919 9077
rect 20529 9072 24919 9074
rect 20529 9016 20534 9072
rect 20590 9016 24858 9072
rect 24914 9016 24919 9072
rect 20529 9014 24919 9016
rect 20529 9011 20595 9014
rect 24853 9011 24919 9014
rect 3233 8938 3299 8941
rect 5165 8938 5231 8941
rect 3233 8936 5231 8938
rect 3233 8880 3238 8936
rect 3294 8880 5170 8936
rect 5226 8880 5231 8936
rect 3233 8878 5231 8880
rect 3233 8875 3299 8878
rect 5165 8875 5231 8878
rect 7097 8938 7163 8941
rect 8109 8938 8175 8941
rect 7097 8936 8175 8938
rect 7097 8880 7102 8936
rect 7158 8880 8114 8936
rect 8170 8880 8175 8936
rect 7097 8878 8175 8880
rect 7097 8875 7163 8878
rect 8109 8875 8175 8878
rect 8477 8938 8543 8941
rect 9949 8940 10015 8941
rect 9806 8938 9812 8940
rect 8477 8936 9812 8938
rect 8477 8880 8482 8936
rect 8538 8880 9812 8936
rect 8477 8878 9812 8880
rect 8477 8875 8543 8878
rect 9806 8876 9812 8878
rect 9876 8876 9882 8940
rect 9949 8936 9996 8940
rect 10060 8938 10066 8940
rect 10409 8938 10475 8941
rect 12065 8938 12131 8941
rect 9949 8880 9954 8936
rect 9949 8876 9996 8880
rect 10060 8878 10106 8938
rect 10409 8936 12131 8938
rect 10409 8880 10414 8936
rect 10470 8880 12070 8936
rect 12126 8880 12131 8936
rect 10409 8878 12131 8880
rect 10060 8876 10066 8878
rect 9949 8875 10015 8876
rect 10409 8875 10475 8878
rect 12065 8875 12131 8878
rect 16941 8938 17007 8941
rect 24209 8938 24275 8941
rect 16941 8936 24275 8938
rect 16941 8880 16946 8936
rect 17002 8880 24214 8936
rect 24270 8880 24275 8936
rect 16941 8878 24275 8880
rect 16941 8875 17007 8878
rect 24209 8875 24275 8878
rect 6085 8802 6151 8805
rect 7925 8802 7991 8805
rect 9489 8804 9555 8805
rect 9438 8802 9444 8804
rect 6085 8800 7991 8802
rect 6085 8744 6090 8800
rect 6146 8744 7930 8800
rect 7986 8744 7991 8800
rect 6085 8742 7991 8744
rect 9362 8742 9444 8802
rect 9508 8802 9555 8804
rect 10685 8802 10751 8805
rect 9508 8800 10751 8802
rect 9550 8744 10690 8800
rect 10746 8744 10751 8800
rect 6085 8739 6151 8742
rect 7925 8739 7991 8742
rect 9438 8740 9444 8742
rect 9508 8742 10751 8744
rect 9508 8740 9555 8742
rect 9489 8739 9555 8740
rect 10685 8739 10751 8742
rect 11053 8802 11119 8805
rect 11421 8802 11487 8805
rect 11053 8800 11487 8802
rect 11053 8744 11058 8800
rect 11114 8744 11426 8800
rect 11482 8744 11487 8800
rect 11053 8742 11487 8744
rect 11053 8739 11119 8742
rect 11421 8739 11487 8742
rect 4281 8736 4597 8737
rect 4281 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4597 8736
rect 4281 8671 4597 8672
rect 12055 8736 12371 8737
rect 12055 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12371 8736
rect 12055 8671 12371 8672
rect 19829 8736 20145 8737
rect 19829 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20145 8736
rect 19829 8671 20145 8672
rect 27603 8736 27919 8737
rect 27603 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27919 8736
rect 27603 8671 27919 8672
rect 7925 8666 7991 8669
rect 11053 8666 11119 8669
rect 16389 8666 16455 8669
rect 7925 8664 11119 8666
rect 7925 8608 7930 8664
rect 7986 8608 11058 8664
rect 11114 8608 11119 8664
rect 7925 8606 11119 8608
rect 7925 8603 7991 8606
rect 11053 8603 11119 8606
rect 12436 8664 16455 8666
rect 12436 8608 16394 8664
rect 16450 8608 16455 8664
rect 12436 8606 16455 8608
rect 6729 8530 6795 8533
rect 8385 8530 8451 8533
rect 8845 8530 8911 8533
rect 6729 8528 8911 8530
rect 6729 8472 6734 8528
rect 6790 8472 8390 8528
rect 8446 8472 8850 8528
rect 8906 8472 8911 8528
rect 6729 8470 8911 8472
rect 6729 8467 6795 8470
rect 8385 8467 8451 8470
rect 8845 8467 8911 8470
rect 10685 8530 10751 8533
rect 12436 8530 12496 8606
rect 16389 8603 16455 8606
rect 10685 8528 12496 8530
rect 10685 8472 10690 8528
rect 10746 8472 12496 8528
rect 10685 8470 12496 8472
rect 10685 8467 10751 8470
rect 12750 8468 12756 8532
rect 12820 8530 12826 8532
rect 19149 8530 19215 8533
rect 12820 8528 19215 8530
rect 12820 8472 19154 8528
rect 19210 8472 19215 8528
rect 12820 8470 19215 8472
rect 12820 8468 12826 8470
rect 19149 8467 19215 8470
rect 19793 8530 19859 8533
rect 23197 8530 23263 8533
rect 19793 8528 23263 8530
rect 19793 8472 19798 8528
rect 19854 8472 23202 8528
rect 23258 8472 23263 8528
rect 19793 8470 23263 8472
rect 19793 8467 19859 8470
rect 23197 8467 23263 8470
rect 5625 8394 5691 8397
rect 7281 8394 7347 8397
rect 7414 8394 7420 8396
rect 5625 8392 7420 8394
rect 5625 8336 5630 8392
rect 5686 8336 7286 8392
rect 7342 8336 7420 8392
rect 5625 8334 7420 8336
rect 5625 8331 5691 8334
rect 7281 8331 7347 8334
rect 7414 8332 7420 8334
rect 7484 8332 7490 8396
rect 8385 8394 8451 8397
rect 11237 8394 11303 8397
rect 8385 8392 11303 8394
rect 8385 8336 8390 8392
rect 8446 8336 11242 8392
rect 11298 8336 11303 8392
rect 8385 8334 11303 8336
rect 8385 8331 8451 8334
rect 11237 8331 11303 8334
rect 10174 8258 10180 8260
rect 8894 8198 10180 8258
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 2037 8122 2103 8125
rect 2865 8122 2931 8125
rect 2037 8120 2931 8122
rect 2037 8064 2042 8120
rect 2098 8064 2870 8120
rect 2926 8064 2931 8120
rect 2037 8062 2931 8064
rect 2037 8059 2103 8062
rect 2865 8059 2931 8062
rect 4061 8122 4127 8125
rect 6453 8122 6519 8125
rect 4061 8120 6519 8122
rect 4061 8064 4066 8120
rect 4122 8064 6458 8120
rect 6514 8064 6519 8120
rect 4061 8062 6519 8064
rect 4061 8059 4127 8062
rect 6453 8059 6519 8062
rect 8894 7989 8954 8198
rect 10174 8196 10180 8198
rect 10244 8258 10250 8260
rect 11513 8258 11579 8261
rect 10244 8256 11579 8258
rect 10244 8200 11518 8256
rect 11574 8200 11579 8256
rect 10244 8198 11579 8200
rect 10244 8196 10250 8198
rect 11513 8195 11579 8198
rect 12750 8196 12756 8260
rect 12820 8196 12826 8260
rect 9029 8122 9095 8125
rect 9581 8122 9647 8125
rect 9029 8120 9647 8122
rect 9029 8064 9034 8120
rect 9090 8064 9586 8120
rect 9642 8064 9647 8120
rect 9029 8062 9647 8064
rect 9029 8059 9095 8062
rect 9581 8059 9647 8062
rect 9857 8122 9923 8125
rect 9990 8122 9996 8124
rect 9857 8120 9996 8122
rect 9857 8064 9862 8120
rect 9918 8064 9996 8120
rect 9857 8062 9996 8064
rect 9857 8059 9923 8062
rect 9990 8060 9996 8062
rect 10060 8060 10066 8124
rect 10225 8122 10291 8125
rect 12758 8122 12818 8196
rect 15942 8192 16258 8193
rect 15942 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16258 8192
rect 15942 8127 16258 8128
rect 23716 8192 24032 8193
rect 23716 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24032 8192
rect 23716 8127 24032 8128
rect 31490 8192 31806 8193
rect 31490 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31806 8192
rect 31490 8127 31806 8128
rect 10225 8120 12818 8122
rect 10225 8064 10230 8120
rect 10286 8064 12818 8120
rect 10225 8062 12818 8064
rect 20529 8122 20595 8125
rect 22737 8122 22803 8125
rect 20529 8120 22803 8122
rect 20529 8064 20534 8120
rect 20590 8064 22742 8120
rect 22798 8064 22803 8120
rect 20529 8062 22803 8064
rect 10225 8059 10291 8062
rect 20529 8059 20595 8062
rect 22737 8059 22803 8062
rect 5901 7986 5967 7989
rect 7005 7986 7071 7989
rect 8569 7986 8635 7989
rect 5901 7984 7071 7986
rect 5901 7928 5906 7984
rect 5962 7928 7010 7984
rect 7066 7928 7071 7984
rect 5901 7926 7071 7928
rect 5901 7923 5967 7926
rect 7005 7923 7071 7926
rect 8250 7984 8635 7986
rect 8250 7928 8574 7984
rect 8630 7928 8635 7984
rect 8250 7926 8635 7928
rect 8894 7984 9003 7989
rect 8894 7928 8942 7984
rect 8998 7928 9003 7984
rect 8894 7926 9003 7928
rect 8250 7853 8310 7926
rect 8569 7923 8635 7926
rect 8937 7923 9003 7926
rect 9765 7986 9831 7989
rect 19333 7986 19399 7989
rect 9765 7984 19399 7986
rect 9765 7928 9770 7984
rect 9826 7928 19338 7984
rect 19394 7928 19399 7984
rect 9765 7926 19399 7928
rect 9765 7923 9831 7926
rect 19333 7923 19399 7926
rect 22369 7986 22435 7989
rect 25957 7986 26023 7989
rect 22369 7984 26023 7986
rect 22369 7928 22374 7984
rect 22430 7928 25962 7984
rect 26018 7928 26023 7984
rect 22369 7926 26023 7928
rect 22369 7923 22435 7926
rect 25957 7923 26023 7926
rect 5441 7850 5507 7853
rect 8017 7852 8083 7853
rect 6862 7850 6868 7852
rect 5441 7848 6868 7850
rect 5441 7792 5446 7848
rect 5502 7792 6868 7848
rect 5441 7790 6868 7792
rect 5441 7787 5507 7790
rect 6862 7788 6868 7790
rect 6932 7788 6938 7852
rect 7966 7850 7972 7852
rect 7926 7790 7972 7850
rect 8036 7848 8083 7852
rect 8078 7792 8083 7848
rect 7966 7788 7972 7790
rect 8036 7788 8083 7792
rect 8017 7787 8083 7788
rect 8201 7848 8310 7853
rect 8661 7852 8727 7853
rect 8661 7850 8708 7852
rect 8201 7792 8206 7848
rect 8262 7792 8310 7848
rect 8201 7790 8310 7792
rect 8616 7848 8708 7850
rect 8616 7792 8666 7848
rect 8616 7790 8708 7792
rect 8201 7787 8267 7790
rect 8661 7788 8708 7790
rect 8772 7788 8778 7852
rect 20253 7850 20319 7853
rect 8894 7848 20319 7850
rect 8894 7792 20258 7848
rect 20314 7792 20319 7848
rect 8894 7790 20319 7792
rect 8661 7787 8727 7788
rect 5441 7716 5507 7717
rect 5390 7714 5396 7716
rect 5314 7654 5396 7714
rect 5460 7714 5507 7716
rect 8894 7714 8954 7790
rect 20253 7787 20319 7790
rect 21725 7850 21791 7853
rect 25865 7850 25931 7853
rect 28349 7850 28415 7853
rect 21725 7848 28415 7850
rect 21725 7792 21730 7848
rect 21786 7792 25870 7848
rect 25926 7792 28354 7848
rect 28410 7792 28415 7848
rect 21725 7790 28415 7792
rect 21725 7787 21791 7790
rect 25865 7787 25931 7790
rect 28349 7787 28415 7790
rect 9765 7714 9831 7717
rect 10777 7716 10843 7717
rect 10726 7714 10732 7716
rect 5460 7712 8954 7714
rect 5502 7656 8954 7712
rect 5390 7652 5396 7654
rect 5460 7654 8954 7656
rect 9078 7712 9831 7714
rect 9078 7656 9770 7712
rect 9826 7656 9831 7712
rect 9078 7654 9831 7656
rect 10686 7654 10732 7714
rect 10796 7712 10843 7716
rect 10838 7656 10843 7712
rect 5460 7652 5507 7654
rect 5441 7651 5507 7652
rect 4281 7648 4597 7649
rect 4281 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4597 7648
rect 4281 7583 4597 7584
rect 6310 7516 6316 7580
rect 6380 7578 6386 7580
rect 9078 7578 9138 7654
rect 9765 7651 9831 7654
rect 10726 7652 10732 7654
rect 10796 7652 10843 7656
rect 10777 7651 10843 7652
rect 10961 7714 11027 7717
rect 11830 7714 11836 7716
rect 10961 7712 11836 7714
rect 10961 7656 10966 7712
rect 11022 7656 11836 7712
rect 10961 7654 11836 7656
rect 10961 7651 11027 7654
rect 11830 7652 11836 7654
rect 11900 7652 11906 7716
rect 20713 7714 20779 7717
rect 23381 7714 23447 7717
rect 20713 7712 23447 7714
rect 20713 7656 20718 7712
rect 20774 7656 23386 7712
rect 23442 7656 23447 7712
rect 20713 7654 23447 7656
rect 20713 7651 20779 7654
rect 23381 7651 23447 7654
rect 12055 7648 12371 7649
rect 12055 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12371 7648
rect 12055 7583 12371 7584
rect 19829 7648 20145 7649
rect 19829 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20145 7648
rect 19829 7583 20145 7584
rect 27603 7648 27919 7649
rect 27603 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27919 7648
rect 27603 7583 27919 7584
rect 6380 7518 9138 7578
rect 9949 7578 10015 7581
rect 10542 7578 10548 7580
rect 9949 7576 10548 7578
rect 9949 7520 9954 7576
rect 10010 7520 10548 7576
rect 9949 7518 10548 7520
rect 6380 7516 6386 7518
rect 9949 7515 10015 7518
rect 10542 7516 10548 7518
rect 10612 7578 10618 7580
rect 10612 7518 11898 7578
rect 10612 7516 10618 7518
rect 1025 7442 1091 7445
rect 10685 7442 10751 7445
rect 1025 7440 10751 7442
rect 1025 7384 1030 7440
rect 1086 7384 10690 7440
rect 10746 7384 10751 7440
rect 1025 7382 10751 7384
rect 11838 7442 11898 7518
rect 18229 7576 18295 7581
rect 18229 7520 18234 7576
rect 18290 7520 18295 7576
rect 18229 7515 18295 7520
rect 18232 7442 18292 7515
rect 11838 7382 18292 7442
rect 1025 7379 1091 7382
rect 10685 7379 10751 7382
rect 6729 7306 6795 7309
rect 10225 7306 10291 7309
rect 11605 7306 11671 7309
rect 25221 7306 25287 7309
rect 6729 7304 8770 7306
rect 6729 7248 6734 7304
rect 6790 7248 8770 7304
rect 6729 7246 8770 7248
rect 6729 7243 6795 7246
rect 5441 7170 5507 7173
rect 7281 7170 7347 7173
rect 5441 7168 7347 7170
rect 5441 7112 5446 7168
rect 5502 7112 7286 7168
rect 7342 7112 7347 7168
rect 5441 7110 7347 7112
rect 8710 7170 8770 7246
rect 10225 7304 11671 7306
rect 10225 7248 10230 7304
rect 10286 7248 11610 7304
rect 11666 7248 11671 7304
rect 10225 7246 11671 7248
rect 10225 7243 10291 7246
rect 11605 7243 11671 7246
rect 12390 7304 25287 7306
rect 12390 7248 25226 7304
rect 25282 7248 25287 7304
rect 12390 7246 25287 7248
rect 12390 7170 12450 7246
rect 25221 7243 25287 7246
rect 8710 7110 12450 7170
rect 20161 7170 20227 7173
rect 20437 7170 20503 7173
rect 20161 7168 20503 7170
rect 20161 7112 20166 7168
rect 20222 7112 20442 7168
rect 20498 7112 20503 7168
rect 20161 7110 20503 7112
rect 5441 7107 5507 7110
rect 7281 7107 7347 7110
rect 20161 7107 20227 7110
rect 20437 7107 20503 7110
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 15942 7104 16258 7105
rect 15942 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16258 7104
rect 15942 7039 16258 7040
rect 23716 7104 24032 7105
rect 23716 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24032 7104
rect 23716 7039 24032 7040
rect 31490 7104 31806 7105
rect 31490 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31806 7104
rect 31490 7039 31806 7040
rect 3877 7034 3943 7037
rect 8753 7034 8819 7037
rect 9438 7034 9444 7036
rect 3877 7032 5642 7034
rect 3877 6976 3882 7032
rect 3938 6976 5642 7032
rect 3877 6974 5642 6976
rect 3877 6971 3943 6974
rect 1761 6898 1827 6901
rect 5441 6898 5507 6901
rect 1761 6896 5507 6898
rect 1761 6840 1766 6896
rect 1822 6840 5446 6896
rect 5502 6840 5507 6896
rect 1761 6838 5507 6840
rect 5582 6898 5642 6974
rect 8753 7032 9444 7034
rect 8753 6976 8758 7032
rect 8814 6976 9444 7032
rect 8753 6974 9444 6976
rect 8753 6971 8819 6974
rect 9438 6972 9444 6974
rect 9508 6972 9514 7036
rect 10910 6972 10916 7036
rect 10980 7034 10986 7036
rect 20529 7034 20595 7037
rect 10980 6974 15762 7034
rect 10980 6972 10986 6974
rect 10409 6898 10475 6901
rect 5582 6896 10475 6898
rect 5582 6840 10414 6896
rect 10470 6840 10475 6896
rect 5582 6838 10475 6840
rect 1761 6835 1827 6838
rect 5441 6835 5507 6838
rect 10409 6835 10475 6838
rect 1945 6762 2011 6765
rect 4521 6762 4587 6765
rect 1945 6760 4587 6762
rect 1945 6704 1950 6760
rect 2006 6704 4526 6760
rect 4582 6704 4587 6760
rect 1945 6702 4587 6704
rect 1945 6699 2011 6702
rect 4521 6699 4587 6702
rect 5441 6762 5507 6765
rect 8201 6762 8267 6765
rect 5441 6760 8267 6762
rect 5441 6704 5446 6760
rect 5502 6704 8206 6760
rect 8262 6704 8267 6760
rect 5441 6702 8267 6704
rect 5441 6699 5507 6702
rect 8201 6699 8267 6702
rect 8477 6762 8543 6765
rect 8702 6762 8708 6764
rect 8477 6760 8708 6762
rect 8477 6704 8482 6760
rect 8538 6704 8708 6760
rect 8477 6702 8708 6704
rect 8477 6699 8543 6702
rect 8702 6700 8708 6702
rect 8772 6700 8778 6764
rect 9765 6762 9831 6765
rect 10918 6762 10978 6972
rect 11789 6898 11855 6901
rect 12801 6898 12867 6901
rect 11789 6896 12867 6898
rect 11789 6840 11794 6896
rect 11850 6840 12806 6896
rect 12862 6840 12867 6896
rect 11789 6838 12867 6840
rect 15702 6898 15762 6974
rect 16438 7032 20595 7034
rect 16438 6976 20534 7032
rect 20590 6976 20595 7032
rect 16438 6974 20595 6976
rect 16438 6898 16498 6974
rect 20529 6971 20595 6974
rect 15702 6838 16498 6898
rect 16573 6898 16639 6901
rect 22645 6898 22711 6901
rect 16573 6896 22711 6898
rect 16573 6840 16578 6896
rect 16634 6840 22650 6896
rect 22706 6840 22711 6896
rect 16573 6838 22711 6840
rect 11789 6835 11855 6838
rect 12801 6835 12867 6838
rect 16573 6835 16639 6838
rect 22645 6835 22711 6838
rect 13629 6762 13695 6765
rect 9765 6760 10978 6762
rect 9765 6704 9770 6760
rect 9826 6704 10978 6760
rect 9765 6702 10978 6704
rect 11286 6760 13695 6762
rect 11286 6704 13634 6760
rect 13690 6704 13695 6760
rect 11286 6702 13695 6704
rect 9765 6699 9831 6702
rect 4981 6626 5047 6629
rect 6310 6626 6316 6628
rect 4981 6624 6316 6626
rect 4981 6568 4986 6624
rect 5042 6568 6316 6624
rect 4981 6566 6316 6568
rect 4981 6563 5047 6566
rect 6310 6564 6316 6566
rect 6380 6564 6386 6628
rect 6637 6626 6703 6629
rect 10317 6626 10383 6629
rect 6637 6624 10383 6626
rect 6637 6568 6642 6624
rect 6698 6568 10322 6624
rect 10378 6568 10383 6624
rect 6637 6566 10383 6568
rect 6637 6563 6703 6566
rect 10317 6563 10383 6566
rect 4281 6560 4597 6561
rect 4281 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4597 6560
rect 4281 6495 4597 6496
rect 11286 6493 11346 6702
rect 13629 6699 13695 6702
rect 14733 6762 14799 6765
rect 22829 6762 22895 6765
rect 14733 6760 22895 6762
rect 14733 6704 14738 6760
rect 14794 6704 22834 6760
rect 22890 6704 22895 6760
rect 14733 6702 22895 6704
rect 14733 6699 14799 6702
rect 22829 6699 22895 6702
rect 24117 6762 24183 6765
rect 25589 6762 25655 6765
rect 24117 6760 25655 6762
rect 24117 6704 24122 6760
rect 24178 6704 25594 6760
rect 25650 6704 25655 6760
rect 24117 6702 25655 6704
rect 24117 6699 24183 6702
rect 25589 6699 25655 6702
rect 12985 6626 13051 6629
rect 14273 6626 14339 6629
rect 16573 6626 16639 6629
rect 12985 6624 16639 6626
rect 12985 6568 12990 6624
rect 13046 6568 14278 6624
rect 14334 6568 16578 6624
rect 16634 6568 16639 6624
rect 12985 6566 16639 6568
rect 12985 6563 13051 6566
rect 14273 6563 14339 6566
rect 16573 6563 16639 6566
rect 21817 6626 21883 6629
rect 25405 6626 25471 6629
rect 21817 6624 25471 6626
rect 21817 6568 21822 6624
rect 21878 6568 25410 6624
rect 25466 6568 25471 6624
rect 21817 6566 25471 6568
rect 21817 6563 21883 6566
rect 25405 6563 25471 6566
rect 12055 6560 12371 6561
rect 12055 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12371 6560
rect 12055 6495 12371 6496
rect 19829 6560 20145 6561
rect 19829 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20145 6560
rect 19829 6495 20145 6496
rect 27603 6560 27919 6561
rect 27603 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27919 6560
rect 27603 6495 27919 6496
rect 5809 6490 5875 6493
rect 11237 6490 11346 6493
rect 5809 6488 11346 6490
rect 5809 6432 5814 6488
rect 5870 6432 11242 6488
rect 11298 6432 11346 6488
rect 5809 6430 11346 6432
rect 12433 6490 12499 6493
rect 16941 6490 17007 6493
rect 12433 6488 17007 6490
rect 12433 6432 12438 6488
rect 12494 6432 16946 6488
rect 17002 6432 17007 6488
rect 12433 6430 17007 6432
rect 5809 6427 5875 6430
rect 11237 6427 11303 6430
rect 12433 6427 12499 6430
rect 16941 6427 17007 6430
rect 22001 6490 22067 6493
rect 25681 6490 25747 6493
rect 26693 6490 26759 6493
rect 22001 6488 26759 6490
rect 22001 6432 22006 6488
rect 22062 6432 25686 6488
rect 25742 6432 26698 6488
rect 26754 6432 26759 6488
rect 22001 6430 26759 6432
rect 22001 6427 22067 6430
rect 25681 6427 25747 6430
rect 26693 6427 26759 6430
rect 7833 6354 7899 6357
rect 13537 6354 13603 6357
rect 7833 6352 13603 6354
rect 7833 6296 7838 6352
rect 7894 6296 13542 6352
rect 13598 6296 13603 6352
rect 7833 6294 13603 6296
rect 7833 6291 7899 6294
rect 13537 6291 13603 6294
rect 24025 6354 24091 6357
rect 25497 6354 25563 6357
rect 24025 6352 25563 6354
rect 24025 6296 24030 6352
rect 24086 6296 25502 6352
rect 25558 6296 25563 6352
rect 24025 6294 25563 6296
rect 24025 6291 24091 6294
rect 25497 6291 25563 6294
rect 3969 6218 4035 6221
rect 10685 6218 10751 6221
rect 3969 6216 10751 6218
rect 3969 6160 3974 6216
rect 4030 6160 10690 6216
rect 10746 6160 10751 6216
rect 3969 6158 10751 6160
rect 3969 6155 4035 6158
rect 10685 6155 10751 6158
rect 24945 6218 25011 6221
rect 27613 6218 27679 6221
rect 24945 6216 27679 6218
rect 24945 6160 24950 6216
rect 25006 6160 27618 6216
rect 27674 6160 27679 6216
rect 24945 6158 27679 6160
rect 24945 6155 25011 6158
rect 27613 6155 27679 6158
rect 7414 6020 7420 6084
rect 7484 6082 7490 6084
rect 7741 6082 7807 6085
rect 7484 6080 7807 6082
rect 7484 6024 7746 6080
rect 7802 6024 7807 6080
rect 7484 6022 7807 6024
rect 7484 6020 7490 6022
rect 7741 6019 7807 6022
rect 9213 6082 9279 6085
rect 9765 6084 9831 6085
rect 9213 6080 9690 6082
rect 9213 6024 9218 6080
rect 9274 6024 9690 6080
rect 9213 6022 9690 6024
rect 9213 6019 9279 6022
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 6913 5946 6979 5949
rect 7046 5946 7052 5948
rect 6913 5944 7052 5946
rect 6913 5888 6918 5944
rect 6974 5888 7052 5944
rect 6913 5886 7052 5888
rect 6913 5883 6979 5886
rect 7046 5884 7052 5886
rect 7116 5884 7122 5948
rect 9630 5946 9690 6022
rect 9765 6080 9812 6084
rect 9876 6082 9882 6084
rect 14457 6082 14523 6085
rect 9876 6080 14523 6082
rect 9765 6024 9770 6080
rect 9876 6024 14462 6080
rect 14518 6024 14523 6080
rect 9765 6020 9812 6024
rect 9876 6022 14523 6024
rect 9876 6020 9882 6022
rect 9765 6019 9831 6020
rect 14457 6019 14523 6022
rect 19241 6082 19307 6085
rect 22461 6082 22527 6085
rect 19241 6080 22527 6082
rect 19241 6024 19246 6080
rect 19302 6024 22466 6080
rect 22522 6024 22527 6080
rect 19241 6022 22527 6024
rect 19241 6019 19307 6022
rect 22461 6019 22527 6022
rect 24393 6082 24459 6085
rect 25681 6082 25747 6085
rect 24393 6080 25747 6082
rect 24393 6024 24398 6080
rect 24454 6024 25686 6080
rect 25742 6024 25747 6080
rect 24393 6022 25747 6024
rect 24393 6019 24459 6022
rect 25681 6019 25747 6022
rect 15942 6016 16258 6017
rect 15942 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16258 6016
rect 15942 5951 16258 5952
rect 23716 6016 24032 6017
rect 23716 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24032 6016
rect 23716 5951 24032 5952
rect 31490 6016 31806 6017
rect 31490 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31806 6016
rect 31490 5951 31806 5952
rect 10317 5946 10383 5949
rect 13445 5946 13511 5949
rect 9630 5886 9828 5946
rect 6085 5810 6151 5813
rect 9581 5810 9647 5813
rect 6085 5808 9647 5810
rect 6085 5752 6090 5808
rect 6146 5752 9586 5808
rect 9642 5752 9647 5808
rect 6085 5750 9647 5752
rect 9768 5810 9828 5886
rect 10317 5944 13511 5946
rect 10317 5888 10322 5944
rect 10378 5888 13450 5944
rect 13506 5888 13511 5944
rect 10317 5886 13511 5888
rect 10317 5883 10383 5886
rect 13445 5883 13511 5886
rect 24209 5946 24275 5949
rect 26233 5946 26299 5949
rect 24209 5944 26299 5946
rect 24209 5888 24214 5944
rect 24270 5888 26238 5944
rect 26294 5888 26299 5944
rect 24209 5886 26299 5888
rect 24209 5883 24275 5886
rect 26233 5883 26299 5886
rect 10777 5810 10843 5813
rect 9768 5808 10843 5810
rect 9768 5752 10782 5808
rect 10838 5752 10843 5808
rect 9768 5750 10843 5752
rect 6085 5747 6151 5750
rect 9581 5747 9647 5750
rect 10777 5747 10843 5750
rect 11605 5810 11671 5813
rect 19333 5810 19399 5813
rect 11605 5808 19399 5810
rect 11605 5752 11610 5808
rect 11666 5752 19338 5808
rect 19394 5752 19399 5808
rect 11605 5750 19399 5752
rect 11605 5747 11671 5750
rect 19333 5747 19399 5750
rect 24853 5810 24919 5813
rect 26417 5810 26483 5813
rect 24853 5808 26483 5810
rect 24853 5752 24858 5808
rect 24914 5752 26422 5808
rect 26478 5752 26483 5808
rect 24853 5750 26483 5752
rect 24853 5747 24919 5750
rect 26417 5747 26483 5750
rect 6862 5612 6868 5676
rect 6932 5674 6938 5676
rect 24301 5674 24367 5677
rect 26509 5674 26575 5677
rect 6932 5614 12634 5674
rect 6932 5612 6938 5614
rect 10317 5538 10383 5541
rect 11329 5538 11395 5541
rect 10317 5536 11395 5538
rect 10317 5480 10322 5536
rect 10378 5480 11334 5536
rect 11390 5480 11395 5536
rect 10317 5478 11395 5480
rect 10317 5475 10383 5478
rect 11329 5475 11395 5478
rect 4281 5472 4597 5473
rect 4281 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4597 5472
rect 4281 5407 4597 5408
rect 12055 5472 12371 5473
rect 12055 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12371 5472
rect 12055 5407 12371 5408
rect 10593 5132 10659 5133
rect 10542 5068 10548 5132
rect 10612 5130 10659 5132
rect 12574 5130 12634 5614
rect 24301 5672 26575 5674
rect 24301 5616 24306 5672
rect 24362 5616 26514 5672
rect 26570 5616 26575 5672
rect 24301 5614 26575 5616
rect 24301 5611 24367 5614
rect 26509 5611 26575 5614
rect 25497 5538 25563 5541
rect 27061 5538 27127 5541
rect 25497 5536 27127 5538
rect 25497 5480 25502 5536
rect 25558 5480 27066 5536
rect 27122 5480 27127 5536
rect 25497 5478 27127 5480
rect 25497 5475 25563 5478
rect 27061 5475 27127 5478
rect 19829 5472 20145 5473
rect 19829 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20145 5472
rect 19829 5407 20145 5408
rect 27603 5472 27919 5473
rect 27603 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27919 5472
rect 27603 5407 27919 5408
rect 16205 5402 16271 5405
rect 18321 5402 18387 5405
rect 16205 5400 18387 5402
rect 16205 5344 16210 5400
rect 16266 5344 18326 5400
rect 18382 5344 18387 5400
rect 16205 5342 18387 5344
rect 16205 5339 16271 5342
rect 18321 5339 18387 5342
rect 13353 5266 13419 5269
rect 21357 5266 21423 5269
rect 13353 5264 21423 5266
rect 13353 5208 13358 5264
rect 13414 5208 21362 5264
rect 21418 5208 21423 5264
rect 13353 5206 21423 5208
rect 13353 5203 13419 5206
rect 21357 5203 21423 5206
rect 25221 5266 25287 5269
rect 27153 5266 27219 5269
rect 25221 5264 27219 5266
rect 25221 5208 25226 5264
rect 25282 5208 27158 5264
rect 27214 5208 27219 5264
rect 25221 5206 27219 5208
rect 25221 5203 25287 5206
rect 27153 5203 27219 5206
rect 12985 5130 13051 5133
rect 15561 5130 15627 5133
rect 10612 5128 10704 5130
rect 10654 5072 10704 5128
rect 10612 5070 10704 5072
rect 12574 5128 15627 5130
rect 12574 5072 12990 5128
rect 13046 5072 15566 5128
rect 15622 5072 15627 5128
rect 12574 5070 15627 5072
rect 10612 5068 10659 5070
rect 10593 5067 10659 5068
rect 12985 5067 13051 5070
rect 15561 5067 15627 5070
rect 15745 5130 15811 5133
rect 18321 5130 18387 5133
rect 15745 5128 18387 5130
rect 15745 5072 15750 5128
rect 15806 5072 18326 5128
rect 18382 5072 18387 5128
rect 15745 5070 18387 5072
rect 15745 5067 15811 5070
rect 18321 5067 18387 5070
rect 22093 5130 22159 5133
rect 23933 5130 23999 5133
rect 25957 5130 26023 5133
rect 22093 5128 26023 5130
rect 22093 5072 22098 5128
rect 22154 5072 23938 5128
rect 23994 5072 25962 5128
rect 26018 5072 26023 5128
rect 22093 5070 26023 5072
rect 22093 5067 22159 5070
rect 23933 5067 23999 5070
rect 25957 5067 26023 5070
rect 10317 4994 10383 4997
rect 12893 4994 12959 4997
rect 10317 4992 12959 4994
rect 10317 4936 10322 4992
rect 10378 4936 12898 4992
rect 12954 4936 12959 4992
rect 10317 4934 12959 4936
rect 10317 4931 10383 4934
rect 12893 4931 12959 4934
rect 14181 4994 14247 4997
rect 15469 4994 15535 4997
rect 14181 4992 15535 4994
rect 14181 4936 14186 4992
rect 14242 4936 15474 4992
rect 15530 4936 15535 4992
rect 14181 4934 15535 4936
rect 14181 4931 14247 4934
rect 15469 4931 15535 4934
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 15942 4928 16258 4929
rect 15942 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16258 4928
rect 15942 4863 16258 4864
rect 23716 4928 24032 4929
rect 23716 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24032 4928
rect 23716 4863 24032 4864
rect 31490 4928 31806 4929
rect 31490 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31806 4928
rect 31490 4863 31806 4864
rect 10409 4858 10475 4861
rect 15745 4858 15811 4861
rect 10409 4856 15811 4858
rect 10409 4800 10414 4856
rect 10470 4800 15750 4856
rect 15806 4800 15811 4856
rect 10409 4798 15811 4800
rect 10409 4795 10475 4798
rect 15745 4795 15811 4798
rect 16573 4858 16639 4861
rect 22369 4858 22435 4861
rect 16573 4856 22435 4858
rect 16573 4800 16578 4856
rect 16634 4800 22374 4856
rect 22430 4800 22435 4856
rect 16573 4798 22435 4800
rect 16573 4795 16639 4798
rect 22369 4795 22435 4798
rect 13905 4722 13971 4725
rect 23473 4722 23539 4725
rect 13905 4720 23539 4722
rect 13905 4664 13910 4720
rect 13966 4664 23478 4720
rect 23534 4664 23539 4720
rect 13905 4662 23539 4664
rect 13905 4659 13971 4662
rect 23473 4659 23539 4662
rect 25773 4722 25839 4725
rect 26877 4722 26943 4725
rect 25773 4720 26943 4722
rect 25773 4664 25778 4720
rect 25834 4664 26882 4720
rect 26938 4664 26943 4720
rect 25773 4662 26943 4664
rect 25773 4659 25839 4662
rect 26877 4659 26943 4662
rect 24761 4586 24827 4589
rect 26877 4586 26943 4589
rect 27613 4586 27679 4589
rect 24761 4584 27679 4586
rect 24761 4528 24766 4584
rect 24822 4528 26882 4584
rect 26938 4528 27618 4584
rect 27674 4528 27679 4584
rect 24761 4526 27679 4528
rect 24761 4523 24827 4526
rect 26877 4523 26943 4526
rect 27613 4523 27679 4526
rect 4281 4384 4597 4385
rect 4281 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4597 4384
rect 4281 4319 4597 4320
rect 12055 4384 12371 4385
rect 12055 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12371 4384
rect 12055 4319 12371 4320
rect 19829 4384 20145 4385
rect 19829 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20145 4384
rect 19829 4319 20145 4320
rect 27603 4384 27919 4385
rect 27603 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27919 4384
rect 27603 4319 27919 4320
rect 20437 4178 20503 4181
rect 24393 4178 24459 4181
rect 20437 4176 24459 4178
rect 20437 4120 20442 4176
rect 20498 4120 24398 4176
rect 24454 4120 24459 4176
rect 20437 4118 24459 4120
rect 20437 4115 20503 4118
rect 24393 4115 24459 4118
rect 21265 4042 21331 4045
rect 21909 4042 21975 4045
rect 21265 4040 21975 4042
rect 21265 3984 21270 4040
rect 21326 3984 21914 4040
rect 21970 3984 21975 4040
rect 21265 3982 21975 3984
rect 21265 3979 21331 3982
rect 21909 3979 21975 3982
rect 23013 4042 23079 4045
rect 23289 4042 23355 4045
rect 25037 4042 25103 4045
rect 23013 4040 25103 4042
rect 23013 3984 23018 4040
rect 23074 3984 23294 4040
rect 23350 3984 25042 4040
rect 25098 3984 25103 4040
rect 23013 3982 25103 3984
rect 23013 3979 23079 3982
rect 23289 3979 23355 3982
rect 25037 3979 25103 3982
rect 25589 4042 25655 4045
rect 27153 4042 27219 4045
rect 25589 4040 27219 4042
rect 25589 3984 25594 4040
rect 25650 3984 27158 4040
rect 27214 3984 27219 4040
rect 25589 3982 27219 3984
rect 25589 3979 25655 3982
rect 27153 3979 27219 3982
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 15942 3840 16258 3841
rect 15942 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16258 3840
rect 15942 3775 16258 3776
rect 23716 3840 24032 3841
rect 23716 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24032 3840
rect 23716 3775 24032 3776
rect 31490 3840 31806 3841
rect 31490 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31806 3840
rect 31490 3775 31806 3776
rect 25129 3770 25195 3773
rect 28257 3770 28323 3773
rect 25086 3768 28323 3770
rect 25086 3712 25134 3768
rect 25190 3712 28262 3768
rect 28318 3712 28323 3768
rect 25086 3710 28323 3712
rect 25086 3707 25195 3710
rect 28257 3707 28323 3710
rect 20989 3634 21055 3637
rect 25086 3634 25146 3707
rect 20989 3632 25146 3634
rect 20989 3576 20994 3632
rect 21050 3576 25146 3632
rect 20989 3574 25146 3576
rect 20989 3571 21055 3574
rect 24025 3498 24091 3501
rect 25221 3498 25287 3501
rect 24025 3496 25287 3498
rect 24025 3440 24030 3496
rect 24086 3440 25226 3496
rect 25282 3440 25287 3496
rect 24025 3438 25287 3440
rect 24025 3435 24091 3438
rect 25221 3435 25287 3438
rect 21449 3362 21515 3365
rect 24853 3362 24919 3365
rect 21449 3360 24919 3362
rect 21449 3304 21454 3360
rect 21510 3304 24858 3360
rect 24914 3304 24919 3360
rect 21449 3302 24919 3304
rect 21449 3299 21515 3302
rect 24853 3299 24919 3302
rect 4281 3296 4597 3297
rect 4281 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4597 3296
rect 4281 3231 4597 3232
rect 12055 3296 12371 3297
rect 12055 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12371 3296
rect 12055 3231 12371 3232
rect 19829 3296 20145 3297
rect 19829 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20145 3296
rect 19829 3231 20145 3232
rect 27603 3296 27919 3297
rect 27603 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27919 3296
rect 27603 3231 27919 3232
rect 21725 3090 21791 3093
rect 24669 3090 24735 3093
rect 28625 3090 28691 3093
rect 21725 3088 28691 3090
rect 21725 3032 21730 3088
rect 21786 3032 24674 3088
rect 24730 3032 28630 3088
rect 28686 3032 28691 3088
rect 21725 3030 28691 3032
rect 21725 3027 21791 3030
rect 24669 3027 24735 3030
rect 28625 3027 28691 3030
rect 14181 2954 14247 2957
rect 20069 2954 20135 2957
rect 14181 2952 20135 2954
rect 14181 2896 14186 2952
rect 14242 2896 20074 2952
rect 20130 2896 20135 2952
rect 14181 2894 20135 2896
rect 14181 2891 14247 2894
rect 20069 2891 20135 2894
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 15942 2752 16258 2753
rect 15942 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16258 2752
rect 15942 2687 16258 2688
rect 23716 2752 24032 2753
rect 23716 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24032 2752
rect 23716 2687 24032 2688
rect 31490 2752 31806 2753
rect 31490 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31806 2752
rect 31490 2687 31806 2688
rect 4281 2208 4597 2209
rect 4281 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4597 2208
rect 4281 2143 4597 2144
rect 12055 2208 12371 2209
rect 12055 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12371 2208
rect 12055 2143 12371 2144
rect 19829 2208 20145 2209
rect 19829 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20145 2208
rect 19829 2143 20145 2144
rect 27603 2208 27919 2209
rect 27603 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27919 2208
rect 27603 2143 27919 2144
rect 8168 1664 8484 1665
rect 8168 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8484 1664
rect 8168 1599 8484 1600
rect 15942 1664 16258 1665
rect 15942 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16258 1664
rect 15942 1599 16258 1600
rect 23716 1664 24032 1665
rect 23716 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24032 1664
rect 23716 1599 24032 1600
rect 31490 1664 31806 1665
rect 31490 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31806 1664
rect 31490 1599 31806 1600
rect 4281 1120 4597 1121
rect 4281 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4597 1120
rect 4281 1055 4597 1056
rect 12055 1120 12371 1121
rect 12055 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12371 1120
rect 12055 1055 12371 1056
rect 19829 1120 20145 1121
rect 19829 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20145 1120
rect 19829 1055 20145 1056
rect 27603 1120 27919 1121
rect 27603 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27919 1120
rect 27603 1055 27919 1056
rect 8168 576 8484 577
rect 8168 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8484 576
rect 8168 511 8484 512
rect 15942 576 16258 577
rect 15942 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16258 576
rect 15942 511 16258 512
rect 23716 576 24032 577
rect 23716 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24032 576
rect 23716 511 24032 512
rect 31490 576 31806 577
rect 31490 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31806 576
rect 31490 511 31806 512
<< via3 >>
rect 14780 22068 14844 22132
rect 4476 21992 4540 21996
rect 4476 21936 4526 21992
rect 4526 21936 4540 21992
rect 4476 21932 4540 21936
rect 9628 21932 9692 21996
rect 16252 21932 16316 21996
rect 25084 21932 25148 21996
rect 28764 21932 28828 21996
rect 6684 21796 6748 21860
rect 7420 21796 7484 21860
rect 12572 21796 12636 21860
rect 24348 21796 24412 21860
rect 25820 21796 25884 21860
rect 28028 21856 28092 21860
rect 28028 21800 28078 21856
rect 28078 21800 28092 21856
rect 28028 21796 28092 21800
rect 29500 21796 29564 21860
rect 30236 21856 30300 21860
rect 30236 21800 30286 21856
rect 30286 21800 30300 21856
rect 30236 21796 30300 21800
rect 4287 21788 4351 21792
rect 4287 21732 4291 21788
rect 4291 21732 4347 21788
rect 4347 21732 4351 21788
rect 4287 21728 4351 21732
rect 4367 21788 4431 21792
rect 4367 21732 4371 21788
rect 4371 21732 4427 21788
rect 4427 21732 4431 21788
rect 4367 21728 4431 21732
rect 4447 21788 4511 21792
rect 4447 21732 4451 21788
rect 4451 21732 4507 21788
rect 4507 21732 4511 21788
rect 4447 21728 4511 21732
rect 4527 21788 4591 21792
rect 4527 21732 4531 21788
rect 4531 21732 4587 21788
rect 4587 21732 4591 21788
rect 4527 21728 4591 21732
rect 12061 21788 12125 21792
rect 12061 21732 12065 21788
rect 12065 21732 12121 21788
rect 12121 21732 12125 21788
rect 12061 21728 12125 21732
rect 12141 21788 12205 21792
rect 12141 21732 12145 21788
rect 12145 21732 12201 21788
rect 12201 21732 12205 21788
rect 12141 21728 12205 21732
rect 12221 21788 12285 21792
rect 12221 21732 12225 21788
rect 12225 21732 12281 21788
rect 12281 21732 12285 21788
rect 12221 21728 12285 21732
rect 12301 21788 12365 21792
rect 12301 21732 12305 21788
rect 12305 21732 12361 21788
rect 12361 21732 12365 21788
rect 12301 21728 12365 21732
rect 19835 21788 19899 21792
rect 19835 21732 19839 21788
rect 19839 21732 19895 21788
rect 19895 21732 19899 21788
rect 19835 21728 19899 21732
rect 19915 21788 19979 21792
rect 19915 21732 19919 21788
rect 19919 21732 19975 21788
rect 19975 21732 19979 21788
rect 19915 21728 19979 21732
rect 19995 21788 20059 21792
rect 19995 21732 19999 21788
rect 19999 21732 20055 21788
rect 20055 21732 20059 21788
rect 19995 21728 20059 21732
rect 20075 21788 20139 21792
rect 20075 21732 20079 21788
rect 20079 21732 20135 21788
rect 20135 21732 20139 21788
rect 20075 21728 20139 21732
rect 27609 21788 27673 21792
rect 27609 21732 27613 21788
rect 27613 21732 27669 21788
rect 27669 21732 27673 21788
rect 27609 21728 27673 21732
rect 27689 21788 27753 21792
rect 27689 21732 27693 21788
rect 27693 21732 27749 21788
rect 27749 21732 27753 21788
rect 27689 21728 27753 21732
rect 27769 21788 27833 21792
rect 27769 21732 27773 21788
rect 27773 21732 27829 21788
rect 27829 21732 27833 21788
rect 27769 21728 27833 21732
rect 27849 21788 27913 21792
rect 27849 21732 27853 21788
rect 27853 21732 27909 21788
rect 27909 21732 27913 21788
rect 27849 21728 27913 21732
rect 13308 21720 13372 21724
rect 13308 21664 13358 21720
rect 13358 21664 13372 21720
rect 13308 21660 13372 21664
rect 26556 21660 26620 21724
rect 3740 21524 3804 21588
rect 14044 21524 14108 21588
rect 17724 21524 17788 21588
rect 27292 21524 27356 21588
rect 15516 21388 15580 21452
rect 796 21252 860 21316
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 15948 21244 16012 21248
rect 15948 21188 15952 21244
rect 15952 21188 16008 21244
rect 16008 21188 16012 21244
rect 15948 21184 16012 21188
rect 16028 21244 16092 21248
rect 16028 21188 16032 21244
rect 16032 21188 16088 21244
rect 16088 21188 16092 21244
rect 16028 21184 16092 21188
rect 16108 21244 16172 21248
rect 16108 21188 16112 21244
rect 16112 21188 16168 21244
rect 16168 21188 16172 21244
rect 16108 21184 16172 21188
rect 16188 21244 16252 21248
rect 16188 21188 16192 21244
rect 16192 21188 16248 21244
rect 16248 21188 16252 21244
rect 16188 21184 16252 21188
rect 23722 21244 23786 21248
rect 23722 21188 23726 21244
rect 23726 21188 23782 21244
rect 23782 21188 23786 21244
rect 23722 21184 23786 21188
rect 23802 21244 23866 21248
rect 23802 21188 23806 21244
rect 23806 21188 23862 21244
rect 23862 21188 23866 21244
rect 23802 21184 23866 21188
rect 23882 21244 23946 21248
rect 23882 21188 23886 21244
rect 23886 21188 23942 21244
rect 23942 21188 23946 21244
rect 23882 21184 23946 21188
rect 23962 21244 24026 21248
rect 23962 21188 23966 21244
rect 23966 21188 24022 21244
rect 24022 21188 24026 21244
rect 23962 21184 24026 21188
rect 31496 21244 31560 21248
rect 31496 21188 31500 21244
rect 31500 21188 31556 21244
rect 31556 21188 31560 21244
rect 31496 21184 31560 21188
rect 31576 21244 31640 21248
rect 31576 21188 31580 21244
rect 31580 21188 31636 21244
rect 31636 21188 31640 21244
rect 31576 21184 31640 21188
rect 31656 21244 31720 21248
rect 31656 21188 31660 21244
rect 31660 21188 31716 21244
rect 31716 21188 31720 21244
rect 31656 21184 31720 21188
rect 31736 21244 31800 21248
rect 31736 21188 31740 21244
rect 31740 21188 31796 21244
rect 31796 21188 31800 21244
rect 31736 21184 31800 21188
rect 1532 21116 1596 21180
rect 3004 21116 3068 21180
rect 5948 21116 6012 21180
rect 10364 21040 10428 21044
rect 10364 20984 10414 21040
rect 10414 20984 10428 21040
rect 10364 20980 10428 20984
rect 12756 20980 12820 21044
rect 19380 20980 19444 21044
rect 2268 20708 2332 20772
rect 6316 20768 6380 20772
rect 6316 20712 6366 20768
rect 6366 20712 6380 20768
rect 6316 20708 6380 20712
rect 10916 20708 10980 20772
rect 30052 20708 30116 20772
rect 4287 20700 4351 20704
rect 4287 20644 4291 20700
rect 4291 20644 4347 20700
rect 4347 20644 4351 20700
rect 4287 20640 4351 20644
rect 4367 20700 4431 20704
rect 4367 20644 4371 20700
rect 4371 20644 4427 20700
rect 4427 20644 4431 20700
rect 4367 20640 4431 20644
rect 4447 20700 4511 20704
rect 4447 20644 4451 20700
rect 4451 20644 4507 20700
rect 4507 20644 4511 20700
rect 4447 20640 4511 20644
rect 4527 20700 4591 20704
rect 4527 20644 4531 20700
rect 4531 20644 4587 20700
rect 4587 20644 4591 20700
rect 4527 20640 4591 20644
rect 12061 20700 12125 20704
rect 12061 20644 12065 20700
rect 12065 20644 12121 20700
rect 12121 20644 12125 20700
rect 12061 20640 12125 20644
rect 12141 20700 12205 20704
rect 12141 20644 12145 20700
rect 12145 20644 12201 20700
rect 12201 20644 12205 20700
rect 12141 20640 12205 20644
rect 12221 20700 12285 20704
rect 12221 20644 12225 20700
rect 12225 20644 12281 20700
rect 12281 20644 12285 20700
rect 12221 20640 12285 20644
rect 12301 20700 12365 20704
rect 12301 20644 12305 20700
rect 12305 20644 12361 20700
rect 12361 20644 12365 20700
rect 12301 20640 12365 20644
rect 19835 20700 19899 20704
rect 19835 20644 19839 20700
rect 19839 20644 19895 20700
rect 19895 20644 19899 20700
rect 19835 20640 19899 20644
rect 19915 20700 19979 20704
rect 19915 20644 19919 20700
rect 19919 20644 19975 20700
rect 19975 20644 19979 20700
rect 19915 20640 19979 20644
rect 19995 20700 20059 20704
rect 19995 20644 19999 20700
rect 19999 20644 20055 20700
rect 20055 20644 20059 20700
rect 19995 20640 20059 20644
rect 20075 20700 20139 20704
rect 20075 20644 20079 20700
rect 20079 20644 20135 20700
rect 20135 20644 20139 20700
rect 20075 20640 20139 20644
rect 27609 20700 27673 20704
rect 27609 20644 27613 20700
rect 27613 20644 27669 20700
rect 27669 20644 27673 20700
rect 27609 20640 27673 20644
rect 27689 20700 27753 20704
rect 27689 20644 27693 20700
rect 27693 20644 27749 20700
rect 27749 20644 27753 20700
rect 27689 20640 27753 20644
rect 27769 20700 27833 20704
rect 27769 20644 27773 20700
rect 27773 20644 27829 20700
rect 27829 20644 27833 20700
rect 27769 20640 27833 20644
rect 27849 20700 27913 20704
rect 27849 20644 27853 20700
rect 27853 20644 27909 20700
rect 27909 20644 27913 20700
rect 27849 20640 27913 20644
rect 7972 20632 8036 20636
rect 7972 20576 7986 20632
rect 7986 20576 8036 20632
rect 7972 20572 8036 20576
rect 9628 20572 9692 20636
rect 11836 20632 11900 20636
rect 11836 20576 11850 20632
rect 11850 20576 11900 20632
rect 11836 20572 11900 20576
rect 16988 20572 17052 20636
rect 17724 20300 17788 20364
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 15948 20156 16012 20160
rect 15948 20100 15952 20156
rect 15952 20100 16008 20156
rect 16008 20100 16012 20156
rect 15948 20096 16012 20100
rect 16028 20156 16092 20160
rect 16028 20100 16032 20156
rect 16032 20100 16088 20156
rect 16088 20100 16092 20156
rect 16028 20096 16092 20100
rect 16108 20156 16172 20160
rect 16108 20100 16112 20156
rect 16112 20100 16168 20156
rect 16168 20100 16172 20156
rect 16108 20096 16172 20100
rect 16188 20156 16252 20160
rect 16188 20100 16192 20156
rect 16192 20100 16248 20156
rect 16248 20100 16252 20156
rect 16188 20096 16252 20100
rect 23722 20156 23786 20160
rect 23722 20100 23726 20156
rect 23726 20100 23782 20156
rect 23782 20100 23786 20156
rect 23722 20096 23786 20100
rect 23802 20156 23866 20160
rect 23802 20100 23806 20156
rect 23806 20100 23862 20156
rect 23862 20100 23866 20156
rect 23802 20096 23866 20100
rect 23882 20156 23946 20160
rect 23882 20100 23886 20156
rect 23886 20100 23942 20156
rect 23942 20100 23946 20156
rect 23882 20096 23946 20100
rect 23962 20156 24026 20160
rect 23962 20100 23966 20156
rect 23966 20100 24022 20156
rect 24022 20100 24026 20156
rect 23962 20096 24026 20100
rect 31496 20156 31560 20160
rect 31496 20100 31500 20156
rect 31500 20100 31556 20156
rect 31556 20100 31560 20156
rect 31496 20096 31560 20100
rect 31576 20156 31640 20160
rect 31576 20100 31580 20156
rect 31580 20100 31636 20156
rect 31636 20100 31640 20156
rect 31576 20096 31640 20100
rect 31656 20156 31720 20160
rect 31656 20100 31660 20156
rect 31660 20100 31716 20156
rect 31716 20100 31720 20156
rect 31656 20096 31720 20100
rect 31736 20156 31800 20160
rect 31736 20100 31740 20156
rect 31740 20100 31796 20156
rect 31796 20100 31800 20156
rect 31736 20096 31800 20100
rect 10180 19680 10244 19684
rect 10180 19624 10194 19680
rect 10194 19624 10244 19680
rect 10180 19620 10244 19624
rect 4287 19612 4351 19616
rect 4287 19556 4291 19612
rect 4291 19556 4347 19612
rect 4347 19556 4351 19612
rect 4287 19552 4351 19556
rect 4367 19612 4431 19616
rect 4367 19556 4371 19612
rect 4371 19556 4427 19612
rect 4427 19556 4431 19612
rect 4367 19552 4431 19556
rect 4447 19612 4511 19616
rect 4447 19556 4451 19612
rect 4451 19556 4507 19612
rect 4507 19556 4511 19612
rect 4447 19552 4511 19556
rect 4527 19612 4591 19616
rect 4527 19556 4531 19612
rect 4531 19556 4587 19612
rect 4587 19556 4591 19612
rect 4527 19552 4591 19556
rect 12061 19612 12125 19616
rect 12061 19556 12065 19612
rect 12065 19556 12121 19612
rect 12121 19556 12125 19612
rect 12061 19552 12125 19556
rect 12141 19612 12205 19616
rect 12141 19556 12145 19612
rect 12145 19556 12201 19612
rect 12201 19556 12205 19612
rect 12141 19552 12205 19556
rect 12221 19612 12285 19616
rect 12221 19556 12225 19612
rect 12225 19556 12281 19612
rect 12281 19556 12285 19612
rect 12221 19552 12285 19556
rect 12301 19612 12365 19616
rect 12301 19556 12305 19612
rect 12305 19556 12361 19612
rect 12361 19556 12365 19612
rect 12301 19552 12365 19556
rect 5396 19348 5460 19412
rect 13492 19348 13556 19412
rect 19835 19612 19899 19616
rect 19835 19556 19839 19612
rect 19839 19556 19895 19612
rect 19895 19556 19899 19612
rect 19835 19552 19899 19556
rect 19915 19612 19979 19616
rect 19915 19556 19919 19612
rect 19919 19556 19975 19612
rect 19975 19556 19979 19612
rect 19915 19552 19979 19556
rect 19995 19612 20059 19616
rect 19995 19556 19999 19612
rect 19999 19556 20055 19612
rect 20055 19556 20059 19612
rect 19995 19552 20059 19556
rect 20075 19612 20139 19616
rect 20075 19556 20079 19612
rect 20079 19556 20135 19612
rect 20135 19556 20139 19612
rect 20075 19552 20139 19556
rect 27609 19612 27673 19616
rect 27609 19556 27613 19612
rect 27613 19556 27669 19612
rect 27669 19556 27673 19612
rect 27609 19552 27673 19556
rect 27689 19612 27753 19616
rect 27689 19556 27693 19612
rect 27693 19556 27749 19612
rect 27749 19556 27753 19612
rect 27689 19552 27753 19556
rect 27769 19612 27833 19616
rect 27769 19556 27773 19612
rect 27773 19556 27829 19612
rect 27829 19556 27833 19612
rect 27769 19552 27833 19556
rect 27849 19612 27913 19616
rect 27849 19556 27853 19612
rect 27853 19556 27909 19612
rect 27909 19556 27913 19612
rect 27849 19552 27913 19556
rect 21404 19544 21468 19548
rect 21404 19488 21454 19544
rect 21454 19488 21468 19544
rect 21404 19484 21468 19488
rect 21956 19544 22020 19548
rect 21956 19488 21970 19544
rect 21970 19488 22020 19544
rect 21956 19484 22020 19488
rect 23428 19544 23492 19548
rect 23428 19488 23478 19544
rect 23478 19488 23492 19544
rect 23428 19484 23492 19488
rect 5212 19212 5276 19276
rect 11100 19212 11164 19276
rect 27108 19348 27172 19412
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 15948 19068 16012 19072
rect 15948 19012 15952 19068
rect 15952 19012 16008 19068
rect 16008 19012 16012 19068
rect 15948 19008 16012 19012
rect 16028 19068 16092 19072
rect 16028 19012 16032 19068
rect 16032 19012 16088 19068
rect 16088 19012 16092 19068
rect 16028 19008 16092 19012
rect 16108 19068 16172 19072
rect 16108 19012 16112 19068
rect 16112 19012 16168 19068
rect 16168 19012 16172 19068
rect 16108 19008 16172 19012
rect 16188 19068 16252 19072
rect 16188 19012 16192 19068
rect 16192 19012 16248 19068
rect 16248 19012 16252 19068
rect 16188 19008 16252 19012
rect 23722 19068 23786 19072
rect 23722 19012 23726 19068
rect 23726 19012 23782 19068
rect 23782 19012 23786 19068
rect 23722 19008 23786 19012
rect 23802 19068 23866 19072
rect 23802 19012 23806 19068
rect 23806 19012 23862 19068
rect 23862 19012 23866 19068
rect 23802 19008 23866 19012
rect 23882 19068 23946 19072
rect 23882 19012 23886 19068
rect 23886 19012 23942 19068
rect 23942 19012 23946 19068
rect 23882 19008 23946 19012
rect 23962 19068 24026 19072
rect 23962 19012 23966 19068
rect 23966 19012 24022 19068
rect 24022 19012 24026 19068
rect 23962 19008 24026 19012
rect 31496 19068 31560 19072
rect 31496 19012 31500 19068
rect 31500 19012 31556 19068
rect 31556 19012 31560 19068
rect 31496 19008 31560 19012
rect 31576 19068 31640 19072
rect 31576 19012 31580 19068
rect 31580 19012 31636 19068
rect 31636 19012 31640 19068
rect 31576 19008 31640 19012
rect 31656 19068 31720 19072
rect 31656 19012 31660 19068
rect 31660 19012 31716 19068
rect 31716 19012 31720 19068
rect 31656 19008 31720 19012
rect 31736 19068 31800 19072
rect 31736 19012 31740 19068
rect 31740 19012 31796 19068
rect 31796 19012 31800 19068
rect 31736 19008 31800 19012
rect 16804 18940 16868 19004
rect 11836 18804 11900 18868
rect 20484 18940 20548 19004
rect 4287 18524 4351 18528
rect 4287 18468 4291 18524
rect 4291 18468 4347 18524
rect 4347 18468 4351 18524
rect 4287 18464 4351 18468
rect 4367 18524 4431 18528
rect 4367 18468 4371 18524
rect 4371 18468 4427 18524
rect 4427 18468 4431 18524
rect 4367 18464 4431 18468
rect 4447 18524 4511 18528
rect 4447 18468 4451 18524
rect 4451 18468 4507 18524
rect 4507 18468 4511 18524
rect 4447 18464 4511 18468
rect 4527 18524 4591 18528
rect 4527 18468 4531 18524
rect 4531 18468 4587 18524
rect 4587 18468 4591 18524
rect 4527 18464 4591 18468
rect 12061 18524 12125 18528
rect 12061 18468 12065 18524
rect 12065 18468 12121 18524
rect 12121 18468 12125 18524
rect 12061 18464 12125 18468
rect 12141 18524 12205 18528
rect 12141 18468 12145 18524
rect 12145 18468 12201 18524
rect 12201 18468 12205 18524
rect 12141 18464 12205 18468
rect 12221 18524 12285 18528
rect 12221 18468 12225 18524
rect 12225 18468 12281 18524
rect 12281 18468 12285 18524
rect 12221 18464 12285 18468
rect 12301 18524 12365 18528
rect 12301 18468 12305 18524
rect 12305 18468 12361 18524
rect 12361 18468 12365 18524
rect 12301 18464 12365 18468
rect 19835 18524 19899 18528
rect 19835 18468 19839 18524
rect 19839 18468 19895 18524
rect 19895 18468 19899 18524
rect 19835 18464 19899 18468
rect 19915 18524 19979 18528
rect 19915 18468 19919 18524
rect 19919 18468 19975 18524
rect 19975 18468 19979 18524
rect 19915 18464 19979 18468
rect 19995 18524 20059 18528
rect 19995 18468 19999 18524
rect 19999 18468 20055 18524
rect 20055 18468 20059 18524
rect 19995 18464 20059 18468
rect 20075 18524 20139 18528
rect 20075 18468 20079 18524
rect 20079 18468 20135 18524
rect 20135 18468 20139 18524
rect 20075 18464 20139 18468
rect 27609 18524 27673 18528
rect 27609 18468 27613 18524
rect 27613 18468 27669 18524
rect 27669 18468 27673 18524
rect 27609 18464 27673 18468
rect 27689 18524 27753 18528
rect 27689 18468 27693 18524
rect 27693 18468 27749 18524
rect 27749 18468 27753 18524
rect 27689 18464 27753 18468
rect 27769 18524 27833 18528
rect 27769 18468 27773 18524
rect 27773 18468 27829 18524
rect 27829 18468 27833 18524
rect 27769 18464 27833 18468
rect 27849 18524 27913 18528
rect 27849 18468 27853 18524
rect 27853 18468 27909 18524
rect 27909 18468 27913 18524
rect 27849 18464 27913 18468
rect 9812 18260 9876 18324
rect 18276 18124 18340 18188
rect 18644 17988 18708 18052
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 15948 17980 16012 17984
rect 15948 17924 15952 17980
rect 15952 17924 16008 17980
rect 16008 17924 16012 17980
rect 15948 17920 16012 17924
rect 16028 17980 16092 17984
rect 16028 17924 16032 17980
rect 16032 17924 16088 17980
rect 16088 17924 16092 17980
rect 16028 17920 16092 17924
rect 16108 17980 16172 17984
rect 16108 17924 16112 17980
rect 16112 17924 16168 17980
rect 16168 17924 16172 17980
rect 16108 17920 16172 17924
rect 16188 17980 16252 17984
rect 16188 17924 16192 17980
rect 16192 17924 16248 17980
rect 16248 17924 16252 17980
rect 16188 17920 16252 17924
rect 23722 17980 23786 17984
rect 23722 17924 23726 17980
rect 23726 17924 23782 17980
rect 23782 17924 23786 17980
rect 23722 17920 23786 17924
rect 23802 17980 23866 17984
rect 23802 17924 23806 17980
rect 23806 17924 23862 17980
rect 23862 17924 23866 17980
rect 23802 17920 23866 17924
rect 23882 17980 23946 17984
rect 23882 17924 23886 17980
rect 23886 17924 23942 17980
rect 23942 17924 23946 17980
rect 23882 17920 23946 17924
rect 23962 17980 24026 17984
rect 23962 17924 23966 17980
rect 23966 17924 24022 17980
rect 24022 17924 24026 17980
rect 23962 17920 24026 17924
rect 31496 17980 31560 17984
rect 31496 17924 31500 17980
rect 31500 17924 31556 17980
rect 31556 17924 31560 17980
rect 31496 17920 31560 17924
rect 31576 17980 31640 17984
rect 31576 17924 31580 17980
rect 31580 17924 31636 17980
rect 31636 17924 31640 17980
rect 31576 17920 31640 17924
rect 31656 17980 31720 17984
rect 31656 17924 31660 17980
rect 31660 17924 31716 17980
rect 31716 17924 31720 17980
rect 31656 17920 31720 17924
rect 31736 17980 31800 17984
rect 31736 17924 31740 17980
rect 31740 17924 31796 17980
rect 31796 17924 31800 17980
rect 31736 17920 31800 17924
rect 4287 17436 4351 17440
rect 4287 17380 4291 17436
rect 4291 17380 4347 17436
rect 4347 17380 4351 17436
rect 4287 17376 4351 17380
rect 4367 17436 4431 17440
rect 4367 17380 4371 17436
rect 4371 17380 4427 17436
rect 4427 17380 4431 17436
rect 4367 17376 4431 17380
rect 4447 17436 4511 17440
rect 4447 17380 4451 17436
rect 4451 17380 4507 17436
rect 4507 17380 4511 17436
rect 4447 17376 4511 17380
rect 4527 17436 4591 17440
rect 4527 17380 4531 17436
rect 4531 17380 4587 17436
rect 4587 17380 4591 17436
rect 4527 17376 4591 17380
rect 12061 17436 12125 17440
rect 12061 17380 12065 17436
rect 12065 17380 12121 17436
rect 12121 17380 12125 17436
rect 12061 17376 12125 17380
rect 12141 17436 12205 17440
rect 12141 17380 12145 17436
rect 12145 17380 12201 17436
rect 12201 17380 12205 17436
rect 12141 17376 12205 17380
rect 12221 17436 12285 17440
rect 12221 17380 12225 17436
rect 12225 17380 12281 17436
rect 12281 17380 12285 17436
rect 12221 17376 12285 17380
rect 12301 17436 12365 17440
rect 12301 17380 12305 17436
rect 12305 17380 12361 17436
rect 12361 17380 12365 17436
rect 12301 17376 12365 17380
rect 19835 17436 19899 17440
rect 19835 17380 19839 17436
rect 19839 17380 19895 17436
rect 19895 17380 19899 17436
rect 19835 17376 19899 17380
rect 19915 17436 19979 17440
rect 19915 17380 19919 17436
rect 19919 17380 19975 17436
rect 19975 17380 19979 17436
rect 19915 17376 19979 17380
rect 19995 17436 20059 17440
rect 19995 17380 19999 17436
rect 19999 17380 20055 17436
rect 20055 17380 20059 17436
rect 19995 17376 20059 17380
rect 20075 17436 20139 17440
rect 20075 17380 20079 17436
rect 20079 17380 20135 17436
rect 20135 17380 20139 17436
rect 20075 17376 20139 17380
rect 27609 17436 27673 17440
rect 27609 17380 27613 17436
rect 27613 17380 27669 17436
rect 27669 17380 27673 17436
rect 27609 17376 27673 17380
rect 27689 17436 27753 17440
rect 27689 17380 27693 17436
rect 27693 17380 27749 17436
rect 27749 17380 27753 17436
rect 27689 17376 27753 17380
rect 27769 17436 27833 17440
rect 27769 17380 27773 17436
rect 27773 17380 27829 17436
rect 27829 17380 27833 17436
rect 27769 17376 27833 17380
rect 27849 17436 27913 17440
rect 27849 17380 27853 17436
rect 27853 17380 27909 17436
rect 27909 17380 27913 17436
rect 27849 17376 27913 17380
rect 17172 17368 17236 17372
rect 17172 17312 17186 17368
rect 17186 17312 17236 17368
rect 17172 17308 17236 17312
rect 10732 17172 10796 17236
rect 19564 17232 19628 17236
rect 19564 17176 19614 17232
rect 19614 17176 19628 17232
rect 19564 17172 19628 17176
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 15948 16892 16012 16896
rect 15948 16836 15952 16892
rect 15952 16836 16008 16892
rect 16008 16836 16012 16892
rect 15948 16832 16012 16836
rect 16028 16892 16092 16896
rect 16028 16836 16032 16892
rect 16032 16836 16088 16892
rect 16088 16836 16092 16892
rect 16028 16832 16092 16836
rect 16108 16892 16172 16896
rect 16108 16836 16112 16892
rect 16112 16836 16168 16892
rect 16168 16836 16172 16892
rect 16108 16832 16172 16836
rect 16188 16892 16252 16896
rect 16188 16836 16192 16892
rect 16192 16836 16248 16892
rect 16248 16836 16252 16892
rect 16188 16832 16252 16836
rect 23722 16892 23786 16896
rect 23722 16836 23726 16892
rect 23726 16836 23782 16892
rect 23782 16836 23786 16892
rect 23722 16832 23786 16836
rect 23802 16892 23866 16896
rect 23802 16836 23806 16892
rect 23806 16836 23862 16892
rect 23862 16836 23866 16892
rect 23802 16832 23866 16836
rect 23882 16892 23946 16896
rect 23882 16836 23886 16892
rect 23886 16836 23942 16892
rect 23942 16836 23946 16892
rect 23882 16832 23946 16836
rect 23962 16892 24026 16896
rect 23962 16836 23966 16892
rect 23966 16836 24022 16892
rect 24022 16836 24026 16892
rect 23962 16832 24026 16836
rect 31496 16892 31560 16896
rect 31496 16836 31500 16892
rect 31500 16836 31556 16892
rect 31556 16836 31560 16892
rect 31496 16832 31560 16836
rect 31576 16892 31640 16896
rect 31576 16836 31580 16892
rect 31580 16836 31636 16892
rect 31636 16836 31640 16892
rect 31576 16832 31640 16836
rect 31656 16892 31720 16896
rect 31656 16836 31660 16892
rect 31660 16836 31716 16892
rect 31716 16836 31720 16892
rect 31656 16832 31720 16836
rect 31736 16892 31800 16896
rect 31736 16836 31740 16892
rect 31740 16836 31796 16892
rect 31796 16836 31800 16892
rect 31736 16832 31800 16836
rect 9628 16764 9692 16828
rect 21404 16492 21468 16556
rect 13492 16356 13556 16420
rect 4287 16348 4351 16352
rect 4287 16292 4291 16348
rect 4291 16292 4347 16348
rect 4347 16292 4351 16348
rect 4287 16288 4351 16292
rect 4367 16348 4431 16352
rect 4367 16292 4371 16348
rect 4371 16292 4427 16348
rect 4427 16292 4431 16348
rect 4367 16288 4431 16292
rect 4447 16348 4511 16352
rect 4447 16292 4451 16348
rect 4451 16292 4507 16348
rect 4507 16292 4511 16348
rect 4447 16288 4511 16292
rect 4527 16348 4591 16352
rect 4527 16292 4531 16348
rect 4531 16292 4587 16348
rect 4587 16292 4591 16348
rect 4527 16288 4591 16292
rect 12061 16348 12125 16352
rect 12061 16292 12065 16348
rect 12065 16292 12121 16348
rect 12121 16292 12125 16348
rect 12061 16288 12125 16292
rect 12141 16348 12205 16352
rect 12141 16292 12145 16348
rect 12145 16292 12201 16348
rect 12201 16292 12205 16348
rect 12141 16288 12205 16292
rect 12221 16348 12285 16352
rect 12221 16292 12225 16348
rect 12225 16292 12281 16348
rect 12281 16292 12285 16348
rect 12221 16288 12285 16292
rect 12301 16348 12365 16352
rect 12301 16292 12305 16348
rect 12305 16292 12361 16348
rect 12361 16292 12365 16348
rect 12301 16288 12365 16292
rect 19835 16348 19899 16352
rect 19835 16292 19839 16348
rect 19839 16292 19895 16348
rect 19895 16292 19899 16348
rect 19835 16288 19899 16292
rect 19915 16348 19979 16352
rect 19915 16292 19919 16348
rect 19919 16292 19975 16348
rect 19975 16292 19979 16348
rect 19915 16288 19979 16292
rect 19995 16348 20059 16352
rect 19995 16292 19999 16348
rect 19999 16292 20055 16348
rect 20055 16292 20059 16348
rect 19995 16288 20059 16292
rect 20075 16348 20139 16352
rect 20075 16292 20079 16348
rect 20079 16292 20135 16348
rect 20135 16292 20139 16348
rect 20075 16288 20139 16292
rect 27609 16348 27673 16352
rect 27609 16292 27613 16348
rect 27613 16292 27669 16348
rect 27669 16292 27673 16348
rect 27609 16288 27673 16292
rect 27689 16348 27753 16352
rect 27689 16292 27693 16348
rect 27693 16292 27749 16348
rect 27749 16292 27753 16348
rect 27689 16288 27753 16292
rect 27769 16348 27833 16352
rect 27769 16292 27773 16348
rect 27773 16292 27829 16348
rect 27829 16292 27833 16348
rect 27769 16288 27833 16292
rect 27849 16348 27913 16352
rect 27849 16292 27853 16348
rect 27853 16292 27909 16348
rect 27909 16292 27913 16348
rect 27849 16288 27913 16292
rect 18828 16220 18892 16284
rect 30972 15948 31036 16012
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 15948 15804 16012 15808
rect 15948 15748 15952 15804
rect 15952 15748 16008 15804
rect 16008 15748 16012 15804
rect 15948 15744 16012 15748
rect 16028 15804 16092 15808
rect 16028 15748 16032 15804
rect 16032 15748 16088 15804
rect 16088 15748 16092 15804
rect 16028 15744 16092 15748
rect 16108 15804 16172 15808
rect 16108 15748 16112 15804
rect 16112 15748 16168 15804
rect 16168 15748 16172 15804
rect 16108 15744 16172 15748
rect 16188 15804 16252 15808
rect 16188 15748 16192 15804
rect 16192 15748 16248 15804
rect 16248 15748 16252 15804
rect 16188 15744 16252 15748
rect 23722 15804 23786 15808
rect 23722 15748 23726 15804
rect 23726 15748 23782 15804
rect 23782 15748 23786 15804
rect 23722 15744 23786 15748
rect 23802 15804 23866 15808
rect 23802 15748 23806 15804
rect 23806 15748 23862 15804
rect 23862 15748 23866 15804
rect 23802 15744 23866 15748
rect 23882 15804 23946 15808
rect 23882 15748 23886 15804
rect 23886 15748 23942 15804
rect 23942 15748 23946 15804
rect 23882 15744 23946 15748
rect 23962 15804 24026 15808
rect 23962 15748 23966 15804
rect 23966 15748 24022 15804
rect 24022 15748 24026 15804
rect 23962 15744 24026 15748
rect 31496 15804 31560 15808
rect 31496 15748 31500 15804
rect 31500 15748 31556 15804
rect 31556 15748 31560 15804
rect 31496 15744 31560 15748
rect 31576 15804 31640 15808
rect 31576 15748 31580 15804
rect 31580 15748 31636 15804
rect 31636 15748 31640 15804
rect 31576 15744 31640 15748
rect 31656 15804 31720 15808
rect 31656 15748 31660 15804
rect 31660 15748 31716 15804
rect 31716 15748 31720 15804
rect 31656 15744 31720 15748
rect 31736 15804 31800 15808
rect 31736 15748 31740 15804
rect 31740 15748 31796 15804
rect 31796 15748 31800 15804
rect 31736 15744 31800 15748
rect 23428 15600 23492 15604
rect 23428 15544 23442 15600
rect 23442 15544 23492 15600
rect 23428 15540 23492 15544
rect 16804 15268 16868 15332
rect 4287 15260 4351 15264
rect 4287 15204 4291 15260
rect 4291 15204 4347 15260
rect 4347 15204 4351 15260
rect 4287 15200 4351 15204
rect 4367 15260 4431 15264
rect 4367 15204 4371 15260
rect 4371 15204 4427 15260
rect 4427 15204 4431 15260
rect 4367 15200 4431 15204
rect 4447 15260 4511 15264
rect 4447 15204 4451 15260
rect 4451 15204 4507 15260
rect 4507 15204 4511 15260
rect 4447 15200 4511 15204
rect 4527 15260 4591 15264
rect 4527 15204 4531 15260
rect 4531 15204 4587 15260
rect 4587 15204 4591 15260
rect 4527 15200 4591 15204
rect 12061 15260 12125 15264
rect 12061 15204 12065 15260
rect 12065 15204 12121 15260
rect 12121 15204 12125 15260
rect 12061 15200 12125 15204
rect 12141 15260 12205 15264
rect 12141 15204 12145 15260
rect 12145 15204 12201 15260
rect 12201 15204 12205 15260
rect 12141 15200 12205 15204
rect 12221 15260 12285 15264
rect 12221 15204 12225 15260
rect 12225 15204 12281 15260
rect 12281 15204 12285 15260
rect 12221 15200 12285 15204
rect 12301 15260 12365 15264
rect 12301 15204 12305 15260
rect 12305 15204 12361 15260
rect 12361 15204 12365 15260
rect 12301 15200 12365 15204
rect 7972 15132 8036 15196
rect 18828 15268 18892 15332
rect 19835 15260 19899 15264
rect 19835 15204 19839 15260
rect 19839 15204 19895 15260
rect 19895 15204 19899 15260
rect 19835 15200 19899 15204
rect 19915 15260 19979 15264
rect 19915 15204 19919 15260
rect 19919 15204 19975 15260
rect 19975 15204 19979 15260
rect 19915 15200 19979 15204
rect 19995 15260 20059 15264
rect 19995 15204 19999 15260
rect 19999 15204 20055 15260
rect 20055 15204 20059 15260
rect 19995 15200 20059 15204
rect 20075 15260 20139 15264
rect 20075 15204 20079 15260
rect 20079 15204 20135 15260
rect 20135 15204 20139 15260
rect 20075 15200 20139 15204
rect 27609 15260 27673 15264
rect 27609 15204 27613 15260
rect 27613 15204 27669 15260
rect 27669 15204 27673 15260
rect 27609 15200 27673 15204
rect 27689 15260 27753 15264
rect 27689 15204 27693 15260
rect 27693 15204 27749 15260
rect 27749 15204 27753 15260
rect 27689 15200 27753 15204
rect 27769 15260 27833 15264
rect 27769 15204 27773 15260
rect 27773 15204 27829 15260
rect 27829 15204 27833 15260
rect 27769 15200 27833 15204
rect 27849 15260 27913 15264
rect 27849 15204 27853 15260
rect 27853 15204 27909 15260
rect 27909 15204 27913 15260
rect 27849 15200 27913 15204
rect 19564 14996 19628 15060
rect 21956 15056 22020 15060
rect 21956 15000 22006 15056
rect 22006 15000 22020 15056
rect 21956 14996 22020 15000
rect 9812 14860 9876 14924
rect 18644 14724 18708 14788
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 15948 14716 16012 14720
rect 15948 14660 15952 14716
rect 15952 14660 16008 14716
rect 16008 14660 16012 14716
rect 15948 14656 16012 14660
rect 16028 14716 16092 14720
rect 16028 14660 16032 14716
rect 16032 14660 16088 14716
rect 16088 14660 16092 14716
rect 16028 14656 16092 14660
rect 16108 14716 16172 14720
rect 16108 14660 16112 14716
rect 16112 14660 16168 14716
rect 16168 14660 16172 14716
rect 16108 14656 16172 14660
rect 16188 14716 16252 14720
rect 16188 14660 16192 14716
rect 16192 14660 16248 14716
rect 16248 14660 16252 14716
rect 16188 14656 16252 14660
rect 23722 14716 23786 14720
rect 23722 14660 23726 14716
rect 23726 14660 23782 14716
rect 23782 14660 23786 14716
rect 23722 14656 23786 14660
rect 23802 14716 23866 14720
rect 23802 14660 23806 14716
rect 23806 14660 23862 14716
rect 23862 14660 23866 14716
rect 23802 14656 23866 14660
rect 23882 14716 23946 14720
rect 23882 14660 23886 14716
rect 23886 14660 23942 14716
rect 23942 14660 23946 14716
rect 23882 14656 23946 14660
rect 23962 14716 24026 14720
rect 23962 14660 23966 14716
rect 23966 14660 24022 14716
rect 24022 14660 24026 14716
rect 23962 14656 24026 14660
rect 31496 14716 31560 14720
rect 31496 14660 31500 14716
rect 31500 14660 31556 14716
rect 31556 14660 31560 14716
rect 31496 14656 31560 14660
rect 31576 14716 31640 14720
rect 31576 14660 31580 14716
rect 31580 14660 31636 14716
rect 31636 14660 31640 14716
rect 31576 14656 31640 14660
rect 31656 14716 31720 14720
rect 31656 14660 31660 14716
rect 31660 14660 31716 14716
rect 31716 14660 31720 14716
rect 31656 14656 31720 14660
rect 31736 14716 31800 14720
rect 31736 14660 31740 14716
rect 31740 14660 31796 14716
rect 31796 14660 31800 14716
rect 31736 14656 31800 14660
rect 18276 14588 18340 14652
rect 4287 14172 4351 14176
rect 4287 14116 4291 14172
rect 4291 14116 4347 14172
rect 4347 14116 4351 14172
rect 4287 14112 4351 14116
rect 4367 14172 4431 14176
rect 4367 14116 4371 14172
rect 4371 14116 4427 14172
rect 4427 14116 4431 14172
rect 4367 14112 4431 14116
rect 4447 14172 4511 14176
rect 4447 14116 4451 14172
rect 4451 14116 4507 14172
rect 4507 14116 4511 14172
rect 4447 14112 4511 14116
rect 4527 14172 4591 14176
rect 4527 14116 4531 14172
rect 4531 14116 4587 14172
rect 4587 14116 4591 14172
rect 4527 14112 4591 14116
rect 12061 14172 12125 14176
rect 12061 14116 12065 14172
rect 12065 14116 12121 14172
rect 12121 14116 12125 14172
rect 12061 14112 12125 14116
rect 12141 14172 12205 14176
rect 12141 14116 12145 14172
rect 12145 14116 12201 14172
rect 12201 14116 12205 14172
rect 12141 14112 12205 14116
rect 12221 14172 12285 14176
rect 12221 14116 12225 14172
rect 12225 14116 12281 14172
rect 12281 14116 12285 14172
rect 12221 14112 12285 14116
rect 12301 14172 12365 14176
rect 12301 14116 12305 14172
rect 12305 14116 12361 14172
rect 12361 14116 12365 14172
rect 12301 14112 12365 14116
rect 19835 14172 19899 14176
rect 19835 14116 19839 14172
rect 19839 14116 19895 14172
rect 19895 14116 19899 14172
rect 19835 14112 19899 14116
rect 19915 14172 19979 14176
rect 19915 14116 19919 14172
rect 19919 14116 19975 14172
rect 19975 14116 19979 14172
rect 19915 14112 19979 14116
rect 19995 14172 20059 14176
rect 19995 14116 19999 14172
rect 19999 14116 20055 14172
rect 20055 14116 20059 14172
rect 19995 14112 20059 14116
rect 20075 14172 20139 14176
rect 20075 14116 20079 14172
rect 20079 14116 20135 14172
rect 20135 14116 20139 14172
rect 20075 14112 20139 14116
rect 27609 14172 27673 14176
rect 27609 14116 27613 14172
rect 27613 14116 27669 14172
rect 27669 14116 27673 14172
rect 27609 14112 27673 14116
rect 27689 14172 27753 14176
rect 27689 14116 27693 14172
rect 27693 14116 27749 14172
rect 27749 14116 27753 14172
rect 27689 14112 27753 14116
rect 27769 14172 27833 14176
rect 27769 14116 27773 14172
rect 27773 14116 27829 14172
rect 27829 14116 27833 14172
rect 27769 14112 27833 14116
rect 27849 14172 27913 14176
rect 27849 14116 27853 14172
rect 27853 14116 27909 14172
rect 27909 14116 27913 14172
rect 27849 14112 27913 14116
rect 17172 14044 17236 14108
rect 8892 13908 8956 13972
rect 17724 13696 17788 13700
rect 17724 13640 17774 13696
rect 17774 13640 17788 13696
rect 17724 13636 17788 13640
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 15948 13628 16012 13632
rect 15948 13572 15952 13628
rect 15952 13572 16008 13628
rect 16008 13572 16012 13628
rect 15948 13568 16012 13572
rect 16028 13628 16092 13632
rect 16028 13572 16032 13628
rect 16032 13572 16088 13628
rect 16088 13572 16092 13628
rect 16028 13568 16092 13572
rect 16108 13628 16172 13632
rect 16108 13572 16112 13628
rect 16112 13572 16168 13628
rect 16168 13572 16172 13628
rect 16108 13568 16172 13572
rect 16188 13628 16252 13632
rect 16188 13572 16192 13628
rect 16192 13572 16248 13628
rect 16248 13572 16252 13628
rect 16188 13568 16252 13572
rect 9628 13364 9692 13428
rect 23722 13628 23786 13632
rect 23722 13572 23726 13628
rect 23726 13572 23782 13628
rect 23782 13572 23786 13628
rect 23722 13568 23786 13572
rect 23802 13628 23866 13632
rect 23802 13572 23806 13628
rect 23806 13572 23862 13628
rect 23862 13572 23866 13628
rect 23802 13568 23866 13572
rect 23882 13628 23946 13632
rect 23882 13572 23886 13628
rect 23886 13572 23942 13628
rect 23942 13572 23946 13628
rect 23882 13568 23946 13572
rect 23962 13628 24026 13632
rect 23962 13572 23966 13628
rect 23966 13572 24022 13628
rect 24022 13572 24026 13628
rect 23962 13568 24026 13572
rect 31496 13628 31560 13632
rect 31496 13572 31500 13628
rect 31500 13572 31556 13628
rect 31556 13572 31560 13628
rect 31496 13568 31560 13572
rect 31576 13628 31640 13632
rect 31576 13572 31580 13628
rect 31580 13572 31636 13628
rect 31636 13572 31640 13628
rect 31576 13568 31640 13572
rect 31656 13628 31720 13632
rect 31656 13572 31660 13628
rect 31660 13572 31716 13628
rect 31716 13572 31720 13628
rect 31656 13568 31720 13572
rect 31736 13628 31800 13632
rect 31736 13572 31740 13628
rect 31740 13572 31796 13628
rect 31796 13572 31800 13628
rect 31736 13568 31800 13572
rect 4287 13084 4351 13088
rect 4287 13028 4291 13084
rect 4291 13028 4347 13084
rect 4347 13028 4351 13084
rect 4287 13024 4351 13028
rect 4367 13084 4431 13088
rect 4367 13028 4371 13084
rect 4371 13028 4427 13084
rect 4427 13028 4431 13084
rect 4367 13024 4431 13028
rect 4447 13084 4511 13088
rect 4447 13028 4451 13084
rect 4451 13028 4507 13084
rect 4507 13028 4511 13084
rect 4447 13024 4511 13028
rect 4527 13084 4591 13088
rect 4527 13028 4531 13084
rect 4531 13028 4587 13084
rect 4587 13028 4591 13084
rect 4527 13024 4591 13028
rect 12061 13084 12125 13088
rect 12061 13028 12065 13084
rect 12065 13028 12121 13084
rect 12121 13028 12125 13084
rect 12061 13024 12125 13028
rect 12141 13084 12205 13088
rect 12141 13028 12145 13084
rect 12145 13028 12201 13084
rect 12201 13028 12205 13084
rect 12141 13024 12205 13028
rect 12221 13084 12285 13088
rect 12221 13028 12225 13084
rect 12225 13028 12281 13084
rect 12281 13028 12285 13084
rect 12221 13024 12285 13028
rect 12301 13084 12365 13088
rect 12301 13028 12305 13084
rect 12305 13028 12361 13084
rect 12361 13028 12365 13084
rect 12301 13024 12365 13028
rect 19835 13084 19899 13088
rect 19835 13028 19839 13084
rect 19839 13028 19895 13084
rect 19895 13028 19899 13084
rect 19835 13024 19899 13028
rect 19915 13084 19979 13088
rect 19915 13028 19919 13084
rect 19919 13028 19975 13084
rect 19975 13028 19979 13084
rect 19915 13024 19979 13028
rect 19995 13084 20059 13088
rect 19995 13028 19999 13084
rect 19999 13028 20055 13084
rect 20055 13028 20059 13084
rect 19995 13024 20059 13028
rect 20075 13084 20139 13088
rect 20075 13028 20079 13084
rect 20079 13028 20135 13084
rect 20135 13028 20139 13084
rect 20075 13024 20139 13028
rect 27609 13084 27673 13088
rect 27609 13028 27613 13084
rect 27613 13028 27669 13084
rect 27669 13028 27673 13084
rect 27609 13024 27673 13028
rect 27689 13084 27753 13088
rect 27689 13028 27693 13084
rect 27693 13028 27749 13084
rect 27749 13028 27753 13084
rect 27689 13024 27753 13028
rect 27769 13084 27833 13088
rect 27769 13028 27773 13084
rect 27773 13028 27829 13084
rect 27829 13028 27833 13084
rect 27769 13024 27833 13028
rect 27849 13084 27913 13088
rect 27849 13028 27853 13084
rect 27853 13028 27909 13084
rect 27909 13028 27913 13084
rect 27849 13024 27913 13028
rect 9628 12548 9692 12612
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 15948 12540 16012 12544
rect 15948 12484 15952 12540
rect 15952 12484 16008 12540
rect 16008 12484 16012 12540
rect 15948 12480 16012 12484
rect 16028 12540 16092 12544
rect 16028 12484 16032 12540
rect 16032 12484 16088 12540
rect 16088 12484 16092 12540
rect 16028 12480 16092 12484
rect 16108 12540 16172 12544
rect 16108 12484 16112 12540
rect 16112 12484 16168 12540
rect 16168 12484 16172 12540
rect 16108 12480 16172 12484
rect 16188 12540 16252 12544
rect 16188 12484 16192 12540
rect 16192 12484 16248 12540
rect 16248 12484 16252 12540
rect 16188 12480 16252 12484
rect 23722 12540 23786 12544
rect 23722 12484 23726 12540
rect 23726 12484 23782 12540
rect 23782 12484 23786 12540
rect 23722 12480 23786 12484
rect 23802 12540 23866 12544
rect 23802 12484 23806 12540
rect 23806 12484 23862 12540
rect 23862 12484 23866 12540
rect 23802 12480 23866 12484
rect 23882 12540 23946 12544
rect 23882 12484 23886 12540
rect 23886 12484 23942 12540
rect 23942 12484 23946 12540
rect 23882 12480 23946 12484
rect 23962 12540 24026 12544
rect 23962 12484 23966 12540
rect 23966 12484 24022 12540
rect 24022 12484 24026 12540
rect 23962 12480 24026 12484
rect 31496 12540 31560 12544
rect 31496 12484 31500 12540
rect 31500 12484 31556 12540
rect 31556 12484 31560 12540
rect 31496 12480 31560 12484
rect 31576 12540 31640 12544
rect 31576 12484 31580 12540
rect 31580 12484 31636 12540
rect 31636 12484 31640 12540
rect 31576 12480 31640 12484
rect 31656 12540 31720 12544
rect 31656 12484 31660 12540
rect 31660 12484 31716 12540
rect 31716 12484 31720 12540
rect 31656 12480 31720 12484
rect 31736 12540 31800 12544
rect 31736 12484 31740 12540
rect 31740 12484 31796 12540
rect 31796 12484 31800 12540
rect 31736 12480 31800 12484
rect 4287 11996 4351 12000
rect 4287 11940 4291 11996
rect 4291 11940 4347 11996
rect 4347 11940 4351 11996
rect 4287 11936 4351 11940
rect 4367 11996 4431 12000
rect 4367 11940 4371 11996
rect 4371 11940 4427 11996
rect 4427 11940 4431 11996
rect 4367 11936 4431 11940
rect 4447 11996 4511 12000
rect 4447 11940 4451 11996
rect 4451 11940 4507 11996
rect 4507 11940 4511 11996
rect 4447 11936 4511 11940
rect 4527 11996 4591 12000
rect 4527 11940 4531 11996
rect 4531 11940 4587 11996
rect 4587 11940 4591 11996
rect 4527 11936 4591 11940
rect 12061 11996 12125 12000
rect 12061 11940 12065 11996
rect 12065 11940 12121 11996
rect 12121 11940 12125 11996
rect 12061 11936 12125 11940
rect 12141 11996 12205 12000
rect 12141 11940 12145 11996
rect 12145 11940 12201 11996
rect 12201 11940 12205 11996
rect 12141 11936 12205 11940
rect 12221 11996 12285 12000
rect 12221 11940 12225 11996
rect 12225 11940 12281 11996
rect 12281 11940 12285 11996
rect 12221 11936 12285 11940
rect 12301 11996 12365 12000
rect 12301 11940 12305 11996
rect 12305 11940 12361 11996
rect 12361 11940 12365 11996
rect 12301 11936 12365 11940
rect 19835 11996 19899 12000
rect 19835 11940 19839 11996
rect 19839 11940 19895 11996
rect 19895 11940 19899 11996
rect 19835 11936 19899 11940
rect 19915 11996 19979 12000
rect 19915 11940 19919 11996
rect 19919 11940 19975 11996
rect 19975 11940 19979 11996
rect 19915 11936 19979 11940
rect 19995 11996 20059 12000
rect 19995 11940 19999 11996
rect 19999 11940 20055 11996
rect 20055 11940 20059 11996
rect 19995 11936 20059 11940
rect 20075 11996 20139 12000
rect 20075 11940 20079 11996
rect 20079 11940 20135 11996
rect 20135 11940 20139 11996
rect 20075 11936 20139 11940
rect 27609 11996 27673 12000
rect 27609 11940 27613 11996
rect 27613 11940 27669 11996
rect 27669 11940 27673 11996
rect 27609 11936 27673 11940
rect 27689 11996 27753 12000
rect 27689 11940 27693 11996
rect 27693 11940 27749 11996
rect 27749 11940 27753 11996
rect 27689 11936 27753 11940
rect 27769 11996 27833 12000
rect 27769 11940 27773 11996
rect 27773 11940 27829 11996
rect 27829 11940 27833 11996
rect 27769 11936 27833 11940
rect 27849 11996 27913 12000
rect 27849 11940 27853 11996
rect 27853 11940 27909 11996
rect 27909 11940 27913 11996
rect 27849 11936 27913 11940
rect 30052 11732 30116 11796
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 15948 11452 16012 11456
rect 15948 11396 15952 11452
rect 15952 11396 16008 11452
rect 16008 11396 16012 11452
rect 15948 11392 16012 11396
rect 16028 11452 16092 11456
rect 16028 11396 16032 11452
rect 16032 11396 16088 11452
rect 16088 11396 16092 11452
rect 16028 11392 16092 11396
rect 16108 11452 16172 11456
rect 16108 11396 16112 11452
rect 16112 11396 16168 11452
rect 16168 11396 16172 11452
rect 16108 11392 16172 11396
rect 16188 11452 16252 11456
rect 16188 11396 16192 11452
rect 16192 11396 16248 11452
rect 16248 11396 16252 11452
rect 16188 11392 16252 11396
rect 23722 11452 23786 11456
rect 23722 11396 23726 11452
rect 23726 11396 23782 11452
rect 23782 11396 23786 11452
rect 23722 11392 23786 11396
rect 23802 11452 23866 11456
rect 23802 11396 23806 11452
rect 23806 11396 23862 11452
rect 23862 11396 23866 11452
rect 23802 11392 23866 11396
rect 23882 11452 23946 11456
rect 23882 11396 23886 11452
rect 23886 11396 23942 11452
rect 23942 11396 23946 11452
rect 23882 11392 23946 11396
rect 23962 11452 24026 11456
rect 23962 11396 23966 11452
rect 23966 11396 24022 11452
rect 24022 11396 24026 11452
rect 23962 11392 24026 11396
rect 31496 11452 31560 11456
rect 31496 11396 31500 11452
rect 31500 11396 31556 11452
rect 31556 11396 31560 11452
rect 31496 11392 31560 11396
rect 31576 11452 31640 11456
rect 31576 11396 31580 11452
rect 31580 11396 31636 11452
rect 31636 11396 31640 11452
rect 31576 11392 31640 11396
rect 31656 11452 31720 11456
rect 31656 11396 31660 11452
rect 31660 11396 31716 11452
rect 31716 11396 31720 11452
rect 31656 11392 31720 11396
rect 31736 11452 31800 11456
rect 31736 11396 31740 11452
rect 31740 11396 31796 11452
rect 31796 11396 31800 11452
rect 31736 11392 31800 11396
rect 8892 10976 8956 10980
rect 8892 10920 8942 10976
rect 8942 10920 8956 10976
rect 8892 10916 8956 10920
rect 4287 10908 4351 10912
rect 4287 10852 4291 10908
rect 4291 10852 4347 10908
rect 4347 10852 4351 10908
rect 4287 10848 4351 10852
rect 4367 10908 4431 10912
rect 4367 10852 4371 10908
rect 4371 10852 4427 10908
rect 4427 10852 4431 10908
rect 4367 10848 4431 10852
rect 4447 10908 4511 10912
rect 4447 10852 4451 10908
rect 4451 10852 4507 10908
rect 4507 10852 4511 10908
rect 4447 10848 4511 10852
rect 4527 10908 4591 10912
rect 4527 10852 4531 10908
rect 4531 10852 4587 10908
rect 4587 10852 4591 10908
rect 4527 10848 4591 10852
rect 12061 10908 12125 10912
rect 12061 10852 12065 10908
rect 12065 10852 12121 10908
rect 12121 10852 12125 10908
rect 12061 10848 12125 10852
rect 12141 10908 12205 10912
rect 12141 10852 12145 10908
rect 12145 10852 12201 10908
rect 12201 10852 12205 10908
rect 12141 10848 12205 10852
rect 12221 10908 12285 10912
rect 12221 10852 12225 10908
rect 12225 10852 12281 10908
rect 12281 10852 12285 10908
rect 12221 10848 12285 10852
rect 12301 10908 12365 10912
rect 12301 10852 12305 10908
rect 12305 10852 12361 10908
rect 12361 10852 12365 10908
rect 12301 10848 12365 10852
rect 19835 10908 19899 10912
rect 19835 10852 19839 10908
rect 19839 10852 19895 10908
rect 19895 10852 19899 10908
rect 19835 10848 19899 10852
rect 19915 10908 19979 10912
rect 19915 10852 19919 10908
rect 19919 10852 19975 10908
rect 19975 10852 19979 10908
rect 19915 10848 19979 10852
rect 19995 10908 20059 10912
rect 19995 10852 19999 10908
rect 19999 10852 20055 10908
rect 20055 10852 20059 10908
rect 19995 10848 20059 10852
rect 20075 10908 20139 10912
rect 20075 10852 20079 10908
rect 20079 10852 20135 10908
rect 20135 10852 20139 10908
rect 20075 10848 20139 10852
rect 27609 10908 27673 10912
rect 27609 10852 27613 10908
rect 27613 10852 27669 10908
rect 27669 10852 27673 10908
rect 27609 10848 27673 10852
rect 27689 10908 27753 10912
rect 27689 10852 27693 10908
rect 27693 10852 27749 10908
rect 27749 10852 27753 10908
rect 27689 10848 27753 10852
rect 27769 10908 27833 10912
rect 27769 10852 27773 10908
rect 27773 10852 27829 10908
rect 27829 10852 27833 10908
rect 27769 10848 27833 10852
rect 27849 10908 27913 10912
rect 27849 10852 27853 10908
rect 27853 10852 27909 10908
rect 27909 10852 27913 10908
rect 27849 10848 27913 10852
rect 10732 10780 10796 10844
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 15948 10364 16012 10368
rect 15948 10308 15952 10364
rect 15952 10308 16008 10364
rect 16008 10308 16012 10364
rect 15948 10304 16012 10308
rect 16028 10364 16092 10368
rect 16028 10308 16032 10364
rect 16032 10308 16088 10364
rect 16088 10308 16092 10364
rect 16028 10304 16092 10308
rect 16108 10364 16172 10368
rect 16108 10308 16112 10364
rect 16112 10308 16168 10364
rect 16168 10308 16172 10364
rect 16108 10304 16172 10308
rect 16188 10364 16252 10368
rect 16188 10308 16192 10364
rect 16192 10308 16248 10364
rect 16248 10308 16252 10364
rect 16188 10304 16252 10308
rect 23722 10364 23786 10368
rect 23722 10308 23726 10364
rect 23726 10308 23782 10364
rect 23782 10308 23786 10364
rect 23722 10304 23786 10308
rect 23802 10364 23866 10368
rect 23802 10308 23806 10364
rect 23806 10308 23862 10364
rect 23862 10308 23866 10364
rect 23802 10304 23866 10308
rect 23882 10364 23946 10368
rect 23882 10308 23886 10364
rect 23886 10308 23942 10364
rect 23942 10308 23946 10364
rect 23882 10304 23946 10308
rect 23962 10364 24026 10368
rect 23962 10308 23966 10364
rect 23966 10308 24022 10364
rect 24022 10308 24026 10364
rect 23962 10304 24026 10308
rect 31496 10364 31560 10368
rect 31496 10308 31500 10364
rect 31500 10308 31556 10364
rect 31556 10308 31560 10364
rect 31496 10304 31560 10308
rect 31576 10364 31640 10368
rect 31576 10308 31580 10364
rect 31580 10308 31636 10364
rect 31636 10308 31640 10364
rect 31576 10304 31640 10308
rect 31656 10364 31720 10368
rect 31656 10308 31660 10364
rect 31660 10308 31716 10364
rect 31716 10308 31720 10364
rect 31656 10304 31720 10308
rect 31736 10364 31800 10368
rect 31736 10308 31740 10364
rect 31740 10308 31796 10364
rect 31796 10308 31800 10364
rect 31736 10304 31800 10308
rect 7052 9964 7116 10028
rect 27108 9964 27172 10028
rect 4287 9820 4351 9824
rect 4287 9764 4291 9820
rect 4291 9764 4347 9820
rect 4347 9764 4351 9820
rect 4287 9760 4351 9764
rect 4367 9820 4431 9824
rect 4367 9764 4371 9820
rect 4371 9764 4427 9820
rect 4427 9764 4431 9820
rect 4367 9760 4431 9764
rect 4447 9820 4511 9824
rect 4447 9764 4451 9820
rect 4451 9764 4507 9820
rect 4507 9764 4511 9820
rect 4447 9760 4511 9764
rect 4527 9820 4591 9824
rect 4527 9764 4531 9820
rect 4531 9764 4587 9820
rect 4587 9764 4591 9820
rect 4527 9760 4591 9764
rect 12061 9820 12125 9824
rect 12061 9764 12065 9820
rect 12065 9764 12121 9820
rect 12121 9764 12125 9820
rect 12061 9760 12125 9764
rect 12141 9820 12205 9824
rect 12141 9764 12145 9820
rect 12145 9764 12201 9820
rect 12201 9764 12205 9820
rect 12141 9760 12205 9764
rect 12221 9820 12285 9824
rect 12221 9764 12225 9820
rect 12225 9764 12281 9820
rect 12281 9764 12285 9820
rect 12221 9760 12285 9764
rect 12301 9820 12365 9824
rect 12301 9764 12305 9820
rect 12305 9764 12361 9820
rect 12361 9764 12365 9820
rect 12301 9760 12365 9764
rect 19835 9820 19899 9824
rect 19835 9764 19839 9820
rect 19839 9764 19895 9820
rect 19895 9764 19899 9820
rect 19835 9760 19899 9764
rect 19915 9820 19979 9824
rect 19915 9764 19919 9820
rect 19919 9764 19975 9820
rect 19975 9764 19979 9820
rect 19915 9760 19979 9764
rect 19995 9820 20059 9824
rect 19995 9764 19999 9820
rect 19999 9764 20055 9820
rect 20055 9764 20059 9820
rect 19995 9760 20059 9764
rect 20075 9820 20139 9824
rect 20075 9764 20079 9820
rect 20079 9764 20135 9820
rect 20135 9764 20139 9820
rect 20075 9760 20139 9764
rect 27609 9820 27673 9824
rect 27609 9764 27613 9820
rect 27613 9764 27669 9820
rect 27669 9764 27673 9820
rect 27609 9760 27673 9764
rect 27689 9820 27753 9824
rect 27689 9764 27693 9820
rect 27693 9764 27749 9820
rect 27749 9764 27753 9820
rect 27689 9760 27753 9764
rect 27769 9820 27833 9824
rect 27769 9764 27773 9820
rect 27773 9764 27829 9820
rect 27829 9764 27833 9820
rect 27769 9760 27833 9764
rect 27849 9820 27913 9824
rect 27849 9764 27853 9820
rect 27853 9764 27909 9820
rect 27909 9764 27913 9820
rect 27849 9760 27913 9764
rect 20484 9556 20548 9620
rect 11836 9420 11900 9484
rect 9628 9284 9692 9348
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 15948 9276 16012 9280
rect 15948 9220 15952 9276
rect 15952 9220 16008 9276
rect 16008 9220 16012 9276
rect 15948 9216 16012 9220
rect 16028 9276 16092 9280
rect 16028 9220 16032 9276
rect 16032 9220 16088 9276
rect 16088 9220 16092 9276
rect 16028 9216 16092 9220
rect 16108 9276 16172 9280
rect 16108 9220 16112 9276
rect 16112 9220 16168 9276
rect 16168 9220 16172 9276
rect 16108 9216 16172 9220
rect 16188 9276 16252 9280
rect 16188 9220 16192 9276
rect 16192 9220 16248 9276
rect 16248 9220 16252 9276
rect 16188 9216 16252 9220
rect 23722 9276 23786 9280
rect 23722 9220 23726 9276
rect 23726 9220 23782 9276
rect 23782 9220 23786 9276
rect 23722 9216 23786 9220
rect 23802 9276 23866 9280
rect 23802 9220 23806 9276
rect 23806 9220 23862 9276
rect 23862 9220 23866 9276
rect 23802 9216 23866 9220
rect 23882 9276 23946 9280
rect 23882 9220 23886 9276
rect 23886 9220 23942 9276
rect 23942 9220 23946 9276
rect 23882 9216 23946 9220
rect 23962 9276 24026 9280
rect 23962 9220 23966 9276
rect 23966 9220 24022 9276
rect 24022 9220 24026 9276
rect 23962 9216 24026 9220
rect 31496 9276 31560 9280
rect 31496 9220 31500 9276
rect 31500 9220 31556 9276
rect 31556 9220 31560 9276
rect 31496 9216 31560 9220
rect 31576 9276 31640 9280
rect 31576 9220 31580 9276
rect 31580 9220 31636 9276
rect 31636 9220 31640 9276
rect 31576 9216 31640 9220
rect 31656 9276 31720 9280
rect 31656 9220 31660 9276
rect 31660 9220 31716 9276
rect 31716 9220 31720 9276
rect 31656 9216 31720 9220
rect 31736 9276 31800 9280
rect 31736 9220 31740 9276
rect 31740 9220 31796 9276
rect 31796 9220 31800 9276
rect 31736 9216 31800 9220
rect 10732 9208 10796 9212
rect 10732 9152 10746 9208
rect 10746 9152 10796 9208
rect 10732 9148 10796 9152
rect 9812 8876 9876 8940
rect 9996 8936 10060 8940
rect 9996 8880 10010 8936
rect 10010 8880 10060 8936
rect 9996 8876 10060 8880
rect 9444 8800 9508 8804
rect 9444 8744 9494 8800
rect 9494 8744 9508 8800
rect 9444 8740 9508 8744
rect 4287 8732 4351 8736
rect 4287 8676 4291 8732
rect 4291 8676 4347 8732
rect 4347 8676 4351 8732
rect 4287 8672 4351 8676
rect 4367 8732 4431 8736
rect 4367 8676 4371 8732
rect 4371 8676 4427 8732
rect 4427 8676 4431 8732
rect 4367 8672 4431 8676
rect 4447 8732 4511 8736
rect 4447 8676 4451 8732
rect 4451 8676 4507 8732
rect 4507 8676 4511 8732
rect 4447 8672 4511 8676
rect 4527 8732 4591 8736
rect 4527 8676 4531 8732
rect 4531 8676 4587 8732
rect 4587 8676 4591 8732
rect 4527 8672 4591 8676
rect 12061 8732 12125 8736
rect 12061 8676 12065 8732
rect 12065 8676 12121 8732
rect 12121 8676 12125 8732
rect 12061 8672 12125 8676
rect 12141 8732 12205 8736
rect 12141 8676 12145 8732
rect 12145 8676 12201 8732
rect 12201 8676 12205 8732
rect 12141 8672 12205 8676
rect 12221 8732 12285 8736
rect 12221 8676 12225 8732
rect 12225 8676 12281 8732
rect 12281 8676 12285 8732
rect 12221 8672 12285 8676
rect 12301 8732 12365 8736
rect 12301 8676 12305 8732
rect 12305 8676 12361 8732
rect 12361 8676 12365 8732
rect 12301 8672 12365 8676
rect 19835 8732 19899 8736
rect 19835 8676 19839 8732
rect 19839 8676 19895 8732
rect 19895 8676 19899 8732
rect 19835 8672 19899 8676
rect 19915 8732 19979 8736
rect 19915 8676 19919 8732
rect 19919 8676 19975 8732
rect 19975 8676 19979 8732
rect 19915 8672 19979 8676
rect 19995 8732 20059 8736
rect 19995 8676 19999 8732
rect 19999 8676 20055 8732
rect 20055 8676 20059 8732
rect 19995 8672 20059 8676
rect 20075 8732 20139 8736
rect 20075 8676 20079 8732
rect 20079 8676 20135 8732
rect 20135 8676 20139 8732
rect 20075 8672 20139 8676
rect 27609 8732 27673 8736
rect 27609 8676 27613 8732
rect 27613 8676 27669 8732
rect 27669 8676 27673 8732
rect 27609 8672 27673 8676
rect 27689 8732 27753 8736
rect 27689 8676 27693 8732
rect 27693 8676 27749 8732
rect 27749 8676 27753 8732
rect 27689 8672 27753 8676
rect 27769 8732 27833 8736
rect 27769 8676 27773 8732
rect 27773 8676 27829 8732
rect 27829 8676 27833 8732
rect 27769 8672 27833 8676
rect 27849 8732 27913 8736
rect 27849 8676 27853 8732
rect 27853 8676 27909 8732
rect 27909 8676 27913 8732
rect 27849 8672 27913 8676
rect 12756 8468 12820 8532
rect 7420 8332 7484 8396
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 10180 8196 10244 8260
rect 12756 8196 12820 8260
rect 9996 8060 10060 8124
rect 15948 8188 16012 8192
rect 15948 8132 15952 8188
rect 15952 8132 16008 8188
rect 16008 8132 16012 8188
rect 15948 8128 16012 8132
rect 16028 8188 16092 8192
rect 16028 8132 16032 8188
rect 16032 8132 16088 8188
rect 16088 8132 16092 8188
rect 16028 8128 16092 8132
rect 16108 8188 16172 8192
rect 16108 8132 16112 8188
rect 16112 8132 16168 8188
rect 16168 8132 16172 8188
rect 16108 8128 16172 8132
rect 16188 8188 16252 8192
rect 16188 8132 16192 8188
rect 16192 8132 16248 8188
rect 16248 8132 16252 8188
rect 16188 8128 16252 8132
rect 23722 8188 23786 8192
rect 23722 8132 23726 8188
rect 23726 8132 23782 8188
rect 23782 8132 23786 8188
rect 23722 8128 23786 8132
rect 23802 8188 23866 8192
rect 23802 8132 23806 8188
rect 23806 8132 23862 8188
rect 23862 8132 23866 8188
rect 23802 8128 23866 8132
rect 23882 8188 23946 8192
rect 23882 8132 23886 8188
rect 23886 8132 23942 8188
rect 23942 8132 23946 8188
rect 23882 8128 23946 8132
rect 23962 8188 24026 8192
rect 23962 8132 23966 8188
rect 23966 8132 24022 8188
rect 24022 8132 24026 8188
rect 23962 8128 24026 8132
rect 31496 8188 31560 8192
rect 31496 8132 31500 8188
rect 31500 8132 31556 8188
rect 31556 8132 31560 8188
rect 31496 8128 31560 8132
rect 31576 8188 31640 8192
rect 31576 8132 31580 8188
rect 31580 8132 31636 8188
rect 31636 8132 31640 8188
rect 31576 8128 31640 8132
rect 31656 8188 31720 8192
rect 31656 8132 31660 8188
rect 31660 8132 31716 8188
rect 31716 8132 31720 8188
rect 31656 8128 31720 8132
rect 31736 8188 31800 8192
rect 31736 8132 31740 8188
rect 31740 8132 31796 8188
rect 31796 8132 31800 8188
rect 31736 8128 31800 8132
rect 6868 7788 6932 7852
rect 7972 7848 8036 7852
rect 7972 7792 8022 7848
rect 8022 7792 8036 7848
rect 7972 7788 8036 7792
rect 8708 7848 8772 7852
rect 8708 7792 8722 7848
rect 8722 7792 8772 7848
rect 8708 7788 8772 7792
rect 5396 7712 5460 7716
rect 5396 7656 5446 7712
rect 5446 7656 5460 7712
rect 5396 7652 5460 7656
rect 10732 7712 10796 7716
rect 10732 7656 10782 7712
rect 10782 7656 10796 7712
rect 4287 7644 4351 7648
rect 4287 7588 4291 7644
rect 4291 7588 4347 7644
rect 4347 7588 4351 7644
rect 4287 7584 4351 7588
rect 4367 7644 4431 7648
rect 4367 7588 4371 7644
rect 4371 7588 4427 7644
rect 4427 7588 4431 7644
rect 4367 7584 4431 7588
rect 4447 7644 4511 7648
rect 4447 7588 4451 7644
rect 4451 7588 4507 7644
rect 4507 7588 4511 7644
rect 4447 7584 4511 7588
rect 4527 7644 4591 7648
rect 4527 7588 4531 7644
rect 4531 7588 4587 7644
rect 4587 7588 4591 7644
rect 4527 7584 4591 7588
rect 6316 7516 6380 7580
rect 10732 7652 10796 7656
rect 11836 7652 11900 7716
rect 12061 7644 12125 7648
rect 12061 7588 12065 7644
rect 12065 7588 12121 7644
rect 12121 7588 12125 7644
rect 12061 7584 12125 7588
rect 12141 7644 12205 7648
rect 12141 7588 12145 7644
rect 12145 7588 12201 7644
rect 12201 7588 12205 7644
rect 12141 7584 12205 7588
rect 12221 7644 12285 7648
rect 12221 7588 12225 7644
rect 12225 7588 12281 7644
rect 12281 7588 12285 7644
rect 12221 7584 12285 7588
rect 12301 7644 12365 7648
rect 12301 7588 12305 7644
rect 12305 7588 12361 7644
rect 12361 7588 12365 7644
rect 12301 7584 12365 7588
rect 19835 7644 19899 7648
rect 19835 7588 19839 7644
rect 19839 7588 19895 7644
rect 19895 7588 19899 7644
rect 19835 7584 19899 7588
rect 19915 7644 19979 7648
rect 19915 7588 19919 7644
rect 19919 7588 19975 7644
rect 19975 7588 19979 7644
rect 19915 7584 19979 7588
rect 19995 7644 20059 7648
rect 19995 7588 19999 7644
rect 19999 7588 20055 7644
rect 20055 7588 20059 7644
rect 19995 7584 20059 7588
rect 20075 7644 20139 7648
rect 20075 7588 20079 7644
rect 20079 7588 20135 7644
rect 20135 7588 20139 7644
rect 20075 7584 20139 7588
rect 27609 7644 27673 7648
rect 27609 7588 27613 7644
rect 27613 7588 27669 7644
rect 27669 7588 27673 7644
rect 27609 7584 27673 7588
rect 27689 7644 27753 7648
rect 27689 7588 27693 7644
rect 27693 7588 27749 7644
rect 27749 7588 27753 7644
rect 27689 7584 27753 7588
rect 27769 7644 27833 7648
rect 27769 7588 27773 7644
rect 27773 7588 27829 7644
rect 27829 7588 27833 7644
rect 27769 7584 27833 7588
rect 27849 7644 27913 7648
rect 27849 7588 27853 7644
rect 27853 7588 27909 7644
rect 27909 7588 27913 7644
rect 27849 7584 27913 7588
rect 10548 7516 10612 7580
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 15948 7100 16012 7104
rect 15948 7044 15952 7100
rect 15952 7044 16008 7100
rect 16008 7044 16012 7100
rect 15948 7040 16012 7044
rect 16028 7100 16092 7104
rect 16028 7044 16032 7100
rect 16032 7044 16088 7100
rect 16088 7044 16092 7100
rect 16028 7040 16092 7044
rect 16108 7100 16172 7104
rect 16108 7044 16112 7100
rect 16112 7044 16168 7100
rect 16168 7044 16172 7100
rect 16108 7040 16172 7044
rect 16188 7100 16252 7104
rect 16188 7044 16192 7100
rect 16192 7044 16248 7100
rect 16248 7044 16252 7100
rect 16188 7040 16252 7044
rect 23722 7100 23786 7104
rect 23722 7044 23726 7100
rect 23726 7044 23782 7100
rect 23782 7044 23786 7100
rect 23722 7040 23786 7044
rect 23802 7100 23866 7104
rect 23802 7044 23806 7100
rect 23806 7044 23862 7100
rect 23862 7044 23866 7100
rect 23802 7040 23866 7044
rect 23882 7100 23946 7104
rect 23882 7044 23886 7100
rect 23886 7044 23942 7100
rect 23942 7044 23946 7100
rect 23882 7040 23946 7044
rect 23962 7100 24026 7104
rect 23962 7044 23966 7100
rect 23966 7044 24022 7100
rect 24022 7044 24026 7100
rect 23962 7040 24026 7044
rect 31496 7100 31560 7104
rect 31496 7044 31500 7100
rect 31500 7044 31556 7100
rect 31556 7044 31560 7100
rect 31496 7040 31560 7044
rect 31576 7100 31640 7104
rect 31576 7044 31580 7100
rect 31580 7044 31636 7100
rect 31636 7044 31640 7100
rect 31576 7040 31640 7044
rect 31656 7100 31720 7104
rect 31656 7044 31660 7100
rect 31660 7044 31716 7100
rect 31716 7044 31720 7100
rect 31656 7040 31720 7044
rect 31736 7100 31800 7104
rect 31736 7044 31740 7100
rect 31740 7044 31796 7100
rect 31796 7044 31800 7100
rect 31736 7040 31800 7044
rect 9444 6972 9508 7036
rect 10916 6972 10980 7036
rect 8708 6700 8772 6764
rect 6316 6564 6380 6628
rect 4287 6556 4351 6560
rect 4287 6500 4291 6556
rect 4291 6500 4347 6556
rect 4347 6500 4351 6556
rect 4287 6496 4351 6500
rect 4367 6556 4431 6560
rect 4367 6500 4371 6556
rect 4371 6500 4427 6556
rect 4427 6500 4431 6556
rect 4367 6496 4431 6500
rect 4447 6556 4511 6560
rect 4447 6500 4451 6556
rect 4451 6500 4507 6556
rect 4507 6500 4511 6556
rect 4447 6496 4511 6500
rect 4527 6556 4591 6560
rect 4527 6500 4531 6556
rect 4531 6500 4587 6556
rect 4587 6500 4591 6556
rect 4527 6496 4591 6500
rect 12061 6556 12125 6560
rect 12061 6500 12065 6556
rect 12065 6500 12121 6556
rect 12121 6500 12125 6556
rect 12061 6496 12125 6500
rect 12141 6556 12205 6560
rect 12141 6500 12145 6556
rect 12145 6500 12201 6556
rect 12201 6500 12205 6556
rect 12141 6496 12205 6500
rect 12221 6556 12285 6560
rect 12221 6500 12225 6556
rect 12225 6500 12281 6556
rect 12281 6500 12285 6556
rect 12221 6496 12285 6500
rect 12301 6556 12365 6560
rect 12301 6500 12305 6556
rect 12305 6500 12361 6556
rect 12361 6500 12365 6556
rect 12301 6496 12365 6500
rect 19835 6556 19899 6560
rect 19835 6500 19839 6556
rect 19839 6500 19895 6556
rect 19895 6500 19899 6556
rect 19835 6496 19899 6500
rect 19915 6556 19979 6560
rect 19915 6500 19919 6556
rect 19919 6500 19975 6556
rect 19975 6500 19979 6556
rect 19915 6496 19979 6500
rect 19995 6556 20059 6560
rect 19995 6500 19999 6556
rect 19999 6500 20055 6556
rect 20055 6500 20059 6556
rect 19995 6496 20059 6500
rect 20075 6556 20139 6560
rect 20075 6500 20079 6556
rect 20079 6500 20135 6556
rect 20135 6500 20139 6556
rect 20075 6496 20139 6500
rect 27609 6556 27673 6560
rect 27609 6500 27613 6556
rect 27613 6500 27669 6556
rect 27669 6500 27673 6556
rect 27609 6496 27673 6500
rect 27689 6556 27753 6560
rect 27689 6500 27693 6556
rect 27693 6500 27749 6556
rect 27749 6500 27753 6556
rect 27689 6496 27753 6500
rect 27769 6556 27833 6560
rect 27769 6500 27773 6556
rect 27773 6500 27829 6556
rect 27829 6500 27833 6556
rect 27769 6496 27833 6500
rect 27849 6556 27913 6560
rect 27849 6500 27853 6556
rect 27853 6500 27909 6556
rect 27909 6500 27913 6556
rect 27849 6496 27913 6500
rect 7420 6020 7484 6084
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 7052 5884 7116 5948
rect 9812 6080 9876 6084
rect 9812 6024 9826 6080
rect 9826 6024 9876 6080
rect 9812 6020 9876 6024
rect 15948 6012 16012 6016
rect 15948 5956 15952 6012
rect 15952 5956 16008 6012
rect 16008 5956 16012 6012
rect 15948 5952 16012 5956
rect 16028 6012 16092 6016
rect 16028 5956 16032 6012
rect 16032 5956 16088 6012
rect 16088 5956 16092 6012
rect 16028 5952 16092 5956
rect 16108 6012 16172 6016
rect 16108 5956 16112 6012
rect 16112 5956 16168 6012
rect 16168 5956 16172 6012
rect 16108 5952 16172 5956
rect 16188 6012 16252 6016
rect 16188 5956 16192 6012
rect 16192 5956 16248 6012
rect 16248 5956 16252 6012
rect 16188 5952 16252 5956
rect 23722 6012 23786 6016
rect 23722 5956 23726 6012
rect 23726 5956 23782 6012
rect 23782 5956 23786 6012
rect 23722 5952 23786 5956
rect 23802 6012 23866 6016
rect 23802 5956 23806 6012
rect 23806 5956 23862 6012
rect 23862 5956 23866 6012
rect 23802 5952 23866 5956
rect 23882 6012 23946 6016
rect 23882 5956 23886 6012
rect 23886 5956 23942 6012
rect 23942 5956 23946 6012
rect 23882 5952 23946 5956
rect 23962 6012 24026 6016
rect 23962 5956 23966 6012
rect 23966 5956 24022 6012
rect 24022 5956 24026 6012
rect 23962 5952 24026 5956
rect 31496 6012 31560 6016
rect 31496 5956 31500 6012
rect 31500 5956 31556 6012
rect 31556 5956 31560 6012
rect 31496 5952 31560 5956
rect 31576 6012 31640 6016
rect 31576 5956 31580 6012
rect 31580 5956 31636 6012
rect 31636 5956 31640 6012
rect 31576 5952 31640 5956
rect 31656 6012 31720 6016
rect 31656 5956 31660 6012
rect 31660 5956 31716 6012
rect 31716 5956 31720 6012
rect 31656 5952 31720 5956
rect 31736 6012 31800 6016
rect 31736 5956 31740 6012
rect 31740 5956 31796 6012
rect 31796 5956 31800 6012
rect 31736 5952 31800 5956
rect 6868 5612 6932 5676
rect 4287 5468 4351 5472
rect 4287 5412 4291 5468
rect 4291 5412 4347 5468
rect 4347 5412 4351 5468
rect 4287 5408 4351 5412
rect 4367 5468 4431 5472
rect 4367 5412 4371 5468
rect 4371 5412 4427 5468
rect 4427 5412 4431 5468
rect 4367 5408 4431 5412
rect 4447 5468 4511 5472
rect 4447 5412 4451 5468
rect 4451 5412 4507 5468
rect 4507 5412 4511 5468
rect 4447 5408 4511 5412
rect 4527 5468 4591 5472
rect 4527 5412 4531 5468
rect 4531 5412 4587 5468
rect 4587 5412 4591 5468
rect 4527 5408 4591 5412
rect 12061 5468 12125 5472
rect 12061 5412 12065 5468
rect 12065 5412 12121 5468
rect 12121 5412 12125 5468
rect 12061 5408 12125 5412
rect 12141 5468 12205 5472
rect 12141 5412 12145 5468
rect 12145 5412 12201 5468
rect 12201 5412 12205 5468
rect 12141 5408 12205 5412
rect 12221 5468 12285 5472
rect 12221 5412 12225 5468
rect 12225 5412 12281 5468
rect 12281 5412 12285 5468
rect 12221 5408 12285 5412
rect 12301 5468 12365 5472
rect 12301 5412 12305 5468
rect 12305 5412 12361 5468
rect 12361 5412 12365 5468
rect 12301 5408 12365 5412
rect 10548 5128 10612 5132
rect 19835 5468 19899 5472
rect 19835 5412 19839 5468
rect 19839 5412 19895 5468
rect 19895 5412 19899 5468
rect 19835 5408 19899 5412
rect 19915 5468 19979 5472
rect 19915 5412 19919 5468
rect 19919 5412 19975 5468
rect 19975 5412 19979 5468
rect 19915 5408 19979 5412
rect 19995 5468 20059 5472
rect 19995 5412 19999 5468
rect 19999 5412 20055 5468
rect 20055 5412 20059 5468
rect 19995 5408 20059 5412
rect 20075 5468 20139 5472
rect 20075 5412 20079 5468
rect 20079 5412 20135 5468
rect 20135 5412 20139 5468
rect 20075 5408 20139 5412
rect 27609 5468 27673 5472
rect 27609 5412 27613 5468
rect 27613 5412 27669 5468
rect 27669 5412 27673 5468
rect 27609 5408 27673 5412
rect 27689 5468 27753 5472
rect 27689 5412 27693 5468
rect 27693 5412 27749 5468
rect 27749 5412 27753 5468
rect 27689 5408 27753 5412
rect 27769 5468 27833 5472
rect 27769 5412 27773 5468
rect 27773 5412 27829 5468
rect 27829 5412 27833 5468
rect 27769 5408 27833 5412
rect 27849 5468 27913 5472
rect 27849 5412 27853 5468
rect 27853 5412 27909 5468
rect 27909 5412 27913 5468
rect 27849 5408 27913 5412
rect 10548 5072 10598 5128
rect 10598 5072 10612 5128
rect 10548 5068 10612 5072
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 15948 4924 16012 4928
rect 15948 4868 15952 4924
rect 15952 4868 16008 4924
rect 16008 4868 16012 4924
rect 15948 4864 16012 4868
rect 16028 4924 16092 4928
rect 16028 4868 16032 4924
rect 16032 4868 16088 4924
rect 16088 4868 16092 4924
rect 16028 4864 16092 4868
rect 16108 4924 16172 4928
rect 16108 4868 16112 4924
rect 16112 4868 16168 4924
rect 16168 4868 16172 4924
rect 16108 4864 16172 4868
rect 16188 4924 16252 4928
rect 16188 4868 16192 4924
rect 16192 4868 16248 4924
rect 16248 4868 16252 4924
rect 16188 4864 16252 4868
rect 23722 4924 23786 4928
rect 23722 4868 23726 4924
rect 23726 4868 23782 4924
rect 23782 4868 23786 4924
rect 23722 4864 23786 4868
rect 23802 4924 23866 4928
rect 23802 4868 23806 4924
rect 23806 4868 23862 4924
rect 23862 4868 23866 4924
rect 23802 4864 23866 4868
rect 23882 4924 23946 4928
rect 23882 4868 23886 4924
rect 23886 4868 23942 4924
rect 23942 4868 23946 4924
rect 23882 4864 23946 4868
rect 23962 4924 24026 4928
rect 23962 4868 23966 4924
rect 23966 4868 24022 4924
rect 24022 4868 24026 4924
rect 23962 4864 24026 4868
rect 31496 4924 31560 4928
rect 31496 4868 31500 4924
rect 31500 4868 31556 4924
rect 31556 4868 31560 4924
rect 31496 4864 31560 4868
rect 31576 4924 31640 4928
rect 31576 4868 31580 4924
rect 31580 4868 31636 4924
rect 31636 4868 31640 4924
rect 31576 4864 31640 4868
rect 31656 4924 31720 4928
rect 31656 4868 31660 4924
rect 31660 4868 31716 4924
rect 31716 4868 31720 4924
rect 31656 4864 31720 4868
rect 31736 4924 31800 4928
rect 31736 4868 31740 4924
rect 31740 4868 31796 4924
rect 31796 4868 31800 4924
rect 31736 4864 31800 4868
rect 4287 4380 4351 4384
rect 4287 4324 4291 4380
rect 4291 4324 4347 4380
rect 4347 4324 4351 4380
rect 4287 4320 4351 4324
rect 4367 4380 4431 4384
rect 4367 4324 4371 4380
rect 4371 4324 4427 4380
rect 4427 4324 4431 4380
rect 4367 4320 4431 4324
rect 4447 4380 4511 4384
rect 4447 4324 4451 4380
rect 4451 4324 4507 4380
rect 4507 4324 4511 4380
rect 4447 4320 4511 4324
rect 4527 4380 4591 4384
rect 4527 4324 4531 4380
rect 4531 4324 4587 4380
rect 4587 4324 4591 4380
rect 4527 4320 4591 4324
rect 12061 4380 12125 4384
rect 12061 4324 12065 4380
rect 12065 4324 12121 4380
rect 12121 4324 12125 4380
rect 12061 4320 12125 4324
rect 12141 4380 12205 4384
rect 12141 4324 12145 4380
rect 12145 4324 12201 4380
rect 12201 4324 12205 4380
rect 12141 4320 12205 4324
rect 12221 4380 12285 4384
rect 12221 4324 12225 4380
rect 12225 4324 12281 4380
rect 12281 4324 12285 4380
rect 12221 4320 12285 4324
rect 12301 4380 12365 4384
rect 12301 4324 12305 4380
rect 12305 4324 12361 4380
rect 12361 4324 12365 4380
rect 12301 4320 12365 4324
rect 19835 4380 19899 4384
rect 19835 4324 19839 4380
rect 19839 4324 19895 4380
rect 19895 4324 19899 4380
rect 19835 4320 19899 4324
rect 19915 4380 19979 4384
rect 19915 4324 19919 4380
rect 19919 4324 19975 4380
rect 19975 4324 19979 4380
rect 19915 4320 19979 4324
rect 19995 4380 20059 4384
rect 19995 4324 19999 4380
rect 19999 4324 20055 4380
rect 20055 4324 20059 4380
rect 19995 4320 20059 4324
rect 20075 4380 20139 4384
rect 20075 4324 20079 4380
rect 20079 4324 20135 4380
rect 20135 4324 20139 4380
rect 20075 4320 20139 4324
rect 27609 4380 27673 4384
rect 27609 4324 27613 4380
rect 27613 4324 27669 4380
rect 27669 4324 27673 4380
rect 27609 4320 27673 4324
rect 27689 4380 27753 4384
rect 27689 4324 27693 4380
rect 27693 4324 27749 4380
rect 27749 4324 27753 4380
rect 27689 4320 27753 4324
rect 27769 4380 27833 4384
rect 27769 4324 27773 4380
rect 27773 4324 27829 4380
rect 27829 4324 27833 4380
rect 27769 4320 27833 4324
rect 27849 4380 27913 4384
rect 27849 4324 27853 4380
rect 27853 4324 27909 4380
rect 27909 4324 27913 4380
rect 27849 4320 27913 4324
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 15948 3836 16012 3840
rect 15948 3780 15952 3836
rect 15952 3780 16008 3836
rect 16008 3780 16012 3836
rect 15948 3776 16012 3780
rect 16028 3836 16092 3840
rect 16028 3780 16032 3836
rect 16032 3780 16088 3836
rect 16088 3780 16092 3836
rect 16028 3776 16092 3780
rect 16108 3836 16172 3840
rect 16108 3780 16112 3836
rect 16112 3780 16168 3836
rect 16168 3780 16172 3836
rect 16108 3776 16172 3780
rect 16188 3836 16252 3840
rect 16188 3780 16192 3836
rect 16192 3780 16248 3836
rect 16248 3780 16252 3836
rect 16188 3776 16252 3780
rect 23722 3836 23786 3840
rect 23722 3780 23726 3836
rect 23726 3780 23782 3836
rect 23782 3780 23786 3836
rect 23722 3776 23786 3780
rect 23802 3836 23866 3840
rect 23802 3780 23806 3836
rect 23806 3780 23862 3836
rect 23862 3780 23866 3836
rect 23802 3776 23866 3780
rect 23882 3836 23946 3840
rect 23882 3780 23886 3836
rect 23886 3780 23942 3836
rect 23942 3780 23946 3836
rect 23882 3776 23946 3780
rect 23962 3836 24026 3840
rect 23962 3780 23966 3836
rect 23966 3780 24022 3836
rect 24022 3780 24026 3836
rect 23962 3776 24026 3780
rect 31496 3836 31560 3840
rect 31496 3780 31500 3836
rect 31500 3780 31556 3836
rect 31556 3780 31560 3836
rect 31496 3776 31560 3780
rect 31576 3836 31640 3840
rect 31576 3780 31580 3836
rect 31580 3780 31636 3836
rect 31636 3780 31640 3836
rect 31576 3776 31640 3780
rect 31656 3836 31720 3840
rect 31656 3780 31660 3836
rect 31660 3780 31716 3836
rect 31716 3780 31720 3836
rect 31656 3776 31720 3780
rect 31736 3836 31800 3840
rect 31736 3780 31740 3836
rect 31740 3780 31796 3836
rect 31796 3780 31800 3836
rect 31736 3776 31800 3780
rect 4287 3292 4351 3296
rect 4287 3236 4291 3292
rect 4291 3236 4347 3292
rect 4347 3236 4351 3292
rect 4287 3232 4351 3236
rect 4367 3292 4431 3296
rect 4367 3236 4371 3292
rect 4371 3236 4427 3292
rect 4427 3236 4431 3292
rect 4367 3232 4431 3236
rect 4447 3292 4511 3296
rect 4447 3236 4451 3292
rect 4451 3236 4507 3292
rect 4507 3236 4511 3292
rect 4447 3232 4511 3236
rect 4527 3292 4591 3296
rect 4527 3236 4531 3292
rect 4531 3236 4587 3292
rect 4587 3236 4591 3292
rect 4527 3232 4591 3236
rect 12061 3292 12125 3296
rect 12061 3236 12065 3292
rect 12065 3236 12121 3292
rect 12121 3236 12125 3292
rect 12061 3232 12125 3236
rect 12141 3292 12205 3296
rect 12141 3236 12145 3292
rect 12145 3236 12201 3292
rect 12201 3236 12205 3292
rect 12141 3232 12205 3236
rect 12221 3292 12285 3296
rect 12221 3236 12225 3292
rect 12225 3236 12281 3292
rect 12281 3236 12285 3292
rect 12221 3232 12285 3236
rect 12301 3292 12365 3296
rect 12301 3236 12305 3292
rect 12305 3236 12361 3292
rect 12361 3236 12365 3292
rect 12301 3232 12365 3236
rect 19835 3292 19899 3296
rect 19835 3236 19839 3292
rect 19839 3236 19895 3292
rect 19895 3236 19899 3292
rect 19835 3232 19899 3236
rect 19915 3292 19979 3296
rect 19915 3236 19919 3292
rect 19919 3236 19975 3292
rect 19975 3236 19979 3292
rect 19915 3232 19979 3236
rect 19995 3292 20059 3296
rect 19995 3236 19999 3292
rect 19999 3236 20055 3292
rect 20055 3236 20059 3292
rect 19995 3232 20059 3236
rect 20075 3292 20139 3296
rect 20075 3236 20079 3292
rect 20079 3236 20135 3292
rect 20135 3236 20139 3292
rect 20075 3232 20139 3236
rect 27609 3292 27673 3296
rect 27609 3236 27613 3292
rect 27613 3236 27669 3292
rect 27669 3236 27673 3292
rect 27609 3232 27673 3236
rect 27689 3292 27753 3296
rect 27689 3236 27693 3292
rect 27693 3236 27749 3292
rect 27749 3236 27753 3292
rect 27689 3232 27753 3236
rect 27769 3292 27833 3296
rect 27769 3236 27773 3292
rect 27773 3236 27829 3292
rect 27829 3236 27833 3292
rect 27769 3232 27833 3236
rect 27849 3292 27913 3296
rect 27849 3236 27853 3292
rect 27853 3236 27909 3292
rect 27909 3236 27913 3292
rect 27849 3232 27913 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 15948 2748 16012 2752
rect 15948 2692 15952 2748
rect 15952 2692 16008 2748
rect 16008 2692 16012 2748
rect 15948 2688 16012 2692
rect 16028 2748 16092 2752
rect 16028 2692 16032 2748
rect 16032 2692 16088 2748
rect 16088 2692 16092 2748
rect 16028 2688 16092 2692
rect 16108 2748 16172 2752
rect 16108 2692 16112 2748
rect 16112 2692 16168 2748
rect 16168 2692 16172 2748
rect 16108 2688 16172 2692
rect 16188 2748 16252 2752
rect 16188 2692 16192 2748
rect 16192 2692 16248 2748
rect 16248 2692 16252 2748
rect 16188 2688 16252 2692
rect 23722 2748 23786 2752
rect 23722 2692 23726 2748
rect 23726 2692 23782 2748
rect 23782 2692 23786 2748
rect 23722 2688 23786 2692
rect 23802 2748 23866 2752
rect 23802 2692 23806 2748
rect 23806 2692 23862 2748
rect 23862 2692 23866 2748
rect 23802 2688 23866 2692
rect 23882 2748 23946 2752
rect 23882 2692 23886 2748
rect 23886 2692 23942 2748
rect 23942 2692 23946 2748
rect 23882 2688 23946 2692
rect 23962 2748 24026 2752
rect 23962 2692 23966 2748
rect 23966 2692 24022 2748
rect 24022 2692 24026 2748
rect 23962 2688 24026 2692
rect 31496 2748 31560 2752
rect 31496 2692 31500 2748
rect 31500 2692 31556 2748
rect 31556 2692 31560 2748
rect 31496 2688 31560 2692
rect 31576 2748 31640 2752
rect 31576 2692 31580 2748
rect 31580 2692 31636 2748
rect 31636 2692 31640 2748
rect 31576 2688 31640 2692
rect 31656 2748 31720 2752
rect 31656 2692 31660 2748
rect 31660 2692 31716 2748
rect 31716 2692 31720 2748
rect 31656 2688 31720 2692
rect 31736 2748 31800 2752
rect 31736 2692 31740 2748
rect 31740 2692 31796 2748
rect 31796 2692 31800 2748
rect 31736 2688 31800 2692
rect 4287 2204 4351 2208
rect 4287 2148 4291 2204
rect 4291 2148 4347 2204
rect 4347 2148 4351 2204
rect 4287 2144 4351 2148
rect 4367 2204 4431 2208
rect 4367 2148 4371 2204
rect 4371 2148 4427 2204
rect 4427 2148 4431 2204
rect 4367 2144 4431 2148
rect 4447 2204 4511 2208
rect 4447 2148 4451 2204
rect 4451 2148 4507 2204
rect 4507 2148 4511 2204
rect 4447 2144 4511 2148
rect 4527 2204 4591 2208
rect 4527 2148 4531 2204
rect 4531 2148 4587 2204
rect 4587 2148 4591 2204
rect 4527 2144 4591 2148
rect 12061 2204 12125 2208
rect 12061 2148 12065 2204
rect 12065 2148 12121 2204
rect 12121 2148 12125 2204
rect 12061 2144 12125 2148
rect 12141 2204 12205 2208
rect 12141 2148 12145 2204
rect 12145 2148 12201 2204
rect 12201 2148 12205 2204
rect 12141 2144 12205 2148
rect 12221 2204 12285 2208
rect 12221 2148 12225 2204
rect 12225 2148 12281 2204
rect 12281 2148 12285 2204
rect 12221 2144 12285 2148
rect 12301 2204 12365 2208
rect 12301 2148 12305 2204
rect 12305 2148 12361 2204
rect 12361 2148 12365 2204
rect 12301 2144 12365 2148
rect 19835 2204 19899 2208
rect 19835 2148 19839 2204
rect 19839 2148 19895 2204
rect 19895 2148 19899 2204
rect 19835 2144 19899 2148
rect 19915 2204 19979 2208
rect 19915 2148 19919 2204
rect 19919 2148 19975 2204
rect 19975 2148 19979 2204
rect 19915 2144 19979 2148
rect 19995 2204 20059 2208
rect 19995 2148 19999 2204
rect 19999 2148 20055 2204
rect 20055 2148 20059 2204
rect 19995 2144 20059 2148
rect 20075 2204 20139 2208
rect 20075 2148 20079 2204
rect 20079 2148 20135 2204
rect 20135 2148 20139 2204
rect 20075 2144 20139 2148
rect 27609 2204 27673 2208
rect 27609 2148 27613 2204
rect 27613 2148 27669 2204
rect 27669 2148 27673 2204
rect 27609 2144 27673 2148
rect 27689 2204 27753 2208
rect 27689 2148 27693 2204
rect 27693 2148 27749 2204
rect 27749 2148 27753 2204
rect 27689 2144 27753 2148
rect 27769 2204 27833 2208
rect 27769 2148 27773 2204
rect 27773 2148 27829 2204
rect 27829 2148 27833 2204
rect 27769 2144 27833 2148
rect 27849 2204 27913 2208
rect 27849 2148 27853 2204
rect 27853 2148 27909 2204
rect 27909 2148 27913 2204
rect 27849 2144 27913 2148
rect 8174 1660 8238 1664
rect 8174 1604 8178 1660
rect 8178 1604 8234 1660
rect 8234 1604 8238 1660
rect 8174 1600 8238 1604
rect 8254 1660 8318 1664
rect 8254 1604 8258 1660
rect 8258 1604 8314 1660
rect 8314 1604 8318 1660
rect 8254 1600 8318 1604
rect 8334 1660 8398 1664
rect 8334 1604 8338 1660
rect 8338 1604 8394 1660
rect 8394 1604 8398 1660
rect 8334 1600 8398 1604
rect 8414 1660 8478 1664
rect 8414 1604 8418 1660
rect 8418 1604 8474 1660
rect 8474 1604 8478 1660
rect 8414 1600 8478 1604
rect 15948 1660 16012 1664
rect 15948 1604 15952 1660
rect 15952 1604 16008 1660
rect 16008 1604 16012 1660
rect 15948 1600 16012 1604
rect 16028 1660 16092 1664
rect 16028 1604 16032 1660
rect 16032 1604 16088 1660
rect 16088 1604 16092 1660
rect 16028 1600 16092 1604
rect 16108 1660 16172 1664
rect 16108 1604 16112 1660
rect 16112 1604 16168 1660
rect 16168 1604 16172 1660
rect 16108 1600 16172 1604
rect 16188 1660 16252 1664
rect 16188 1604 16192 1660
rect 16192 1604 16248 1660
rect 16248 1604 16252 1660
rect 16188 1600 16252 1604
rect 23722 1660 23786 1664
rect 23722 1604 23726 1660
rect 23726 1604 23782 1660
rect 23782 1604 23786 1660
rect 23722 1600 23786 1604
rect 23802 1660 23866 1664
rect 23802 1604 23806 1660
rect 23806 1604 23862 1660
rect 23862 1604 23866 1660
rect 23802 1600 23866 1604
rect 23882 1660 23946 1664
rect 23882 1604 23886 1660
rect 23886 1604 23942 1660
rect 23942 1604 23946 1660
rect 23882 1600 23946 1604
rect 23962 1660 24026 1664
rect 23962 1604 23966 1660
rect 23966 1604 24022 1660
rect 24022 1604 24026 1660
rect 23962 1600 24026 1604
rect 31496 1660 31560 1664
rect 31496 1604 31500 1660
rect 31500 1604 31556 1660
rect 31556 1604 31560 1660
rect 31496 1600 31560 1604
rect 31576 1660 31640 1664
rect 31576 1604 31580 1660
rect 31580 1604 31636 1660
rect 31636 1604 31640 1660
rect 31576 1600 31640 1604
rect 31656 1660 31720 1664
rect 31656 1604 31660 1660
rect 31660 1604 31716 1660
rect 31716 1604 31720 1660
rect 31656 1600 31720 1604
rect 31736 1660 31800 1664
rect 31736 1604 31740 1660
rect 31740 1604 31796 1660
rect 31796 1604 31800 1660
rect 31736 1600 31800 1604
rect 4287 1116 4351 1120
rect 4287 1060 4291 1116
rect 4291 1060 4347 1116
rect 4347 1060 4351 1116
rect 4287 1056 4351 1060
rect 4367 1116 4431 1120
rect 4367 1060 4371 1116
rect 4371 1060 4427 1116
rect 4427 1060 4431 1116
rect 4367 1056 4431 1060
rect 4447 1116 4511 1120
rect 4447 1060 4451 1116
rect 4451 1060 4507 1116
rect 4507 1060 4511 1116
rect 4447 1056 4511 1060
rect 4527 1116 4591 1120
rect 4527 1060 4531 1116
rect 4531 1060 4587 1116
rect 4587 1060 4591 1116
rect 4527 1056 4591 1060
rect 12061 1116 12125 1120
rect 12061 1060 12065 1116
rect 12065 1060 12121 1116
rect 12121 1060 12125 1116
rect 12061 1056 12125 1060
rect 12141 1116 12205 1120
rect 12141 1060 12145 1116
rect 12145 1060 12201 1116
rect 12201 1060 12205 1116
rect 12141 1056 12205 1060
rect 12221 1116 12285 1120
rect 12221 1060 12225 1116
rect 12225 1060 12281 1116
rect 12281 1060 12285 1116
rect 12221 1056 12285 1060
rect 12301 1116 12365 1120
rect 12301 1060 12305 1116
rect 12305 1060 12361 1116
rect 12361 1060 12365 1116
rect 12301 1056 12365 1060
rect 19835 1116 19899 1120
rect 19835 1060 19839 1116
rect 19839 1060 19895 1116
rect 19895 1060 19899 1116
rect 19835 1056 19899 1060
rect 19915 1116 19979 1120
rect 19915 1060 19919 1116
rect 19919 1060 19975 1116
rect 19975 1060 19979 1116
rect 19915 1056 19979 1060
rect 19995 1116 20059 1120
rect 19995 1060 19999 1116
rect 19999 1060 20055 1116
rect 20055 1060 20059 1116
rect 19995 1056 20059 1060
rect 20075 1116 20139 1120
rect 20075 1060 20079 1116
rect 20079 1060 20135 1116
rect 20135 1060 20139 1116
rect 20075 1056 20139 1060
rect 27609 1116 27673 1120
rect 27609 1060 27613 1116
rect 27613 1060 27669 1116
rect 27669 1060 27673 1116
rect 27609 1056 27673 1060
rect 27689 1116 27753 1120
rect 27689 1060 27693 1116
rect 27693 1060 27749 1116
rect 27749 1060 27753 1116
rect 27689 1056 27753 1060
rect 27769 1116 27833 1120
rect 27769 1060 27773 1116
rect 27773 1060 27829 1116
rect 27829 1060 27833 1116
rect 27769 1056 27833 1060
rect 27849 1116 27913 1120
rect 27849 1060 27853 1116
rect 27853 1060 27909 1116
rect 27909 1060 27913 1116
rect 27849 1056 27913 1060
rect 8174 572 8238 576
rect 8174 516 8178 572
rect 8178 516 8234 572
rect 8234 516 8238 572
rect 8174 512 8238 516
rect 8254 572 8318 576
rect 8254 516 8258 572
rect 8258 516 8314 572
rect 8314 516 8318 572
rect 8254 512 8318 516
rect 8334 572 8398 576
rect 8334 516 8338 572
rect 8338 516 8394 572
rect 8394 516 8398 572
rect 8334 512 8398 516
rect 8414 572 8478 576
rect 8414 516 8418 572
rect 8418 516 8474 572
rect 8474 516 8478 572
rect 8414 512 8478 516
rect 15948 572 16012 576
rect 15948 516 15952 572
rect 15952 516 16008 572
rect 16008 516 16012 572
rect 15948 512 16012 516
rect 16028 572 16092 576
rect 16028 516 16032 572
rect 16032 516 16088 572
rect 16088 516 16092 572
rect 16028 512 16092 516
rect 16108 572 16172 576
rect 16108 516 16112 572
rect 16112 516 16168 572
rect 16168 516 16172 572
rect 16108 512 16172 516
rect 16188 572 16252 576
rect 16188 516 16192 572
rect 16192 516 16248 572
rect 16248 516 16252 572
rect 16188 512 16252 516
rect 23722 572 23786 576
rect 23722 516 23726 572
rect 23726 516 23782 572
rect 23782 516 23786 572
rect 23722 512 23786 516
rect 23802 572 23866 576
rect 23802 516 23806 572
rect 23806 516 23862 572
rect 23862 516 23866 572
rect 23802 512 23866 516
rect 23882 572 23946 576
rect 23882 516 23886 572
rect 23886 516 23942 572
rect 23942 516 23946 572
rect 23882 512 23946 516
rect 23962 572 24026 576
rect 23962 516 23966 572
rect 23966 516 24022 572
rect 24022 516 24026 572
rect 23962 512 24026 516
rect 31496 572 31560 576
rect 31496 516 31500 572
rect 31500 516 31556 572
rect 31556 516 31560 572
rect 31496 512 31560 516
rect 31576 572 31640 576
rect 31576 516 31580 572
rect 31580 516 31636 572
rect 31636 516 31640 572
rect 31576 512 31640 516
rect 31656 572 31720 576
rect 31656 516 31660 572
rect 31660 516 31716 572
rect 31716 516 31720 572
rect 31656 512 31720 516
rect 31736 572 31800 576
rect 31736 516 31740 572
rect 31740 516 31796 572
rect 31796 516 31800 572
rect 31736 512 31800 516
<< metal4 >>
rect 798 21317 858 22304
rect 795 21316 861 21317
rect 795 21252 796 21316
rect 860 21252 861 21316
rect 795 21251 861 21252
rect 1534 21181 1594 22304
rect 1531 21180 1597 21181
rect 1531 21116 1532 21180
rect 1596 21116 1597 21180
rect 1531 21115 1597 21116
rect 2270 20773 2330 22304
rect 3006 21181 3066 22304
rect 3742 21589 3802 22304
rect 4478 21997 4538 22304
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 4279 21792 4599 21808
rect 4279 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4599 21792
rect 3739 21588 3805 21589
rect 3739 21524 3740 21588
rect 3804 21524 3805 21588
rect 3739 21523 3805 21524
rect 3003 21180 3069 21181
rect 3003 21116 3004 21180
rect 3068 21116 3069 21180
rect 3003 21115 3069 21116
rect 2267 20772 2333 20773
rect 2267 20708 2268 20772
rect 2332 20708 2333 20772
rect 2267 20707 2333 20708
rect 4279 20704 4599 21728
rect 4279 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4599 20704
rect 4279 19616 4599 20640
rect 4279 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4599 19616
rect 4279 18528 4599 19552
rect 5214 19277 5274 22304
rect 5950 21181 6010 22304
rect 6686 21861 6746 22304
rect 7422 21861 7482 22304
rect 8158 22130 8218 22304
rect 7974 22070 8218 22130
rect 8894 22130 8954 22304
rect 9078 22174 9506 22234
rect 9078 22130 9138 22174
rect 8894 22070 9138 22130
rect 6683 21860 6749 21861
rect 6683 21796 6684 21860
rect 6748 21796 6749 21860
rect 6683 21795 6749 21796
rect 7419 21860 7485 21861
rect 7419 21796 7420 21860
rect 7484 21796 7485 21860
rect 7419 21795 7485 21796
rect 5947 21180 6013 21181
rect 5947 21116 5948 21180
rect 6012 21116 6013 21180
rect 5947 21115 6013 21116
rect 6315 20772 6381 20773
rect 6315 20708 6316 20772
rect 6380 20708 6381 20772
rect 6315 20707 6381 20708
rect 5395 19412 5461 19413
rect 5395 19348 5396 19412
rect 5460 19348 5461 19412
rect 5395 19347 5461 19348
rect 5211 19276 5277 19277
rect 5211 19212 5212 19276
rect 5276 19212 5277 19276
rect 5211 19211 5277 19212
rect 4279 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4599 18528
rect 4279 17440 4599 18464
rect 4279 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4599 17440
rect 4279 16352 4599 17376
rect 4279 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4599 16352
rect 4279 15264 4599 16288
rect 4279 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4599 15264
rect 4279 14176 4599 15200
rect 4279 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4599 14176
rect 4279 13088 4599 14112
rect 4279 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4599 13088
rect 4279 12000 4599 13024
rect 4279 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4599 12000
rect 4279 10912 4599 11936
rect 4279 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4599 10912
rect 4279 9824 4599 10848
rect 4279 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4599 9824
rect 4279 8736 4599 9760
rect 4279 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4599 8736
rect 4279 7648 4599 8672
rect 5398 7717 5458 19347
rect 5395 7716 5461 7717
rect 5395 7652 5396 7716
rect 5460 7652 5461 7716
rect 5395 7651 5461 7652
rect 4279 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4599 7648
rect 4279 6560 4599 7584
rect 6318 7581 6378 20707
rect 7974 20637 8034 22070
rect 9446 21858 9506 22174
rect 9630 22130 9690 22304
rect 9630 22070 9874 22130
rect 9627 21996 9693 21997
rect 9627 21932 9628 21996
rect 9692 21932 9693 21996
rect 9627 21931 9693 21932
rect 9630 21858 9690 21931
rect 8166 21248 8486 21808
rect 9446 21798 9690 21858
rect 9814 21450 9874 22070
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 7971 20636 8037 20637
rect 7971 20572 7972 20636
rect 8036 20572 8037 20636
rect 7971 20571 8037 20572
rect 8166 20160 8486 21184
rect 9630 21390 9874 21450
rect 9630 20637 9690 21390
rect 10366 21045 10426 22304
rect 10363 21044 10429 21045
rect 10363 20980 10364 21044
rect 10428 20980 10429 21044
rect 10363 20979 10429 20980
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 9627 20636 9693 20637
rect 9627 20572 9628 20636
rect 9692 20572 9693 20636
rect 9627 20571 9693 20572
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 10179 19684 10245 19685
rect 10179 19620 10180 19684
rect 10244 19620 10245 19684
rect 10179 19619 10245 19620
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 9811 18324 9877 18325
rect 9811 18260 9812 18324
rect 9876 18260 9877 18324
rect 9811 18259 9877 18260
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 9627 16828 9693 16829
rect 9627 16764 9628 16828
rect 9692 16764 9693 16828
rect 9627 16763 9693 16764
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 7971 15196 8037 15197
rect 7971 15132 7972 15196
rect 8036 15132 8037 15196
rect 7971 15131 8037 15132
rect 7051 10028 7117 10029
rect 7051 9964 7052 10028
rect 7116 9964 7117 10028
rect 7051 9963 7117 9964
rect 6867 7852 6933 7853
rect 6867 7788 6868 7852
rect 6932 7788 6933 7852
rect 6867 7787 6933 7788
rect 6315 7580 6381 7581
rect 6315 7516 6316 7580
rect 6380 7516 6381 7580
rect 6315 7515 6381 7516
rect 6318 6629 6378 7515
rect 6315 6628 6381 6629
rect 6315 6564 6316 6628
rect 6380 6564 6381 6628
rect 6315 6563 6381 6564
rect 4279 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4599 6560
rect 4279 5472 4599 6496
rect 6870 5677 6930 7787
rect 7054 5949 7114 9963
rect 7419 8396 7485 8397
rect 7419 8332 7420 8396
rect 7484 8332 7485 8396
rect 7419 8331 7485 8332
rect 7422 6085 7482 8331
rect 7974 7853 8034 15131
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8891 13972 8957 13973
rect 8891 13908 8892 13972
rect 8956 13908 8957 13972
rect 8891 13907 8957 13908
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8894 10981 8954 13907
rect 9630 13429 9690 16763
rect 9814 14925 9874 18259
rect 9811 14924 9877 14925
rect 9811 14860 9812 14924
rect 9876 14860 9877 14924
rect 9811 14859 9877 14860
rect 9627 13428 9693 13429
rect 9627 13364 9628 13428
rect 9692 13364 9693 13428
rect 9627 13363 9693 13364
rect 9627 12612 9693 12613
rect 9627 12548 9628 12612
rect 9692 12548 9693 12612
rect 9627 12547 9693 12548
rect 8891 10980 8957 10981
rect 8891 10916 8892 10980
rect 8956 10916 8957 10980
rect 8891 10915 8957 10916
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 9630 9349 9690 12547
rect 9627 9348 9693 9349
rect 9627 9284 9628 9348
rect 9692 9284 9693 9348
rect 9627 9283 9693 9284
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 9811 8940 9877 8941
rect 9811 8876 9812 8940
rect 9876 8876 9877 8940
rect 9811 8875 9877 8876
rect 9995 8940 10061 8941
rect 9995 8876 9996 8940
rect 10060 8876 10061 8940
rect 9995 8875 10061 8876
rect 9443 8804 9509 8805
rect 9443 8740 9444 8804
rect 9508 8740 9509 8804
rect 9443 8739 9509 8740
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 7971 7852 8037 7853
rect 7971 7788 7972 7852
rect 8036 7788 8037 7852
rect 7971 7787 8037 7788
rect 8166 7104 8486 8128
rect 8707 7852 8773 7853
rect 8707 7788 8708 7852
rect 8772 7788 8773 7852
rect 8707 7787 8773 7788
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 7419 6084 7485 6085
rect 7419 6020 7420 6084
rect 7484 6020 7485 6084
rect 7419 6019 7485 6020
rect 8166 6016 8486 7040
rect 8710 6765 8770 7787
rect 9446 7037 9506 8739
rect 9443 7036 9509 7037
rect 9443 6972 9444 7036
rect 9508 6972 9509 7036
rect 9443 6971 9509 6972
rect 8707 6764 8773 6765
rect 8707 6700 8708 6764
rect 8772 6700 8773 6764
rect 8707 6699 8773 6700
rect 9814 6085 9874 8875
rect 9998 8125 10058 8875
rect 10182 8261 10242 19619
rect 10731 17236 10797 17237
rect 10731 17172 10732 17236
rect 10796 17172 10797 17236
rect 10731 17171 10797 17172
rect 10734 10845 10794 17171
rect 10731 10844 10797 10845
rect 10731 10780 10732 10844
rect 10796 10780 10797 10844
rect 10731 10779 10797 10780
rect 10731 9212 10797 9213
rect 10731 9148 10732 9212
rect 10796 9148 10797 9212
rect 10731 9147 10797 9148
rect 10179 8260 10245 8261
rect 10179 8196 10180 8260
rect 10244 8196 10245 8260
rect 10179 8195 10245 8196
rect 9995 8124 10061 8125
rect 9995 8060 9996 8124
rect 10060 8060 10061 8124
rect 9995 8059 10061 8060
rect 10734 7717 10794 9147
rect 10731 7716 10797 7717
rect 10731 7652 10732 7716
rect 10796 7652 10797 7716
rect 10731 7651 10797 7652
rect 10547 7580 10613 7581
rect 10547 7516 10548 7580
rect 10612 7516 10613 7580
rect 10547 7515 10613 7516
rect 9811 6084 9877 6085
rect 9811 6020 9812 6084
rect 9876 6020 9877 6084
rect 9811 6019 9877 6020
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 7051 5948 7117 5949
rect 7051 5884 7052 5948
rect 7116 5884 7117 5948
rect 7051 5883 7117 5884
rect 6867 5676 6933 5677
rect 6867 5612 6868 5676
rect 6932 5612 6933 5676
rect 6867 5611 6933 5612
rect 4279 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4599 5472
rect 4279 4384 4599 5408
rect 4279 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4599 4384
rect 4279 3296 4599 4320
rect 4279 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4599 3296
rect 4279 2208 4599 3232
rect 4279 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4599 2208
rect 4279 1120 4599 2144
rect 4279 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4599 1120
rect 4279 496 4599 1056
rect 8166 4928 8486 5952
rect 10550 5133 10610 7515
rect 10918 7037 10978 20707
rect 11102 19277 11162 22304
rect 11838 20637 11898 22304
rect 12574 21861 12634 22304
rect 12571 21860 12637 21861
rect 12053 21792 12373 21808
rect 12571 21796 12572 21860
rect 12636 21796 12637 21860
rect 12571 21795 12637 21796
rect 12053 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12373 21792
rect 12053 20704 12373 21728
rect 13310 21725 13370 22304
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 14046 21589 14106 22304
rect 14782 22133 14842 22304
rect 14779 22132 14845 22133
rect 14779 22068 14780 22132
rect 14844 22068 14845 22132
rect 14779 22067 14845 22068
rect 14043 21588 14109 21589
rect 14043 21524 14044 21588
rect 14108 21524 14109 21588
rect 14043 21523 14109 21524
rect 15518 21453 15578 22304
rect 16254 21997 16314 22304
rect 16251 21996 16317 21997
rect 16251 21932 16252 21996
rect 16316 21932 16317 21996
rect 16251 21931 16317 21932
rect 15515 21452 15581 21453
rect 15515 21388 15516 21452
rect 15580 21388 15581 21452
rect 15515 21387 15581 21388
rect 15940 21248 16260 21808
rect 15940 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16260 21248
rect 12755 21044 12821 21045
rect 12755 20980 12756 21044
rect 12820 20980 12821 21044
rect 12755 20979 12821 20980
rect 12053 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12373 20704
rect 11835 20636 11901 20637
rect 11835 20572 11836 20636
rect 11900 20572 11901 20636
rect 11835 20571 11901 20572
rect 12053 19616 12373 20640
rect 12053 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12373 19616
rect 11099 19276 11165 19277
rect 11099 19212 11100 19276
rect 11164 19212 11165 19276
rect 11099 19211 11165 19212
rect 11835 18868 11901 18869
rect 11835 18804 11836 18868
rect 11900 18804 11901 18868
rect 11835 18803 11901 18804
rect 11838 9485 11898 18803
rect 12053 18528 12373 19552
rect 12053 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12373 18528
rect 12053 17440 12373 18464
rect 12053 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12373 17440
rect 12053 16352 12373 17376
rect 12053 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12373 16352
rect 12053 15264 12373 16288
rect 12053 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12373 15264
rect 12053 14176 12373 15200
rect 12053 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12373 14176
rect 12053 13088 12373 14112
rect 12053 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12373 13088
rect 12053 12000 12373 13024
rect 12053 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12373 12000
rect 12053 10912 12373 11936
rect 12053 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12373 10912
rect 12053 9824 12373 10848
rect 12053 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12373 9824
rect 11835 9484 11901 9485
rect 11835 9420 11836 9484
rect 11900 9420 11901 9484
rect 11835 9419 11901 9420
rect 11838 7717 11898 9419
rect 12053 8736 12373 9760
rect 12053 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12373 8736
rect 11835 7716 11901 7717
rect 11835 7652 11836 7716
rect 11900 7652 11901 7716
rect 11835 7651 11901 7652
rect 12053 7648 12373 8672
rect 12758 8533 12818 20979
rect 15940 20160 16260 21184
rect 16990 20637 17050 22304
rect 17726 21589 17786 22304
rect 18462 22104 18522 22304
rect 19198 22104 19258 22304
rect 19934 22104 19994 22304
rect 20670 22104 20730 22304
rect 21406 22104 21466 22304
rect 22142 22104 22202 22304
rect 22878 22104 22938 22304
rect 23614 22104 23674 22304
rect 24350 21861 24410 22304
rect 25086 21997 25146 22304
rect 25083 21996 25149 21997
rect 25083 21932 25084 21996
rect 25148 21932 25149 21996
rect 25083 21931 25149 21932
rect 25822 21861 25882 22304
rect 24347 21860 24413 21861
rect 19827 21792 20147 21808
rect 19827 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20147 21792
rect 17723 21588 17789 21589
rect 17723 21524 17724 21588
rect 17788 21524 17789 21588
rect 17723 21523 17789 21524
rect 19379 21044 19445 21045
rect 19379 20980 19380 21044
rect 19444 20980 19445 21044
rect 19379 20979 19445 20980
rect 16987 20636 17053 20637
rect 16987 20572 16988 20636
rect 17052 20572 17053 20636
rect 16987 20571 17053 20572
rect 17723 20364 17789 20365
rect 17723 20300 17724 20364
rect 17788 20300 17789 20364
rect 17723 20299 17789 20300
rect 15940 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16260 20160
rect 13491 19412 13557 19413
rect 13491 19348 13492 19412
rect 13556 19348 13557 19412
rect 13491 19347 13557 19348
rect 13494 16421 13554 19347
rect 15940 19072 16260 20096
rect 15940 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16260 19072
rect 15940 17984 16260 19008
rect 16803 19004 16869 19005
rect 16803 18940 16804 19004
rect 16868 18940 16869 19004
rect 16803 18939 16869 18940
rect 15940 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16260 17984
rect 15940 16896 16260 17920
rect 15940 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16260 16896
rect 13491 16420 13557 16421
rect 13491 16356 13492 16420
rect 13556 16356 13557 16420
rect 13491 16355 13557 16356
rect 15940 15808 16260 16832
rect 15940 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16260 15808
rect 15940 14720 16260 15744
rect 16806 15333 16866 18939
rect 17171 17372 17237 17373
rect 17171 17308 17172 17372
rect 17236 17308 17237 17372
rect 17171 17307 17237 17308
rect 16803 15332 16869 15333
rect 16803 15268 16804 15332
rect 16868 15268 16869 15332
rect 16803 15267 16869 15268
rect 15940 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16260 14720
rect 15940 13632 16260 14656
rect 17174 14109 17234 17307
rect 17171 14108 17237 14109
rect 17171 14044 17172 14108
rect 17236 14044 17237 14108
rect 17171 14043 17237 14044
rect 17726 13701 17786 20299
rect 18275 18188 18341 18189
rect 18275 18124 18276 18188
rect 18340 18124 18341 18188
rect 18275 18123 18341 18124
rect 18278 14653 18338 18123
rect 18643 18052 18709 18053
rect 18643 17988 18644 18052
rect 18708 17988 18709 18052
rect 18643 17987 18709 17988
rect 18646 14789 18706 17987
rect 19382 17370 19442 20979
rect 19827 20704 20147 21728
rect 19827 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20147 20704
rect 19827 19616 20147 20640
rect 19827 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20147 19616
rect 19827 18528 20147 19552
rect 23714 21248 24034 21808
rect 24347 21796 24348 21860
rect 24412 21796 24413 21860
rect 24347 21795 24413 21796
rect 25819 21860 25885 21861
rect 25819 21796 25820 21860
rect 25884 21796 25885 21860
rect 25819 21795 25885 21796
rect 26558 21725 26618 22304
rect 26555 21724 26621 21725
rect 26555 21660 26556 21724
rect 26620 21660 26621 21724
rect 26555 21659 26621 21660
rect 27294 21589 27354 22304
rect 28030 21861 28090 22304
rect 28766 21997 28826 22304
rect 28763 21996 28829 21997
rect 28763 21932 28764 21996
rect 28828 21932 28829 21996
rect 28763 21931 28829 21932
rect 29502 21861 29562 22304
rect 30238 21861 30298 22304
rect 28027 21860 28093 21861
rect 27601 21792 27921 21808
rect 28027 21796 28028 21860
rect 28092 21796 28093 21860
rect 28027 21795 28093 21796
rect 29499 21860 29565 21861
rect 29499 21796 29500 21860
rect 29564 21796 29565 21860
rect 29499 21795 29565 21796
rect 30235 21860 30301 21861
rect 30235 21796 30236 21860
rect 30300 21796 30301 21860
rect 30235 21795 30301 21796
rect 27601 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27921 21792
rect 27291 21588 27357 21589
rect 27291 21524 27292 21588
rect 27356 21524 27357 21588
rect 27291 21523 27357 21524
rect 23714 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24034 21248
rect 23714 20160 24034 21184
rect 23714 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24034 20160
rect 21403 19548 21469 19549
rect 21403 19484 21404 19548
rect 21468 19484 21469 19548
rect 21403 19483 21469 19484
rect 21955 19548 22021 19549
rect 21955 19484 21956 19548
rect 22020 19484 22021 19548
rect 21955 19483 22021 19484
rect 23427 19548 23493 19549
rect 23427 19484 23428 19548
rect 23492 19484 23493 19548
rect 23427 19483 23493 19484
rect 20483 19004 20549 19005
rect 20483 18940 20484 19004
rect 20548 18940 20549 19004
rect 20483 18939 20549 18940
rect 19827 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20147 18528
rect 19827 17440 20147 18464
rect 19827 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20147 17440
rect 19382 17310 19626 17370
rect 19566 17237 19626 17310
rect 19563 17236 19629 17237
rect 19563 17172 19564 17236
rect 19628 17172 19629 17236
rect 19563 17171 19629 17172
rect 18827 16284 18893 16285
rect 18827 16220 18828 16284
rect 18892 16220 18893 16284
rect 18827 16219 18893 16220
rect 18830 15333 18890 16219
rect 18827 15332 18893 15333
rect 18827 15268 18828 15332
rect 18892 15268 18893 15332
rect 18827 15267 18893 15268
rect 19566 15061 19626 17171
rect 19827 16352 20147 17376
rect 19827 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20147 16352
rect 19827 15264 20147 16288
rect 19827 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20147 15264
rect 19563 15060 19629 15061
rect 19563 14996 19564 15060
rect 19628 14996 19629 15060
rect 19563 14995 19629 14996
rect 18643 14788 18709 14789
rect 18643 14724 18644 14788
rect 18708 14724 18709 14788
rect 18643 14723 18709 14724
rect 18275 14652 18341 14653
rect 18275 14588 18276 14652
rect 18340 14588 18341 14652
rect 18275 14587 18341 14588
rect 19827 14176 20147 15200
rect 19827 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20147 14176
rect 17723 13700 17789 13701
rect 17723 13636 17724 13700
rect 17788 13636 17789 13700
rect 17723 13635 17789 13636
rect 15940 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16260 13632
rect 15940 12544 16260 13568
rect 15940 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16260 12544
rect 15940 11456 16260 12480
rect 15940 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16260 11456
rect 15940 10368 16260 11392
rect 15940 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16260 10368
rect 15940 9280 16260 10304
rect 15940 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16260 9280
rect 12755 8532 12821 8533
rect 12755 8468 12756 8532
rect 12820 8468 12821 8532
rect 12755 8467 12821 8468
rect 12758 8261 12818 8467
rect 12755 8260 12821 8261
rect 12755 8196 12756 8260
rect 12820 8196 12821 8260
rect 12755 8195 12821 8196
rect 12053 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12373 7648
rect 10915 7036 10981 7037
rect 10915 6972 10916 7036
rect 10980 6972 10981 7036
rect 10915 6971 10981 6972
rect 12053 6560 12373 7584
rect 12053 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12373 6560
rect 12053 5472 12373 6496
rect 12053 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12373 5472
rect 10547 5132 10613 5133
rect 10547 5068 10548 5132
rect 10612 5068 10613 5132
rect 10547 5067 10613 5068
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 1664 8486 2688
rect 8166 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8486 1664
rect 8166 576 8486 1600
rect 8166 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8486 576
rect 8166 496 8486 512
rect 12053 4384 12373 5408
rect 12053 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12373 4384
rect 12053 3296 12373 4320
rect 12053 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12373 3296
rect 12053 2208 12373 3232
rect 12053 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12373 2208
rect 12053 1120 12373 2144
rect 12053 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12373 1120
rect 12053 496 12373 1056
rect 15940 8192 16260 9216
rect 15940 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16260 8192
rect 15940 7104 16260 8128
rect 15940 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16260 7104
rect 15940 6016 16260 7040
rect 15940 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16260 6016
rect 15940 4928 16260 5952
rect 15940 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16260 4928
rect 15940 3840 16260 4864
rect 15940 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16260 3840
rect 15940 2752 16260 3776
rect 15940 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16260 2752
rect 15940 1664 16260 2688
rect 15940 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16260 1664
rect 15940 576 16260 1600
rect 15940 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16260 576
rect 15940 496 16260 512
rect 19827 13088 20147 14112
rect 19827 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20147 13088
rect 19827 12000 20147 13024
rect 19827 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20147 12000
rect 19827 10912 20147 11936
rect 19827 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20147 10912
rect 19827 9824 20147 10848
rect 19827 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20147 9824
rect 19827 8736 20147 9760
rect 20486 9621 20546 18939
rect 21406 16557 21466 19483
rect 21403 16556 21469 16557
rect 21403 16492 21404 16556
rect 21468 16492 21469 16556
rect 21403 16491 21469 16492
rect 21958 15061 22018 19483
rect 23430 15605 23490 19483
rect 23714 19072 24034 20096
rect 27601 20704 27921 21728
rect 30051 20772 30117 20773
rect 30051 20708 30052 20772
rect 30116 20708 30117 20772
rect 30051 20707 30117 20708
rect 27601 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27921 20704
rect 27601 19616 27921 20640
rect 27601 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27921 19616
rect 27107 19412 27173 19413
rect 27107 19348 27108 19412
rect 27172 19348 27173 19412
rect 27107 19347 27173 19348
rect 23714 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24034 19072
rect 23714 17984 24034 19008
rect 23714 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24034 17984
rect 23714 16896 24034 17920
rect 23714 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24034 16896
rect 23714 15808 24034 16832
rect 23714 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24034 15808
rect 23427 15604 23493 15605
rect 23427 15540 23428 15604
rect 23492 15540 23493 15604
rect 23427 15539 23493 15540
rect 21955 15060 22021 15061
rect 21955 14996 21956 15060
rect 22020 14996 22021 15060
rect 21955 14995 22021 14996
rect 23714 14720 24034 15744
rect 23714 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24034 14720
rect 23714 13632 24034 14656
rect 23714 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24034 13632
rect 23714 12544 24034 13568
rect 23714 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24034 12544
rect 23714 11456 24034 12480
rect 23714 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24034 11456
rect 23714 10368 24034 11392
rect 23714 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24034 10368
rect 20483 9620 20549 9621
rect 20483 9556 20484 9620
rect 20548 9556 20549 9620
rect 20483 9555 20549 9556
rect 19827 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20147 8736
rect 19827 7648 20147 8672
rect 19827 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20147 7648
rect 19827 6560 20147 7584
rect 19827 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20147 6560
rect 19827 5472 20147 6496
rect 19827 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20147 5472
rect 19827 4384 20147 5408
rect 19827 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20147 4384
rect 19827 3296 20147 4320
rect 19827 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20147 3296
rect 19827 2208 20147 3232
rect 19827 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20147 2208
rect 19827 1120 20147 2144
rect 19827 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20147 1120
rect 19827 496 20147 1056
rect 23714 9280 24034 10304
rect 27110 10029 27170 19347
rect 27601 18528 27921 19552
rect 27601 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27921 18528
rect 27601 17440 27921 18464
rect 27601 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27921 17440
rect 27601 16352 27921 17376
rect 27601 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27921 16352
rect 27601 15264 27921 16288
rect 27601 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27921 15264
rect 27601 14176 27921 15200
rect 27601 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27921 14176
rect 27601 13088 27921 14112
rect 27601 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27921 13088
rect 27601 12000 27921 13024
rect 27601 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27921 12000
rect 27601 10912 27921 11936
rect 30054 11797 30114 20707
rect 30974 16013 31034 22304
rect 31710 22104 31770 22304
rect 31488 21248 31808 21808
rect 31488 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31808 21248
rect 31488 20160 31808 21184
rect 31488 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31808 20160
rect 31488 19072 31808 20096
rect 31488 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31808 19072
rect 31488 17984 31808 19008
rect 31488 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31808 17984
rect 31488 16896 31808 17920
rect 31488 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31808 16896
rect 30971 16012 31037 16013
rect 30971 15948 30972 16012
rect 31036 15948 31037 16012
rect 30971 15947 31037 15948
rect 31488 15808 31808 16832
rect 31488 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31808 15808
rect 31488 14720 31808 15744
rect 31488 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31808 14720
rect 31488 13632 31808 14656
rect 31488 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31808 13632
rect 31488 12544 31808 13568
rect 31488 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31808 12544
rect 30051 11796 30117 11797
rect 30051 11732 30052 11796
rect 30116 11732 30117 11796
rect 30051 11731 30117 11732
rect 27601 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27921 10912
rect 27107 10028 27173 10029
rect 27107 9964 27108 10028
rect 27172 9964 27173 10028
rect 27107 9963 27173 9964
rect 23714 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24034 9280
rect 23714 8192 24034 9216
rect 23714 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24034 8192
rect 23714 7104 24034 8128
rect 23714 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24034 7104
rect 23714 6016 24034 7040
rect 23714 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24034 6016
rect 23714 4928 24034 5952
rect 23714 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24034 4928
rect 23714 3840 24034 4864
rect 23714 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24034 3840
rect 23714 2752 24034 3776
rect 23714 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24034 2752
rect 23714 1664 24034 2688
rect 23714 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24034 1664
rect 23714 576 24034 1600
rect 23714 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24034 576
rect 23714 496 24034 512
rect 27601 9824 27921 10848
rect 27601 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27921 9824
rect 27601 8736 27921 9760
rect 27601 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27921 8736
rect 27601 7648 27921 8672
rect 27601 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27921 7648
rect 27601 6560 27921 7584
rect 27601 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27921 6560
rect 27601 5472 27921 6496
rect 27601 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27921 5472
rect 27601 4384 27921 5408
rect 27601 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27921 4384
rect 27601 3296 27921 4320
rect 27601 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27921 3296
rect 27601 2208 27921 3232
rect 27601 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27921 2208
rect 27601 1120 27921 2144
rect 27601 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27921 1120
rect 27601 496 27921 1056
rect 31488 11456 31808 12480
rect 31488 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31808 11456
rect 31488 10368 31808 11392
rect 31488 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31808 10368
rect 31488 9280 31808 10304
rect 31488 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31808 9280
rect 31488 8192 31808 9216
rect 31488 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31808 8192
rect 31488 7104 31808 8128
rect 31488 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31808 7104
rect 31488 6016 31808 7040
rect 31488 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31808 6016
rect 31488 4928 31808 5952
rect 31488 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31808 4928
rect 31488 3840 31808 4864
rect 31488 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31808 3840
rect 31488 2752 31808 3776
rect 31488 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31808 2752
rect 31488 1664 31808 2688
rect 31488 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31808 1664
rect 31488 576 31808 1600
rect 31488 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31808 576
rect 31488 496 31808 512
use sky130_fd_sc_hd__inv_2  _0922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21160 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16284 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0926_
timestamp 1704896540
transform 1 0 16560 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15548 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16744 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17756 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0930_
timestamp 1704896540
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0932_
timestamp 1704896540
transform 1 0 19780 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8280 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20148 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1704896540
transform -1 0 18584 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27416 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27416 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 1704896540
transform -1 0 14352 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0939_
timestamp 1704896540
transform 1 0 14628 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1704896540
transform -1 0 12052 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0941_
timestamp 1704896540
transform 1 0 11776 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1704896540
transform -1 0 7452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0944_
timestamp 1704896540
transform -1 0 8280 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1704896540
transform -1 0 5796 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1704896540
transform 1 0 11408 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0947_
timestamp 1704896540
transform -1 0 11592 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1704896540
transform -1 0 8188 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1704896540
transform -1 0 10120 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0950_
timestamp 1704896540
transform 1 0 9752 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 1704896540
transform 1 0 8464 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1704896540
transform -1 0 9200 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0953_
timestamp 1704896540
transform 1 0 9200 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1704896540
transform 1 0 4784 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1704896540
transform -1 0 5336 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0956_
timestamp 1704896540
transform 1 0 6072 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp 1704896540
transform -1 0 5704 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 1704896540
transform -1 0 6164 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0959_
timestamp 1704896540
transform 1 0 8372 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0960_
timestamp 1704896540
transform -1 0 18216 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0961_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17664 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0963_
timestamp 1704896540
transform 1 0 15180 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0964_
timestamp 1704896540
transform 1 0 15640 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1704896540
transform -1 0 4968 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0967_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1704896540
transform -1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0969_
timestamp 1704896540
transform -1 0 9108 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10028 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_2  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7544 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0974_
timestamp 1704896540
transform 1 0 9936 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0975_
timestamp 1704896540
transform -1 0 11500 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0976_
timestamp 1704896540
transform -1 0 10764 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0977_
timestamp 1704896540
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0979_
timestamp 1704896540
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9568 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0981_
timestamp 1704896540
transform -1 0 28520 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21252 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24472 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0984_
timestamp 1704896540
transform -1 0 12788 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1704896540
transform -1 0 21160 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20332 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0987_
timestamp 1704896540
transform 1 0 22540 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16560 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1704896540
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0991_
timestamp 1704896540
transform -1 0 11316 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0992_
timestamp 1704896540
transform 1 0 5152 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0993_
timestamp 1704896540
transform 1 0 5796 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0994_
timestamp 1704896540
transform 1 0 6808 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _0996_
timestamp 1704896540
transform 1 0 6440 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1704896540
transform -1 0 21528 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _0998_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26956 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1704896540
transform -1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1002_
timestamp 1704896540
transform 1 0 23828 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1003_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25116 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1704896540
transform 1 0 10948 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1005_
timestamp 1704896540
transform -1 0 10948 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1006_
timestamp 1704896540
transform -1 0 6440 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1704896540
transform 1 0 4692 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1008_
timestamp 1704896540
transform 1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1009_
timestamp 1704896540
transform 1 0 920 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1010_
timestamp 1704896540
transform 1 0 1012 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1011_
timestamp 1704896540
transform 1 0 10304 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1704896540
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20608 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1014_
timestamp 1704896540
transform 1 0 24380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1015_
timestamp 1704896540
transform -1 0 24380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1704896540
transform -1 0 15180 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1017_
timestamp 1704896540
transform -1 0 22816 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1018_
timestamp 1704896540
transform -1 0 22356 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1019_
timestamp 1704896540
transform 1 0 25392 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1020_
timestamp 1704896540
transform 1 0 30452 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1704896540
transform 1 0 10948 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1022_
timestamp 1704896540
transform -1 0 10856 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1023_
timestamp 1704896540
transform -1 0 10028 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1024_
timestamp 1704896540
transform 1 0 8832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1025_
timestamp 1704896540
transform 1 0 7636 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1026_
timestamp 1704896540
transform -1 0 8280 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1027_
timestamp 1704896540
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1028_
timestamp 1704896540
transform -1 0 15732 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1704896540
transform -1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1030_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15732 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1032_
timestamp 1704896540
transform 1 0 30176 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1033_
timestamp 1704896540
transform -1 0 12420 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp 1704896540
transform 1 0 10028 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1035_
timestamp 1704896540
transform -1 0 8924 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1036_
timestamp 1704896540
transform -1 0 8832 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1037_
timestamp 1704896540
transform -1 0 8280 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1038_
timestamp 1704896540
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1039_
timestamp 1704896540
transform 1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1040_
timestamp 1704896540
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1041_
timestamp 1704896540
transform -1 0 16744 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1704896540
transform -1 0 13248 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1043_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1044_
timestamp 1704896540
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1045_
timestamp 1704896540
transform 1 0 17204 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1046_
timestamp 1704896540
transform 1 0 28980 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1047_
timestamp 1704896540
transform 1 0 29624 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1704896540
transform -1 0 10580 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1049_
timestamp 1704896540
transform 1 0 12328 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1050_
timestamp 1704896540
transform -1 0 5336 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1051_
timestamp 1704896540
transform 1 0 4508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1704896540
transform 1 0 4048 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1053_
timestamp 1704896540
transform -1 0 4784 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1054_
timestamp 1704896540
transform 1 0 4968 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_4  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15088 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 1704896540
transform -1 0 6624 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16100 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1704896540
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1704896540
transform 1 0 14720 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1060_
timestamp 1704896540
transform 1 0 15732 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1061_
timestamp 1704896540
transform 1 0 25024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1062_
timestamp 1704896540
transform 1 0 8924 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1063_
timestamp 1704896540
transform -1 0 8280 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1064_
timestamp 1704896540
transform 1 0 3772 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1065_
timestamp 1704896540
transform 1 0 4784 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1066_
timestamp 1704896540
transform 1 0 3404 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1067_
timestamp 1704896540
transform -1 0 4692 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1068_
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 1704896540
transform -1 0 5244 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10856 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12788 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1072_
timestamp 1704896540
transform 1 0 13248 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1073_
timestamp 1704896540
transform -1 0 10028 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1074_
timestamp 1704896540
transform 1 0 10028 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1075_
timestamp 1704896540
transform 1 0 3772 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1076_
timestamp 1704896540
transform 1 0 4416 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1077_
timestamp 1704896540
transform -1 0 2208 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1078_
timestamp 1704896540
transform -1 0 1932 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1079_
timestamp 1704896540
transform 1 0 4968 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1080_
timestamp 1704896540
transform -1 0 5244 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1081_
timestamp 1704896540
transform 1 0 11040 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _1082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1083_
timestamp 1704896540
transform 1 0 9200 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1084_
timestamp 1704896540
transform -1 0 7452 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1085_
timestamp 1704896540
transform -1 0 3312 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _1087_
timestamp 1704896540
transform 1 0 14076 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1088_
timestamp 1704896540
transform 1 0 13524 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1089_
timestamp 1704896540
transform 1 0 13524 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1090_
timestamp 1704896540
transform -1 0 14628 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1704896540
transform -1 0 13340 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1092_
timestamp 1704896540
transform 1 0 14628 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1093_
timestamp 1704896540
transform -1 0 23276 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1094_
timestamp 1704896540
transform 1 0 23828 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1095_
timestamp 1704896540
transform 1 0 24656 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1704896540
transform 1 0 23552 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19964 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1098_
timestamp 1704896540
transform 1 0 24012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1099_
timestamp 1704896540
transform -1 0 25116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21252 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21068 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1103_
timestamp 1704896540
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_4  _1104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _1105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23644 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _1106_
timestamp 1704896540
transform -1 0 20792 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1107_
timestamp 1704896540
transform 1 0 24748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1108_
timestamp 1704896540
transform -1 0 30912 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1109_
timestamp 1704896540
transform -1 0 28520 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_
timestamp 1704896540
transform 1 0 17848 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1111_
timestamp 1704896540
transform 1 0 19412 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1112_
timestamp 1704896540
transform 1 0 27968 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22080 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1114_
timestamp 1704896540
transform -1 0 20608 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1115_
timestamp 1704896540
transform 1 0 18492 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1116_
timestamp 1704896540
transform 1 0 20516 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1117_
timestamp 1704896540
transform 1 0 23828 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1118_
timestamp 1704896540
transform 1 0 19964 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1704896540
transform 1 0 27876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1121_
timestamp 1704896540
transform -1 0 25392 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1122_
timestamp 1704896540
transform -1 0 27876 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13432 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1124_
timestamp 1704896540
transform -1 0 13984 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _1125_
timestamp 1704896540
transform -1 0 25484 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1704896540
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1127_
timestamp 1704896540
transform -1 0 28060 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1704896540
transform -1 0 16376 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1129_
timestamp 1704896540
transform 1 0 16284 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1130_
timestamp 1704896540
transform 1 0 30636 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1131_
timestamp 1704896540
transform -1 0 25852 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1132_
timestamp 1704896540
transform -1 0 26312 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _1133_
timestamp 1704896540
transform 1 0 19964 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_4  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1704896540
transform -1 0 25852 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1136_
timestamp 1704896540
transform -1 0 24748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1137_
timestamp 1704896540
transform 1 0 27416 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _1138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25852 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1704896540
transform -1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27692 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1141_
timestamp 1704896540
transform 1 0 27416 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1142_
timestamp 1704896540
transform -1 0 21068 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1143_
timestamp 1704896540
transform -1 0 23368 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1144_
timestamp 1704896540
transform 1 0 20516 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_2  _1145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19872 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _1147_
timestamp 1704896540
transform 1 0 19412 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1148_
timestamp 1704896540
transform 1 0 20056 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16008 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21436 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1151_
timestamp 1704896540
transform -1 0 21344 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26588 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1153_
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1154_
timestamp 1704896540
transform -1 0 22632 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1156_
timestamp 1704896540
transform 1 0 17940 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1157_
timestamp 1704896540
transform 1 0 17572 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1158_
timestamp 1704896540
transform 1 0 23092 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1704896540
transform 1 0 23644 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1160_
timestamp 1704896540
transform 1 0 24288 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1161_
timestamp 1704896540
transform -1 0 25024 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _1162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13984 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _1163_
timestamp 1704896540
transform 1 0 24104 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1164_
timestamp 1704896540
transform -1 0 19228 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1165_
timestamp 1704896540
transform 1 0 18768 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 1704896540
transform 1 0 19228 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22632 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1168_
timestamp 1704896540
transform -1 0 25392 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15916 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_1  _1170_
timestamp 1704896540
transform 1 0 26128 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1704896540
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1172_
timestamp 1704896540
transform -1 0 25484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1173_
timestamp 1704896540
transform -1 0 30728 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1174_
timestamp 1704896540
transform 1 0 21896 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27140 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1176_
timestamp 1704896540
transform 1 0 26680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1177_
timestamp 1704896540
transform 1 0 26680 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27140 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1179_
timestamp 1704896540
transform 1 0 26864 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_2  _1180_
timestamp 1704896540
transform 1 0 22172 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1704896540
transform 1 0 22816 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1182_
timestamp 1704896540
transform 1 0 23828 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1183_
timestamp 1704896540
transform 1 0 22080 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24380 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 1704896540
transform 1 0 22356 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1186_
timestamp 1704896540
transform -1 0 23552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1704896540
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1188_
timestamp 1704896540
transform 1 0 17020 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1189_
timestamp 1704896540
transform 1 0 29716 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1190_
timestamp 1704896540
transform 1 0 30452 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17664 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 28244 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1193_
timestamp 1704896540
transform 1 0 28428 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1194_
timestamp 1704896540
transform -1 0 24840 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1195_
timestamp 1704896540
transform -1 0 27140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_4  _1196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28520 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_1  _1197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25392 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1198_
timestamp 1704896540
transform 1 0 24196 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1199_
timestamp 1704896540
transform -1 0 25668 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1200_
timestamp 1704896540
transform 1 0 29900 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20516 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1202_
timestamp 1704896540
transform -1 0 25208 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1203_
timestamp 1704896540
transform 1 0 28060 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1204_
timestamp 1704896540
transform 1 0 29992 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28980 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 1704896540
transform 1 0 26772 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1207_
timestamp 1704896540
transform -1 0 28612 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1208_
timestamp 1704896540
transform 1 0 23828 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1209_
timestamp 1704896540
transform 1 0 23828 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1210_
timestamp 1704896540
transform -1 0 26312 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26588 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1212_
timestamp 1704896540
transform 1 0 27416 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1213_
timestamp 1704896540
transform 1 0 26956 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1214_
timestamp 1704896540
transform 1 0 25208 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1215_
timestamp 1704896540
transform -1 0 23276 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1704896540
transform -1 0 25300 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1217_
timestamp 1704896540
transform 1 0 25208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1704896540
transform 1 0 25668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1219_
timestamp 1704896540
transform -1 0 24564 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1220_
timestamp 1704896540
transform -1 0 25484 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23184 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1222_
timestamp 1704896540
transform 1 0 28060 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1223_
timestamp 1704896540
transform -1 0 29532 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1224_
timestamp 1704896540
transform -1 0 28888 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _1225_
timestamp 1704896540
transform -1 0 21344 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1704896540
transform 1 0 26404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23276 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1704896540
transform -1 0 23736 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23460 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1230_
timestamp 1704896540
transform -1 0 26312 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26680 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1232_
timestamp 1704896540
transform 1 0 26404 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21160 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1234_
timestamp 1704896540
transform -1 0 24288 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28152 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1236_
timestamp 1704896540
transform 1 0 29440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1237_
timestamp 1704896540
transform -1 0 29440 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1238_
timestamp 1704896540
transform -1 0 29716 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1239_
timestamp 1704896540
transform -1 0 28520 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1240_
timestamp 1704896540
transform -1 0 27508 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1704896540
transform 1 0 28612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_4  _1242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 28152 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__a221o_1  _1243_
timestamp 1704896540
transform 1 0 25024 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1244_
timestamp 1704896540
transform 1 0 26404 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1245_
timestamp 1704896540
transform -1 0 28060 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1246_
timestamp 1704896540
transform 1 0 24380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24932 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 1704896540
transform 1 0 22172 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1250_
timestamp 1704896540
transform 1 0 22540 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _1251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23276 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _1252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 1 5984
box -38 -48 1418 592
use sky130_fd_sc_hd__o211a_1  _1253_
timestamp 1704896540
transform -1 0 23644 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24288 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1255_
timestamp 1704896540
transform 1 0 18400 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14260 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1257_
timestamp 1704896540
transform 1 0 14352 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1258_
timestamp 1704896540
transform -1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1704896540
transform -1 0 13800 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_4  _1260_
timestamp 1704896540
transform 1 0 26680 0 1 5984
box -38 -48 1418 592
use sky130_fd_sc_hd__a21o_1  _1261_
timestamp 1704896540
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1262_
timestamp 1704896540
transform 1 0 24564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1263_
timestamp 1704896540
transform -1 0 24564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _1264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21252 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1265_
timestamp 1704896540
transform 1 0 23828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _1266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21620 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21160 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1268_
timestamp 1704896540
transform 1 0 16192 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1704896540
transform -1 0 17848 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1270_
timestamp 1704896540
transform -1 0 17756 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 1704896540
transform -1 0 8924 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1272_
timestamp 1704896540
transform 1 0 8280 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1273_
timestamp 1704896540
transform -1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1274_
timestamp 1704896540
transform 1 0 11592 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1275_
timestamp 1704896540
transform -1 0 21068 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1276_
timestamp 1704896540
transform -1 0 25116 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1277_
timestamp 1704896540
transform 1 0 19504 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19412 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1279_
timestamp 1704896540
transform -1 0 19504 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1280_
timestamp 1704896540
transform -1 0 15640 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1281_
timestamp 1704896540
transform 1 0 20424 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1282_
timestamp 1704896540
transform 1 0 16928 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1283_
timestamp 1704896540
transform 1 0 22172 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1284_
timestamp 1704896540
transform -1 0 17020 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1285_
timestamp 1704896540
transform 1 0 17020 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1286_
timestamp 1704896540
transform 1 0 16836 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1287_
timestamp 1704896540
transform 1 0 13524 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1288_
timestamp 1704896540
transform 1 0 17756 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1704896540
transform -1 0 17020 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1290_
timestamp 1704896540
transform -1 0 18124 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1291_
timestamp 1704896540
transform 1 0 17020 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1292_
timestamp 1704896540
transform -1 0 17664 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1704896540
transform -1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1294_
timestamp 1704896540
transform 1 0 25116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1295_
timestamp 1704896540
transform -1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1296_
timestamp 1704896540
transform 1 0 28888 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1297_
timestamp 1704896540
transform -1 0 17664 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1298_
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1299_
timestamp 1704896540
transform 1 0 28336 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1300_
timestamp 1704896540
transform -1 0 31096 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1301_
timestamp 1704896540
transform -1 0 16652 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1302_
timestamp 1704896540
transform -1 0 29440 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1303_
timestamp 1704896540
transform 1 0 30268 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1304_
timestamp 1704896540
transform 1 0 30636 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1305_
timestamp 1704896540
transform -1 0 31280 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1306_
timestamp 1704896540
transform 1 0 30084 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1307_
timestamp 1704896540
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1308_
timestamp 1704896540
transform 1 0 28980 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1309_
timestamp 1704896540
transform 1 0 28980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _1310_
timestamp 1704896540
transform -1 0 27600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1311_
timestamp 1704896540
transform -1 0 23552 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1704896540
transform 1 0 27784 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27784 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _1314_
timestamp 1704896540
transform 1 0 25300 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25208 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1316_
timestamp 1704896540
transform 1 0 22356 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1317_
timestamp 1704896540
transform -1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1318_
timestamp 1704896540
transform -1 0 24472 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1319_
timestamp 1704896540
transform 1 0 26404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1320_
timestamp 1704896540
transform 1 0 27508 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1321_
timestamp 1704896540
transform 1 0 26864 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1322_
timestamp 1704896540
transform 1 0 26036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1323_
timestamp 1704896540
transform -1 0 25760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1324_
timestamp 1704896540
transform -1 0 27692 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1325_
timestamp 1704896540
transform -1 0 27048 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1326_
timestamp 1704896540
transform -1 0 26312 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1327_
timestamp 1704896540
transform 1 0 27692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23736 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _1329_
timestamp 1704896540
transform 1 0 13340 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1330_
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1704896540
transform -1 0 8280 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1332_
timestamp 1704896540
transform 1 0 20700 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1333_
timestamp 1704896540
transform -1 0 18216 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1334_
timestamp 1704896540
transform 1 0 20332 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1704896540
transform -1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1336_
timestamp 1704896540
transform 1 0 18124 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _1337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18860 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1338_
timestamp 1704896540
transform -1 0 18860 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1339_
timestamp 1704896540
transform -1 0 17480 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1340_
timestamp 1704896540
transform 1 0 16836 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1341_
timestamp 1704896540
transform -1 0 17940 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1704896540
transform -1 0 19412 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1343_
timestamp 1704896540
transform 1 0 21252 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1704896540
transform -1 0 14352 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1345_
timestamp 1704896540
transform 1 0 14352 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1704896540
transform 1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1347_
timestamp 1704896540
transform 1 0 12696 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1348_
timestamp 1704896540
transform 1 0 12512 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1704896540
transform 1 0 22724 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1350_
timestamp 1704896540
transform 1 0 16468 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1351_
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1352_
timestamp 1704896540
transform -1 0 13432 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1353_
timestamp 1704896540
transform 1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1354_
timestamp 1704896540
transform -1 0 12328 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1355_
timestamp 1704896540
transform -1 0 13248 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1356_
timestamp 1704896540
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1357_
timestamp 1704896540
transform -1 0 27232 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1358_
timestamp 1704896540
transform 1 0 21068 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1359_
timestamp 1704896540
transform 1 0 20424 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1360_
timestamp 1704896540
transform -1 0 22080 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _1361_
timestamp 1704896540
transform -1 0 16008 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _1362_
timestamp 1704896540
transform 1 0 24288 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1364_
timestamp 1704896540
transform -1 0 25024 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1365_
timestamp 1704896540
transform 1 0 25392 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1366_
timestamp 1704896540
transform 1 0 26404 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1367_
timestamp 1704896540
transform 1 0 26956 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1368_
timestamp 1704896540
transform -1 0 27600 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1369_
timestamp 1704896540
transform -1 0 26772 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1370_
timestamp 1704896540
transform 1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1704896540
transform -1 0 24380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1372_
timestamp 1704896540
transform -1 0 23736 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1704896540
transform 1 0 25300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1374_
timestamp 1704896540
transform -1 0 25300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1375_
timestamp 1704896540
transform -1 0 29440 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1376_
timestamp 1704896540
transform -1 0 25024 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1377_
timestamp 1704896540
transform 1 0 25484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1378_
timestamp 1704896540
transform 1 0 24380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1379_
timestamp 1704896540
transform -1 0 25760 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1380_
timestamp 1704896540
transform 1 0 23092 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1381_
timestamp 1704896540
transform 1 0 22632 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1382_
timestamp 1704896540
transform -1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1383_
timestamp 1704896540
transform 1 0 9752 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1384_
timestamp 1704896540
transform -1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1385_
timestamp 1704896540
transform -1 0 13248 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1386_
timestamp 1704896540
transform -1 0 12512 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1387_
timestamp 1704896540
transform 1 0 14444 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1388_
timestamp 1704896540
transform -1 0 13248 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1389_
timestamp 1704896540
transform -1 0 15916 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15916 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1704896540
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1392_
timestamp 1704896540
transform 1 0 14444 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1704896540
transform 1 0 13708 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1394_
timestamp 1704896540
transform -1 0 14444 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1395_
timestamp 1704896540
transform 1 0 21988 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1396_
timestamp 1704896540
transform 1 0 22816 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 1704896540
transform -1 0 24380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1398_
timestamp 1704896540
transform 1 0 21160 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1399_
timestamp 1704896540
transform 1 0 22540 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 1704896540
transform 1 0 22540 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1401_
timestamp 1704896540
transform -1 0 24104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1402_
timestamp 1704896540
transform -1 0 15732 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1403_
timestamp 1704896540
transform 1 0 23368 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1404_
timestamp 1704896540
transform 1 0 22816 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1405_
timestamp 1704896540
transform -1 0 23276 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1406_
timestamp 1704896540
transform 1 0 26128 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1704896540
transform -1 0 20148 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1408_
timestamp 1704896540
transform -1 0 22448 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_4  _1409_
timestamp 1704896540
transform 1 0 17940 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _1410_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18768 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _1411_
timestamp 1704896540
transform 1 0 23736 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1412_
timestamp 1704896540
transform 1 0 21804 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1413_
timestamp 1704896540
transform 1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1414_
timestamp 1704896540
transform -1 0 23368 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1415_
timestamp 1704896540
transform -1 0 22448 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1416_
timestamp 1704896540
transform -1 0 27048 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1417_
timestamp 1704896540
transform 1 0 21252 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1418_
timestamp 1704896540
transform -1 0 20608 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1419_
timestamp 1704896540
transform 1 0 20608 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1420_
timestamp 1704896540
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1421_
timestamp 1704896540
transform 1 0 21528 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1422_
timestamp 1704896540
transform -1 0 22448 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1704896540
transform 1 0 20792 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1424_
timestamp 1704896540
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1425_
timestamp 1704896540
transform -1 0 21896 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1426_
timestamp 1704896540
transform -1 0 21620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _1427_
timestamp 1704896540
transform 1 0 21712 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_4  _1428_
timestamp 1704896540
transform -1 0 14628 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1429_
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1430_
timestamp 1704896540
transform 1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1431_
timestamp 1704896540
transform 1 0 25484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1704896540
transform -1 0 23276 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1433_
timestamp 1704896540
transform -1 0 19504 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1434_
timestamp 1704896540
transform 1 0 18492 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1435_
timestamp 1704896540
transform 1 0 22172 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1436_
timestamp 1704896540
transform 1 0 23276 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1437_
timestamp 1704896540
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1438_
timestamp 1704896540
transform 1 0 24932 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1439_
timestamp 1704896540
transform -1 0 24748 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1440_
timestamp 1704896540
transform 1 0 27232 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1441_
timestamp 1704896540
transform -1 0 27784 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1442_
timestamp 1704896540
transform -1 0 25300 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1443_
timestamp 1704896540
transform 1 0 24288 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1704896540
transform -1 0 20424 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1445_
timestamp 1704896540
transform 1 0 15088 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1446_
timestamp 1704896540
transform 1 0 18676 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1447_
timestamp 1704896540
transform 1 0 13800 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1448_
timestamp 1704896540
transform 1 0 16192 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1449_
timestamp 1704896540
transform -1 0 15088 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1450_
timestamp 1704896540
transform 1 0 15272 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1451_
timestamp 1704896540
transform 1 0 14628 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1452_
timestamp 1704896540
transform 1 0 14076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1453_
timestamp 1704896540
transform 1 0 16468 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1454_
timestamp 1704896540
transform -1 0 25852 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1455_
timestamp 1704896540
transform 1 0 23828 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1456_
timestamp 1704896540
transform 1 0 20148 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1457_
timestamp 1704896540
transform -1 0 22816 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _1458_
timestamp 1704896540
transform -1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _1459_
timestamp 1704896540
transform -1 0 17296 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1460_
timestamp 1704896540
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1461_
timestamp 1704896540
transform -1 0 15732 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1704896540
transform -1 0 14996 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1463_
timestamp 1704896540
transform -1 0 15916 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 1704896540
transform 1 0 19504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1465_
timestamp 1704896540
transform -1 0 18768 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1466_
timestamp 1704896540
transform 1 0 16836 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1467_
timestamp 1704896540
transform 1 0 19504 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19412 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1469_
timestamp 1704896540
transform -1 0 18584 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1470_
timestamp 1704896540
transform -1 0 19504 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1471_
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1472_
timestamp 1704896540
transform -1 0 19872 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1473_
timestamp 1704896540
transform 1 0 20792 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1474_
timestamp 1704896540
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1475_
timestamp 1704896540
transform 1 0 20424 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1476_
timestamp 1704896540
transform 1 0 19872 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1478_
timestamp 1704896540
transform 1 0 18860 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1479_
timestamp 1704896540
transform -1 0 15640 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1480_
timestamp 1704896540
transform 1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1481_
timestamp 1704896540
transform -1 0 14904 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1482_
timestamp 1704896540
transform 1 0 6164 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1704896540
transform 1 0 5888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 29900 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_1  _1485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28980 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1486_
timestamp 1704896540
transform 1 0 27692 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1704896540
transform 1 0 24564 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1488_
timestamp 1704896540
transform 1 0 23736 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1489_
timestamp 1704896540
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1490_
timestamp 1704896540
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1491_
timestamp 1704896540
transform 1 0 26404 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1492_
timestamp 1704896540
transform 1 0 25484 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1493_
timestamp 1704896540
transform 1 0 24840 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1494_
timestamp 1704896540
transform -1 0 16192 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1495_
timestamp 1704896540
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1496_
timestamp 1704896540
transform 1 0 11224 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1497_
timestamp 1704896540
transform 1 0 11592 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1498_
timestamp 1704896540
transform 1 0 12236 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1499_
timestamp 1704896540
transform 1 0 11224 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1500_
timestamp 1704896540
transform -1 0 11592 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1501_
timestamp 1704896540
transform -1 0 29348 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1502_
timestamp 1704896540
transform 1 0 29900 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1503_
timestamp 1704896540
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1504_
timestamp 1704896540
transform 1 0 30176 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1505_
timestamp 1704896540
transform 1 0 29900 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1506_
timestamp 1704896540
transform 1 0 26956 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1507_
timestamp 1704896540
transform 1 0 24748 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1508_
timestamp 1704896540
transform 1 0 24380 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 1704896540
transform -1 0 20332 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1510_
timestamp 1704896540
transform -1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1704896540
transform -1 0 17112 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1512_
timestamp 1704896540
transform -1 0 19504 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 1704896540
transform -1 0 17204 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1514_
timestamp 1704896540
transform 1 0 16652 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1515_
timestamp 1704896540
transform -1 0 16836 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1516_
timestamp 1704896540
transform -1 0 15548 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1517_
timestamp 1704896540
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 1704896540
transform -1 0 18216 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1519_
timestamp 1704896540
transform -1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1520_
timestamp 1704896540
transform 1 0 17112 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1521_
timestamp 1704896540
transform 1 0 17572 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1522_
timestamp 1704896540
transform -1 0 18860 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _1523_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18216 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _1524_
timestamp 1704896540
transform 1 0 17756 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1525_
timestamp 1704896540
transform -1 0 20976 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1526_
timestamp 1704896540
transform -1 0 20240 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1527_
timestamp 1704896540
transform 1 0 18952 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1528_
timestamp 1704896540
transform 1 0 15180 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1704896540
transform -1 0 14996 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1530_
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1531_
timestamp 1704896540
transform -1 0 14720 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1704896540
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1704896540
transform 1 0 1472 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1534_
timestamp 1704896540
transform -1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1535_
timestamp 1704896540
transform -1 0 22540 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1536_
timestamp 1704896540
transform 1 0 22080 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1537_
timestamp 1704896540
transform 1 0 21436 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1538_
timestamp 1704896540
transform -1 0 21896 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1539_
timestamp 1704896540
transform 1 0 19964 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1540_
timestamp 1704896540
transform 1 0 20884 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1704896540
transform -1 0 19320 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1542_
timestamp 1704896540
transform -1 0 18584 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1543_
timestamp 1704896540
transform 1 0 19320 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1544_
timestamp 1704896540
transform -1 0 21436 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1545_
timestamp 1704896540
transform -1 0 19412 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1546_
timestamp 1704896540
transform -1 0 19780 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1547_
timestamp 1704896540
transform 1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1548_
timestamp 1704896540
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1549_
timestamp 1704896540
transform -1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1550_
timestamp 1704896540
transform -1 0 20424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1551_
timestamp 1704896540
transform -1 0 20148 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1552_
timestamp 1704896540
transform 1 0 19320 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1553_
timestamp 1704896540
transform -1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1554_
timestamp 1704896540
transform -1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1555_
timestamp 1704896540
transform 1 0 20516 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1556_
timestamp 1704896540
transform -1 0 21896 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1557_
timestamp 1704896540
transform 1 0 20056 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1558_
timestamp 1704896540
transform 1 0 19596 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1559_
timestamp 1704896540
transform -1 0 15180 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1560_
timestamp 1704896540
transform 1 0 17388 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1561_
timestamp 1704896540
transform 1 0 20148 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1562_
timestamp 1704896540
transform -1 0 17848 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1563_
timestamp 1704896540
transform -1 0 16928 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1564_
timestamp 1704896540
transform -1 0 17296 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1565_
timestamp 1704896540
transform 1 0 14352 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1566_
timestamp 1704896540
transform -1 0 17848 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1567_
timestamp 1704896540
transform 1 0 16652 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1568_
timestamp 1704896540
transform 1 0 17756 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1569_
timestamp 1704896540
transform -1 0 18584 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1570_
timestamp 1704896540
transform -1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1571_
timestamp 1704896540
transform 1 0 19596 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1572_
timestamp 1704896540
transform 1 0 19412 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1573_
timestamp 1704896540
transform -1 0 19872 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1574_
timestamp 1704896540
transform 1 0 17848 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1575_
timestamp 1704896540
transform -1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1576_
timestamp 1704896540
transform -1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1577_
timestamp 1704896540
transform -1 0 15180 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1578_
timestamp 1704896540
transform 1 0 13800 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 1704896540
transform 1 0 3680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1704896540
transform -1 0 3772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1581_
timestamp 1704896540
transform 1 0 14996 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1582_
timestamp 1704896540
transform -1 0 14996 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1583_
timestamp 1704896540
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1704896540
transform 1 0 1196 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1704896540
transform -1 0 17480 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1704896540
transform -1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1587_
timestamp 1704896540
transform -1 0 17296 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1704896540
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1589_
timestamp 1704896540
transform -1 0 27232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1590_
timestamp 1704896540
transform -1 0 27508 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1704896540
transform -1 0 26312 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1592_
timestamp 1704896540
transform 1 0 28704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 1704896540
transform -1 0 26128 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1704896540
transform 1 0 28980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 1704896540
transform -1 0 26312 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1596_
timestamp 1704896540
transform 1 0 27876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1597_
timestamp 1704896540
transform -1 0 19964 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1704896540
transform 1 0 19964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1599_
timestamp 1704896540
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1704896540
transform -1 0 22908 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1601_
timestamp 1704896540
transform -1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1602_
timestamp 1704896540
transform 1 0 12880 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1603_
timestamp 1704896540
transform 1 0 15640 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1604_
timestamp 1704896540
transform 1 0 13616 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o41ai_1  _1605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14168 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1606_
timestamp 1704896540
transform -1 0 16560 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1607_
timestamp 1704896540
transform 1 0 11040 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1608_
timestamp 1704896540
transform 1 0 12144 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1609_
timestamp 1704896540
transform -1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1611_
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1704896540
transform -1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1613_
timestamp 1704896540
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1704896540
transform -1 0 10764 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1615_
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1704896540
transform -1 0 11316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1617_
timestamp 1704896540
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1704896540
transform -1 0 8648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1619_
timestamp 1704896540
transform 1 0 10856 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1620_
timestamp 1704896540
transform -1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1704896540
transform -1 0 10856 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1622_
timestamp 1704896540
transform -1 0 10764 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1623_
timestamp 1704896540
transform -1 0 11500 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1704896540
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1625_
timestamp 1704896540
transform -1 0 10028 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1626_
timestamp 1704896540
transform -1 0 8832 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1627_
timestamp 1704896540
transform 1 0 8832 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1628_
timestamp 1704896540
transform -1 0 8280 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1629_
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1630_
timestamp 1704896540
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1631_
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1704896540
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1633_
timestamp 1704896540
transform 1 0 8740 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1704896540
transform 1 0 8464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1635_
timestamp 1704896540
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1636_
timestamp 1704896540
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 1704896540
transform 1 0 1840 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1638_
timestamp 1704896540
transform 1 0 1472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1639_
timestamp 1704896540
transform 1 0 1656 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1640_
timestamp 1704896540
transform -1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1641_
timestamp 1704896540
transform 1 0 2484 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1642_
timestamp 1704896540
transform -1 0 1196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1643_
timestamp 1704896540
transform -1 0 10212 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1644_
timestamp 1704896540
transform -1 0 9752 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1645_
timestamp 1704896540
transform -1 0 8280 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1646_
timestamp 1704896540
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1704896540
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1704896540
transform -1 0 4876 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1649_
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1650_
timestamp 1704896540
transform 1 0 2760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1651_
timestamp 1704896540
transform -1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1652_
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1653_
timestamp 1704896540
transform 1 0 7084 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1704896540
transform -1 0 6256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1655_
timestamp 1704896540
transform 1 0 1656 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1656_
timestamp 1704896540
transform 1 0 1196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1657_
timestamp 1704896540
transform 1 0 1656 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1658_
timestamp 1704896540
transform 1 0 1196 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1704896540
transform 1 0 1288 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1704896540
transform 1 0 1012 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1661_
timestamp 1704896540
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1662_
timestamp 1704896540
transform -1 0 9660 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1663_
timestamp 1704896540
transform 1 0 11592 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1664_
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1665_
timestamp 1704896540
transform -1 0 4968 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1704896540
transform 1 0 4876 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1704896540
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1669_
timestamp 1704896540
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1704896540
transform 1 0 6624 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1671_
timestamp 1704896540
transform -1 0 5060 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1704896540
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1675_
timestamp 1704896540
transform 1 0 2668 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1677_
timestamp 1704896540
transform -1 0 1288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1704896540
transform 1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _1680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9292 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1704896540
transform 1 0 7360 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1704896540
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1704896540
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1704896540
transform 1 0 2300 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1704896540
transform -1 0 1196 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1704896540
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1704896540
transform -1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1704896540
transform 1 0 6256 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1690_
timestamp 1704896540
transform -1 0 6072 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1704896540
transform -1 0 3128 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1704896540
transform 1 0 3220 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1704896540
transform 1 0 3496 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1704896540
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1695_
timestamp 1704896540
transform 1 0 3036 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1704896540
transform -1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1697_
timestamp 1704896540
transform 1 0 8924 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1698_
timestamp 1704896540
transform 1 0 9292 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1699_
timestamp 1704896540
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1700_
timestamp 1704896540
transform -1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 1704896540
transform 1 0 12328 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1702_
timestamp 1704896540
transform -1 0 12604 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1704896540
transform 1 0 12604 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1704896540
transform -1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1704896540
transform 1 0 5612 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1704896540
transform -1 0 5612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1708_
timestamp 1704896540
transform -1 0 11224 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1704896540
transform 1 0 2668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1704896540
transform -1 0 2116 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1704896540
transform 1 0 2668 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1704896540
transform 1 0 3220 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1704896540
transform -1 0 3128 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1715_
timestamp 1704896540
transform 1 0 9476 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1716_
timestamp 1704896540
transform 1 0 10304 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1704896540
transform 1 0 7176 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1704896540
transform -1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 1704896540
transform -1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1704896540
transform 1 0 5152 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 1704896540
transform 1 0 3312 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1704896540
transform -1 0 3404 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1704896540
transform 1 0 5888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1725_
timestamp 1704896540
transform -1 0 7912 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1704896540
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1704896540
transform 1 0 1472 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1704896540
transform 1 0 1196 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 1704896540
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1730_
timestamp 1704896540
transform 1 0 1196 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 1704896540
transform 1 0 1656 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1732_
timestamp 1704896540
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1733_
timestamp 1704896540
transform 1 0 15456 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1734_
timestamp 1704896540
transform -1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1735_
timestamp 1704896540
transform 1 0 17112 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1736_
timestamp 1704896540
transform 1 0 17572 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1737_
timestamp 1704896540
transform -1 0 18492 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1738_
timestamp 1704896540
transform 1 0 16284 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1739_
timestamp 1704896540
transform 1 0 17940 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1740_
timestamp 1704896540
transform 1 0 18676 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1741_
timestamp 1704896540
transform 1 0 17940 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 1704896540
transform -1 0 24196 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1743_
timestamp 1704896540
transform 1 0 25668 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1704896540
transform 1 0 26404 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1745_
timestamp 1704896540
transform -1 0 26312 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1704896540
transform 1 0 27416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1704896540
transform -1 0 27876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1704896540
transform -1 0 25668 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1704896540
transform -1 0 26220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1704896540
transform -1 0 21160 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1704896540
transform 1 0 24196 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1704896540
transform 1 0 25116 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1704896540
transform 1 0 24840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1704896540
transform -1 0 23736 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1704896540
transform 1 0 25944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1704896540
transform 1 0 21252 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1757_
timestamp 1704896540
transform -1 0 20608 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1758_
timestamp 1704896540
transform -1 0 11592 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1759_
timestamp 1704896540
transform -1 0 9568 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1760_
timestamp 1704896540
transform -1 0 12512 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1761_
timestamp 1704896540
transform -1 0 8464 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1762_
timestamp 1704896540
transform -1 0 11408 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1763_
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1764_
timestamp 1704896540
transform 1 0 16836 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1765_
timestamp 1704896540
transform -1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 1704896540
transform 1 0 3128 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1704896540
transform 1 0 17756 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_2  _1768_
timestamp 1704896540
transform 1 0 17664 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1769_
timestamp 1704896540
transform -1 0 18216 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 1704896540
transform 1 0 2024 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1771_
timestamp 1704896540
transform 1 0 1196 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1772_
timestamp 1704896540
transform 1 0 3220 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1773_
timestamp 1704896540
transform 1 0 5704 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1774_
timestamp 1704896540
transform 1 0 5796 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1704896540
transform 1 0 3956 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1704896540
transform 1 0 3680 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1777_
timestamp 1704896540
transform -1 0 3128 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1778_
timestamp 1704896540
transform 1 0 4968 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1779_
timestamp 1704896540
transform 1 0 4232 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1780_
timestamp 1704896540
transform -1 0 4232 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1781_
timestamp 1704896540
transform 1 0 4324 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1704896540
transform -1 0 3128 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1704896540
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1784__1
timestamp 1704896540
transform 1 0 12420 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1785_
timestamp 1704896540
transform -1 0 17940 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1786_
timestamp 1704896540
transform 1 0 18216 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1787_
timestamp 1704896540
transform -1 0 18400 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 1704896540
transform -1 0 16560 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1789_
timestamp 1704896540
transform 1 0 16928 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1790_
timestamp 1704896540
transform -1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1791_
timestamp 1704896540
transform -1 0 15824 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1704896540
transform -1 0 15456 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1793_
timestamp 1704896540
transform -1 0 18584 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1794_
timestamp 1704896540
transform 1 0 18216 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1795_
timestamp 1704896540
transform -1 0 18216 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1796_
timestamp 1704896540
transform -1 0 11776 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1797_
timestamp 1704896540
transform 1 0 10488 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1798_
timestamp 1704896540
transform 1 0 10212 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1799_
timestamp 1704896540
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1800_
timestamp 1704896540
transform -1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1801_
timestamp 1704896540
transform -1 0 10212 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1802_
timestamp 1704896540
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1803_
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1804_
timestamp 1704896540
transform -1 0 10120 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1805_
timestamp 1704896540
transform 1 0 10120 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1806_
timestamp 1704896540
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1807_
timestamp 1704896540
transform -1 0 10488 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1808_
timestamp 1704896540
transform -1 0 9568 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1809_
timestamp 1704896540
transform 1 0 9292 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1810_
timestamp 1704896540
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1811_
timestamp 1704896540
transform 1 0 10488 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1812_
timestamp 1704896540
transform -1 0 8648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1813_
timestamp 1704896540
transform 1 0 9568 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1814_
timestamp 1704896540
transform 1 0 11132 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1815_
timestamp 1704896540
transform 1 0 9292 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1816_
timestamp 1704896540
transform 1 0 8280 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1817_
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1818_
timestamp 1704896540
transform 1 0 9752 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1819_
timestamp 1704896540
transform 1 0 11132 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1820_
timestamp 1704896540
transform 1 0 8648 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1821_
timestamp 1704896540
transform 1 0 9200 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1822_
timestamp 1704896540
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1823_
timestamp 1704896540
transform 1 0 9476 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1824_
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1825_
timestamp 1704896540
transform 1 0 7820 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1826_
timestamp 1704896540
transform 1 0 12236 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1827_
timestamp 1704896540
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1828_
timestamp 1704896540
transform -1 0 9936 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1829_
timestamp 1704896540
transform -1 0 10948 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1830_
timestamp 1704896540
transform -1 0 6716 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1831_
timestamp 1704896540
transform -1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1832_
timestamp 1704896540
transform -1 0 10120 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1833_
timestamp 1704896540
transform -1 0 11408 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1834_
timestamp 1704896540
transform -1 0 12144 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1835_
timestamp 1704896540
transform 1 0 9200 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1836_
timestamp 1704896540
transform -1 0 10488 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1837_
timestamp 1704896540
transform 1 0 10396 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1838_
timestamp 1704896540
transform -1 0 8280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1839_
timestamp 1704896540
transform -1 0 10672 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1840_
timestamp 1704896540
transform -1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1841_
timestamp 1704896540
transform 1 0 15732 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1842_
timestamp 1704896540
transform -1 0 16744 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1843_
timestamp 1704896540
transform -1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 1704896540
transform -1 0 6900 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1845_
timestamp 1704896540
transform -1 0 6900 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 1704896540
transform 1 0 6256 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1847_
timestamp 1704896540
transform -1 0 5704 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1848_
timestamp 1704896540
transform -1 0 8280 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1849_
timestamp 1704896540
transform 1 0 8924 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1850_
timestamp 1704896540
transform 1 0 4600 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1851_
timestamp 1704896540
transform -1 0 3588 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1852_
timestamp 1704896540
transform 1 0 3588 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1853_
timestamp 1704896540
transform -1 0 3312 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 1704896540
transform 1 0 1196 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1855_
timestamp 1704896540
transform -1 0 1196 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1856_
timestamp 1704896540
transform 1 0 1472 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1857_
timestamp 1704896540
transform -1 0 1196 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1858_
timestamp 1704896540
transform 1 0 5796 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1859_
timestamp 1704896540
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12328 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1861_
timestamp 1704896540
transform -1 0 10120 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1862_
timestamp 1704896540
transform 1 0 10580 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1863_
timestamp 1704896540
transform 1 0 7452 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1864_
timestamp 1704896540
transform 1 0 5704 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1865_
timestamp 1704896540
transform 1 0 1012 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1866_
timestamp 1704896540
transform 1 0 3864 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1868_
timestamp 1704896540
transform -1 0 18400 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1869_
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 28336 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1871_
timestamp 1704896540
transform 1 0 26496 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1872_
timestamp 1704896540
transform 1 0 26864 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26772 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1874_
timestamp 1704896540
transform 1 0 19412 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1875_
timestamp 1704896540
transform 1 0 22816 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1876_
timestamp 1704896540
transform 1 0 24932 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1877_
timestamp 1704896540
transform -1 0 29440 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1878_
timestamp 1704896540
transform 1 0 26864 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1879_
timestamp 1704896540
transform 1 0 15732 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1880_
timestamp 1704896540
transform 1 0 13800 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1881_
timestamp 1704896540
transform -1 0 13340 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1882_
timestamp 1704896540
transform 1 0 12512 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1883_
timestamp 1704896540
transform 1 0 11592 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1884_
timestamp 1704896540
transform 1 0 11316 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1885_
timestamp 1704896540
transform 1 0 9844 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1886_
timestamp 1704896540
transform 1 0 11224 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1887_
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1888_
timestamp 1704896540
transform -1 0 13432 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1889_
timestamp 1704896540
transform 1 0 8556 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1890_
timestamp 1704896540
transform 1 0 4416 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1891_
timestamp 1704896540
transform 1 0 2024 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1892_
timestamp 1704896540
transform 1 0 8096 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1893_
timestamp 1704896540
transform 1 0 6256 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1894_
timestamp 1704896540
transform 1 0 1104 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1895_
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1896_
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1897_
timestamp 1704896540
transform -1 0 8280 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1898_
timestamp 1704896540
transform 1 0 4508 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1899_
timestamp 1704896540
transform 1 0 2116 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1900_
timestamp 1704896540
transform -1 0 10212 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1901_
timestamp 1704896540
transform 1 0 6348 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1902_
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1903_
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1904_
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1905_
timestamp 1704896540
transform 1 0 7728 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1906_
timestamp 1704896540
transform 1 0 3864 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1907_
timestamp 1704896540
transform 1 0 2484 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1908_
timestamp 1704896540
transform 1 0 5888 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1909_
timestamp 1704896540
transform 1 0 4784 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1910_
timestamp 1704896540
transform 1 0 2116 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1911_
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1912_
timestamp 1704896540
transform 1 0 2208 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1913_
timestamp 1704896540
transform 1 0 5520 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1914_
timestamp 1704896540
transform 1 0 4508 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1915_
timestamp 1704896540
transform 1 0 1196 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1916_
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1917_
timestamp 1704896540
transform 1 0 6164 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1918_
timestamp 1704896540
transform 1 0 2668 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1919_
timestamp 1704896540
transform 1 0 3036 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1920_
timestamp 1704896540
transform -1 0 5152 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1921_
timestamp 1704896540
transform 1 0 11040 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1922_
timestamp 1704896540
transform 1 0 13616 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1923_
timestamp 1704896540
transform 1 0 12788 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1924_
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1925_
timestamp 1704896540
transform 1 0 13156 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1926_
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1927_
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1928_
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1929_
timestamp 1704896540
transform 1 0 6532 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1930_
timestamp 1704896540
transform -1 0 5244 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1931_
timestamp 1704896540
transform 1 0 3404 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1932_
timestamp 1704896540
transform 1 0 5520 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1933_
timestamp 1704896540
transform -1 0 8464 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1934_
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1935_
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1936_
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1937_
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1938_
timestamp 1704896540
transform -1 0 23736 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1939_
timestamp 1704896540
transform -1 0 28336 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1940_
timestamp 1704896540
transform 1 0 28336 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1941_
timestamp 1704896540
transform -1 0 26404 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1942_
timestamp 1704896540
transform -1 0 23368 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1943_
timestamp 1704896540
transform 1 0 24380 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1944_
timestamp 1704896540
transform -1 0 25208 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1945_
timestamp 1704896540
transform 1 0 20700 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1946_
timestamp 1704896540
transform 1 0 828 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1947_
timestamp 1704896540
transform 1 0 3588 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1948_
timestamp 1704896540
transform 1 0 1012 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1949_
timestamp 1704896540
transform -1 0 13248 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1950_
timestamp 1704896540
transform -1 0 25484 0 -1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1951_
timestamp 1704896540
transform -1 0 20792 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1952_
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1953_
timestamp 1704896540
transform 1 0 11960 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1954_
timestamp 1704896540
transform 1 0 11316 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1955_
timestamp 1704896540
transform 1 0 11684 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1956_
timestamp 1704896540
transform 1 0 11224 0 1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1957_
timestamp 1704896540
transform 1 0 10304 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1958_
timestamp 1704896540
transform 1 0 5796 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1959_
timestamp 1704896540
transform 1 0 9568 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1960_
timestamp 1704896540
transform 1 0 8556 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1961_
timestamp 1704896540
transform 1 0 8004 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1962_
timestamp 1704896540
transform -1 0 7636 0 1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1963_
timestamp 1704896540
transform 1 0 5888 0 -1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1964_
timestamp 1704896540
transform -1 0 9108 0 -1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1965_
timestamp 1704896540
transform 1 0 3588 0 1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1966_
timestamp 1704896540
transform 1 0 3220 0 1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1967_
timestamp 1704896540
transform 1 0 920 0 -1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1968_
timestamp 1704896540
transform 1 0 828 0 -1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_4  _1969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3128 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform -1 0 21620 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1704896540
transform -1 0 19504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1704896540
transform -1 0 20976 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1704896540
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1704896540
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17020 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1704896540
transform -1 0 8280 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1704896540
transform -1 0 8280 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1704896540
transform -1 0 8188 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1704896540
transform -1 0 9108 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1704896540
transform -1 0 15732 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1704896540
transform 1 0 21528 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1704896540
transform 1 0 21896 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1704896540
transform -1 0 6348 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1704896540
transform -1 0 7176 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1704896540
transform -1 0 15640 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1704896540
transform 1 0 16560 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1704896540
transform -1 0 16008 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1704896540
transform -1 0 5428 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1704896540
transform -1 0 9568 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1704896540
transform -1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1704896540
transform -1 0 10304 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1704896540
transform -1 0 13432 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1704896540
transform -1 0 29532 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1704896540
transform -1 0 29900 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1704896540
transform 1 0 29992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1704896540
transform -1 0 29992 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1704896540
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1704896540
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1704896540
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1704896540
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1704896540
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1704896540
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1704896540
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1704896540
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1704896540
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1704896540
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1704896540
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_193
timestamp 1704896540
transform 1 0 18308 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_205
timestamp 1704896540
transform 1 0 19412 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_209
timestamp 1704896540
transform 1 0 19780 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 1704896540
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1704896540
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1704896540
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1704896540
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1704896540
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1704896540
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1704896540
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1704896540
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1704896540
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1704896540
transform 1 0 30820 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_149
timestamp 1704896540
transform 1 0 14260 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1704896540
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_184
timestamp 1704896540
transform 1 0 17480 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_190
timestamp 1704896540
transform 1 0 18032 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1704896540
transform 1 0 19780 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_228
timestamp 1704896540
transform 1 0 21528 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_238
timestamp 1704896540
transform 1 0 22448 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1704896540
transform 1 0 23552 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_253
timestamp 1704896540
transform 1 0 23828 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_272
timestamp 1704896540
transform 1 0 25576 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_280
timestamp 1704896540
transform 1 0 26312 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_285
timestamp 1704896540
transform 1 0 26772 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_297
timestamp 1704896540
transform 1 0 27876 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_305
timestamp 1704896540
transform 1 0 28612 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1704896540
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1704896540
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1704896540
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_77
timestamp 1704896540
transform 1 0 7636 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_86
timestamp 1704896540
transform 1 0 8464 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1704896540
transform 1 0 10304 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_153
timestamp 1704896540
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_206
timestamp 1704896540
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_210
timestamp 1704896540
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_229
timestamp 1704896540
transform 1 0 21620 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_251
timestamp 1704896540
transform 1 0 23644 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_274
timestamp 1704896540
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_294
timestamp 1704896540
transform 1 0 27600 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_306
timestamp 1704896540
transform 1 0 28704 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_318
timestamp 1704896540
transform 1 0 29808 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_330
timestamp 1704896540
transform 1 0 30912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_334
timestamp 1704896540
transform 1 0 31280 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_11
timestamp 1704896540
transform 1 0 1564 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_23
timestamp 1704896540
transform 1 0 2668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_43
timestamp 1704896540
transform 1 0 4508 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_55
timestamp 1704896540
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_79
timestamp 1704896540
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_98
timestamp 1704896540
transform 1 0 9568 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_130
timestamp 1704896540
transform 1 0 12512 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1704896540
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_168
timestamp 1704896540
transform 1 0 16008 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_174
timestamp 1704896540
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_192
timestamp 1704896540
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_202
timestamp 1704896540
transform 1 0 19136 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_214
timestamp 1704896540
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_225
timestamp 1704896540
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_232
timestamp 1704896540
transform 1 0 21896 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_238
timestamp 1704896540
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_274
timestamp 1704896540
transform 1 0 25760 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_280
timestamp 1704896540
transform 1 0 26312 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_292
timestamp 1704896540
transform 1 0 27416 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_304
timestamp 1704896540
transform 1 0 28520 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1704896540
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1704896540
transform 1 0 30084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 1704896540
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1704896540
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_13
timestamp 1704896540
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1704896540
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_143
timestamp 1704896540
transform 1 0 13708 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp 1704896540
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_177
timestamp 1704896540
transform 1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_238
timestamp 1704896540
transform 1 0 22448 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_244
timestamp 1704896540
transform 1 0 23000 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_252
timestamp 1704896540
transform 1 0 23736 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_266
timestamp 1704896540
transform 1 0 25024 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_274
timestamp 1704896540
transform 1 0 25760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26404 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_299
timestamp 1704896540
transform 1 0 28060 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_311
timestamp 1704896540
transform 1 0 29164 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_323
timestamp 1704896540
transform 1 0 30268 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1704896540
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_38
timestamp 1704896540
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_80
timestamp 1704896540
transform 1 0 7912 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_165
timestamp 1704896540
transform 1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_169
timestamp 1704896540
transform 1 0 16100 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_181
timestamp 1704896540
transform 1 0 17204 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp 1704896540
transform 1 0 18124 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_197
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_207
timestamp 1704896540
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_217
timestamp 1704896540
transform 1 0 20516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_234
timestamp 1704896540
transform 1 0 22080 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_260
timestamp 1704896540
transform 1 0 24472 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1704896540
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1704896540
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1704896540
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1704896540
transform 1 0 30084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1704896540
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_10
timestamp 1704896540
transform 1 0 1472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_41
timestamp 1704896540
transform 1 0 4324 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_83
timestamp 1704896540
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_148
timestamp 1704896540
transform 1 0 14168 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_172
timestamp 1704896540
transform 1 0 16376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_186
timestamp 1704896540
transform 1 0 17664 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_196
timestamp 1704896540
transform 1 0 18584 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_202
timestamp 1704896540
transform 1 0 19136 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1704896540
transform 1 0 20976 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_241
timestamp 1704896540
transform 1 0 22724 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_258
timestamp 1704896540
transform 1 0 24288 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_268
timestamp 1704896540
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1704896540
transform 1 0 26036 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_298
timestamp 1704896540
transform 1 0 27968 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_310
timestamp 1704896540
transform 1 0 29072 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_322
timestamp 1704896540
transform 1 0 30176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_334
timestamp 1704896540
transform 1 0 31280 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_23
timestamp 1704896540
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_38
timestamp 1704896540
transform 1 0 4048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_62
timestamp 1704896540
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_107
timestamp 1704896540
transform 1 0 10396 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_157
timestamp 1704896540
transform 1 0 14996 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_161
timestamp 1704896540
transform 1 0 15364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_172
timestamp 1704896540
transform 1 0 16376 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_210
timestamp 1704896540
transform 1 0 19872 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_216
timestamp 1704896540
transform 1 0 20424 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_257
timestamp 1704896540
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26036 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_304
timestamp 1704896540
transform 1 0 28520 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_318
timestamp 1704896540
transform 1 0 29808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_330
timestamp 1704896540
transform 1 0 30912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_334
timestamp 1704896540
transform 1 0 31280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_99
timestamp 1704896540
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_141
timestamp 1704896540
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_182
timestamp 1704896540
transform 1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_195
timestamp 1704896540
transform 1 0 18492 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_203
timestamp 1704896540
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1704896540
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_265
timestamp 1704896540
transform 1 0 24932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_287
timestamp 1704896540
transform 1 0 26956 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1704896540
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1704896540
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_38
timestamp 1704896540
transform 1 0 4048 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1704896540
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_148
timestamp 1704896540
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_157
timestamp 1704896540
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_168
timestamp 1704896540
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_177
timestamp 1704896540
transform 1 0 16836 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1704896540
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_205
timestamp 1704896540
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_216
timestamp 1704896540
transform 1 0 20424 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1704896540
transform 1 0 23552 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_282
timestamp 1704896540
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_315
timestamp 1704896540
transform 1 0 29532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_327
timestamp 1704896540
transform 1 0 30636 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_98
timestamp 1704896540
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_107
timestamp 1704896540
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_116
timestamp 1704896540
transform 1 0 11224 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_178
timestamp 1704896540
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_182
timestamp 1704896540
transform 1 0 17296 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_188
timestamp 1704896540
transform 1 0 17848 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_195
timestamp 1704896540
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_202
timestamp 1704896540
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_206
timestamp 1704896540
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_218
timestamp 1704896540
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1704896540
transform 1 0 20976 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_247
timestamp 1704896540
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_270
timestamp 1704896540
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_285
timestamp 1704896540
transform 1 0 26772 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_312
timestamp 1704896540
transform 1 0 29256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_324
timestamp 1704896540
transform 1 0 30360 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_332
timestamp 1704896540
transform 1 0 31096 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1704896540
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_49
timestamp 1704896540
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_182
timestamp 1704896540
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_188
timestamp 1704896540
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_217
timestamp 1704896540
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_234
timestamp 1704896540
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_247
timestamp 1704896540
transform 1 0 23276 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_253
timestamp 1704896540
transform 1 0 23828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_278
timestamp 1704896540
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_284
timestamp 1704896540
transform 1 0 26680 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1704896540
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1704896540
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1704896540
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_43
timestamp 1704896540
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_72
timestamp 1704896540
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_82
timestamp 1704896540
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_98
timestamp 1704896540
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1704896540
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_201
timestamp 1704896540
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_205
timestamp 1704896540
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1704896540
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1704896540
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1704896540
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_308
timestamp 1704896540
transform 1 0 28888 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_320
timestamp 1704896540
transform 1 0 29992 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_332
timestamp 1704896540
transform 1 0 31096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1704896540
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_45
timestamp 1704896540
transform 1 0 4692 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1704896540
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_103
timestamp 1704896540
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_174
timestamp 1704896540
transform 1 0 16560 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_184
timestamp 1704896540
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_200
timestamp 1704896540
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_204
timestamp 1704896540
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_215
timestamp 1704896540
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_279
timestamp 1704896540
transform 1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_283
timestamp 1704896540
transform 1 0 26588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_300
timestamp 1704896540
transform 1 0 28152 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1704896540
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1704896540
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 1704896540
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1704896540
transform 1 0 1196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_66
timestamp 1704896540
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_83
timestamp 1704896540
transform 1 0 8188 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1704896540
transform 1 0 11500 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_126
timestamp 1704896540
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_157
timestamp 1704896540
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_200
timestamp 1704896540
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_214
timestamp 1704896540
transform 1 0 20240 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_234
timestamp 1704896540
transform 1 0 22080 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_263
timestamp 1704896540
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_276
timestamp 1704896540
transform 1 0 25944 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_323
timestamp 1704896540
transform 1 0 30268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1704896540
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_38
timestamp 1704896540
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_42
timestamp 1704896540
transform 1 0 4416 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_51
timestamp 1704896540
transform 1 0 5244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_66
timestamp 1704896540
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1704896540
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_203
timestamp 1704896540
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_231
timestamp 1704896540
transform 1 0 21804 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_279
timestamp 1704896540
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_290
timestamp 1704896540
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1704896540
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1704896540
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1704896540
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1704896540
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_333
timestamp 1704896540
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1704896540
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_104
timestamp 1704896540
transform 1 0 10120 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_123
timestamp 1704896540
transform 1 0 11868 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_178
timestamp 1704896540
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_195
timestamp 1704896540
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_263
timestamp 1704896540
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1704896540
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_314
timestamp 1704896540
transform 1 0 29440 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_326
timestamp 1704896540
transform 1 0 30544 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_334
timestamp 1704896540
transform 1 0 31280 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_38
timestamp 1704896540
transform 1 0 4048 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_50
timestamp 1704896540
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1704896540
transform 1 0 9108 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1704896540
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_161
timestamp 1704896540
transform 1 0 15364 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_184
timestamp 1704896540
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 1704896540
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_220
timestamp 1704896540
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_259
timestamp 1704896540
transform 1 0 24380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_302
timestamp 1704896540
transform 1 0 28336 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_319
timestamp 1704896540
transform 1 0 29900 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_331
timestamp 1704896540
transform 1 0 31004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_10
timestamp 1704896540
transform 1 0 1472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_38
timestamp 1704896540
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1704896540
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_85
timestamp 1704896540
transform 1 0 8372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_120
timestamp 1704896540
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_144
timestamp 1704896540
transform 1 0 13800 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_183
timestamp 1704896540
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_199
timestamp 1704896540
transform 1 0 18860 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_213
timestamp 1704896540
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_271
timestamp 1704896540
transform 1 0 25484 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_304
timestamp 1704896540
transform 1 0 28520 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_324
timestamp 1704896540
transform 1 0 30360 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_332
timestamp 1704896540
transform 1 0 31096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_23
timestamp 1704896540
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_50
timestamp 1704896540
transform 1 0 5152 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_76
timestamp 1704896540
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_128
timestamp 1704896540
transform 1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_178
timestamp 1704896540
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_190
timestamp 1704896540
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_225
timestamp 1704896540
transform 1 0 21252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_248
timestamp 1704896540
transform 1 0 23368 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1704896540
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1704896540
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1704896540
transform 1 0 30084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_333
timestamp 1704896540
transform 1 0 31188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1704896540
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_13
timestamp 1704896540
transform 1 0 1748 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_25
timestamp 1704896540
transform 1 0 2852 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_33
timestamp 1704896540
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_70
timestamp 1704896540
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_74
timestamp 1704896540
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_124
timestamp 1704896540
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_151
timestamp 1704896540
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_162
timestamp 1704896540
transform 1 0 15456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_179
timestamp 1704896540
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_202
timestamp 1704896540
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_218
timestamp 1704896540
transform 1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp 1704896540
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 1704896540
transform 1 0 25852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1704896540
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_281
timestamp 1704896540
transform 1 0 26404 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_295
timestamp 1704896540
transform 1 0 27692 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_307
timestamp 1704896540
transform 1 0 28796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_319
timestamp 1704896540
transform 1 0 29900 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_331
timestamp 1704896540
transform 1 0 31004 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1704896540
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_51
timestamp 1704896540
transform 1 0 5244 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_63
timestamp 1704896540
transform 1 0 6348 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1704896540
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_94
timestamp 1704896540
transform 1 0 9200 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1704896540
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_141
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_231
timestamp 1704896540
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_237
timestamp 1704896540
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1704896540
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_275
timestamp 1704896540
transform 1 0 25852 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_279
timestamp 1704896540
transform 1 0 26220 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_287
timestamp 1704896540
transform 1 0 26956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_294
timestamp 1704896540
transform 1 0 27600 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_299
timestamp 1704896540
transform 1 0 28060 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1704896540
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_309
timestamp 1704896540
transform 1 0 28980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_317
timestamp 1704896540
transform 1 0 29716 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_324
timestamp 1704896540
transform 1 0 30360 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_332
timestamp 1704896540
transform 1 0 31096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_10
timestamp 1704896540
transform 1 0 1472 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_23
timestamp 1704896540
transform 1 0 2668 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_144
timestamp 1704896540
transform 1 0 13800 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_177
timestamp 1704896540
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1704896540
transform 1 0 20792 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_258
timestamp 1704896540
transform 1 0 24288 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_267
timestamp 1704896540
transform 1 0 25116 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_273
timestamp 1704896540
transform 1 0 25668 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_289
timestamp 1704896540
transform 1 0 27140 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_301
timestamp 1704896540
transform 1 0 28244 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_332
timestamp 1704896540
transform 1 0 31096 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_24
timestamp 1704896540
transform 1 0 2760 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5428 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_114
timestamp 1704896540
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_156
timestamp 1704896540
transform 1 0 14904 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1704896540
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_211
timestamp 1704896540
transform 1 0 19964 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_223
timestamp 1704896540
transform 1 0 21068 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_231
timestamp 1704896540
transform 1 0 21804 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1704896540
transform 1 0 23368 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_260
timestamp 1704896540
transform 1 0 24472 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_268
timestamp 1704896540
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_275
timestamp 1704896540
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_287
timestamp 1704896540
transform 1 0 26956 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_291
timestamp 1704896540
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1704896540
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1704896540
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1704896540
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_321
timestamp 1704896540
transform 1 0 30084 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_328
timestamp 1704896540
transform 1 0 30728 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_334
timestamp 1704896540
transform 1 0 31280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_124
timestamp 1704896540
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_172
timestamp 1704896540
transform 1 0 16376 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_187
timestamp 1704896540
transform 1 0 17756 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_199
timestamp 1704896540
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_210
timestamp 1704896540
transform 1 0 19872 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_216
timestamp 1704896540
transform 1 0 20424 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1704896540
transform 1 0 20976 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1704896540
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_235
timestamp 1704896540
transform 1 0 22172 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_247
timestamp 1704896540
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_251
timestamp 1704896540
transform 1 0 23644 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_259
timestamp 1704896540
transform 1 0 24380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_271
timestamp 1704896540
transform 1 0 25484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_281
timestamp 1704896540
transform 1 0 26404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_289
timestamp 1704896540
transform 1 0 27140 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_299
timestamp 1704896540
transform 1 0 28060 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_308
timestamp 1704896540
transform 1 0 28888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_316
timestamp 1704896540
transform 1 0 29624 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_333
timestamp 1704896540
transform 1 0 31188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_24
timestamp 1704896540
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_33
timestamp 1704896540
transform 1 0 3588 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_126
timestamp 1704896540
transform 1 0 12144 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1704896540
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1704896540
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1704896540
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_203
timestamp 1704896540
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_217
timestamp 1704896540
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_221
timestamp 1704896540
transform 1 0 20884 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_226
timestamp 1704896540
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_234
timestamp 1704896540
transform 1 0 22080 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1704896540
transform 1 0 23552 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 1704896540
transform 1 0 23828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_264
timestamp 1704896540
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_273
timestamp 1704896540
transform 1 0 25668 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_288
timestamp 1704896540
transform 1 0 27048 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_296
timestamp 1704896540
transform 1 0 27784 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_304
timestamp 1704896540
transform 1 0 28520 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1704896540
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_321
timestamp 1704896540
transform 1 0 30084 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_331
timestamp 1704896540
transform 1 0 31004 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1704896540
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 1704896540
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_71
timestamp 1704896540
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_102
timestamp 1704896540
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_144
timestamp 1704896540
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_152
timestamp 1704896540
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp 1704896540
transform 1 0 15640 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_182
timestamp 1704896540
transform 1 0 17296 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_190
timestamp 1704896540
transform 1 0 18032 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_208
timestamp 1704896540
transform 1 0 19688 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_216
timestamp 1704896540
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1704896540
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1704896540
transform 1 0 21252 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_233
timestamp 1704896540
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_244
timestamp 1704896540
transform 1 0 23000 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_252
timestamp 1704896540
transform 1 0 23736 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_261
timestamp 1704896540
transform 1 0 24564 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_305
timestamp 1704896540
transform 1 0 28612 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_317
timestamp 1704896540
transform 1 0 29716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_326
timestamp 1704896540
transform 1 0 30544 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_334
timestamp 1704896540
transform 1 0 31280 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3220 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_77
timestamp 1704896540
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_130
timestamp 1704896540
transform 1 0 12512 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_149
timestamp 1704896540
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_158
timestamp 1704896540
transform 1 0 15088 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_170
timestamp 1704896540
transform 1 0 16192 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_178
timestamp 1704896540
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1704896540
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_213
timestamp 1704896540
transform 1 0 20148 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_221
timestamp 1704896540
transform 1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_230
timestamp 1704896540
transform 1 0 21712 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_238
timestamp 1704896540
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_244
timestamp 1704896540
transform 1 0 23000 0 1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_259
timestamp 1704896540
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_271
timestamp 1704896540
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_283
timestamp 1704896540
transform 1 0 26588 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_296
timestamp 1704896540
transform 1 0 27784 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1704896540
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_321
timestamp 1704896540
transform 1 0 30084 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_328
timestamp 1704896540
transform 1 0 30728 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_334
timestamp 1704896540
transform 1 0 31280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_23
timestamp 1704896540
transform 1 0 2668 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_94
timestamp 1704896540
transform 1 0 9200 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_131
timestamp 1704896540
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_139
timestamp 1704896540
transform 1 0 13340 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_157
timestamp 1704896540
transform 1 0 14996 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1704896540
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_179
timestamp 1704896540
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_184
timestamp 1704896540
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_196
timestamp 1704896540
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_216
timestamp 1704896540
transform 1 0 20424 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_225
timestamp 1704896540
transform 1 0 21252 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_240
timestamp 1704896540
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_250
timestamp 1704896540
transform 1 0 23552 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_277
timestamp 1704896540
transform 1 0 26036 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_292
timestamp 1704896540
transform 1 0 27416 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_302
timestamp 1704896540
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_316
timestamp 1704896540
transform 1 0 29624 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_328
timestamp 1704896540
transform 1 0 30728 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_334
timestamp 1704896540
transform 1 0 31280 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1704896540
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_122
timestamp 1704896540
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1704896540
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_157
timestamp 1704896540
transform 1 0 14996 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_161
timestamp 1704896540
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_170
timestamp 1704896540
transform 1 0 16192 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_178
timestamp 1704896540
transform 1 0 16928 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_186
timestamp 1704896540
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_200
timestamp 1704896540
transform 1 0 18952 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_206
timestamp 1704896540
transform 1 0 19504 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_218
timestamp 1704896540
transform 1 0 20608 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_230
timestamp 1704896540
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_239
timestamp 1704896540
transform 1 0 22540 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1704896540
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1704896540
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_265
timestamp 1704896540
transform 1 0 24932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_272
timestamp 1704896540
transform 1 0 25576 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_280
timestamp 1704896540
transform 1 0 26312 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_289
timestamp 1704896540
transform 1 0 27140 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_300
timestamp 1704896540
transform 1 0 28152 0 1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1704896540
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_329
timestamp 1704896540
transform 1 0 30820 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1704896540
transform 1 0 5796 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1704896540
transform 1 0 6164 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_80
timestamp 1704896540
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1704896540
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_130
timestamp 1704896540
transform 1 0 12512 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_142
timestamp 1704896540
transform 1 0 13616 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_154
timestamp 1704896540
transform 1 0 14720 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1704896540
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_177
timestamp 1704896540
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_192
timestamp 1704896540
transform 1 0 18216 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_200
timestamp 1704896540
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 1704896540
transform 1 0 20240 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1704896540
transform 1 0 20976 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_233
timestamp 1704896540
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_245
timestamp 1704896540
transform 1 0 23092 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_251
timestamp 1704896540
transform 1 0 23644 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_268
timestamp 1704896540
transform 1 0 25208 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1704896540
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_287
timestamp 1704896540
transform 1 0 26956 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_299
timestamp 1704896540
transform 1 0 28060 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_313
timestamp 1704896540
transform 1 0 29348 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_327
timestamp 1704896540
transform 1 0 30636 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_45
timestamp 1704896540
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_60
timestamp 1704896540
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_128
timestamp 1704896540
transform 1 0 12328 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1704896540
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_141
timestamp 1704896540
transform 1 0 13524 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_158
timestamp 1704896540
transform 1 0 15088 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_171
timestamp 1704896540
transform 1 0 16284 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1704896540
transform 1 0 17480 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_209
timestamp 1704896540
transform 1 0 19780 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1704896540
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_233
timestamp 1704896540
transform 1 0 21988 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_239
timestamp 1704896540
transform 1 0 22540 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_247
timestamp 1704896540
transform 1 0 23276 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1704896540
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_253
timestamp 1704896540
transform 1 0 23828 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_269
timestamp 1704896540
transform 1 0 25300 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_277
timestamp 1704896540
transform 1 0 26036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_287
timestamp 1704896540
transform 1 0 26956 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_296
timestamp 1704896540
transform 1 0 27784 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_315
timestamp 1704896540
transform 1 0 29532 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_321
timestamp 1704896540
transform 1 0 30084 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_329
timestamp 1704896540
transform 1 0 30820 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_123
timestamp 1704896540
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_135
timestamp 1704896540
transform 1 0 12972 0 -1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_146
timestamp 1704896540
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_158
timestamp 1704896540
transform 1 0 15088 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1704896540
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_177
timestamp 1704896540
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_186
timestamp 1704896540
transform 1 0 17664 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_194
timestamp 1704896540
transform 1 0 18400 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_200
timestamp 1704896540
transform 1 0 18952 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1704896540
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_244
timestamp 1704896540
transform 1 0 23000 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_256
timestamp 1704896540
transform 1 0 24104 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_262
timestamp 1704896540
transform 1 0 24656 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_270
timestamp 1704896540
transform 1 0 25392 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1704896540
transform 1 0 26128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26404 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_291
timestamp 1704896540
transform 1 0 27324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_303
timestamp 1704896540
transform 1 0 28428 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_314
timestamp 1704896540
transform 1 0 29440 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1704896540
transform 1 0 30544 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_334
timestamp 1704896540
transform 1 0 31280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_23
timestamp 1704896540
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_61
timestamp 1704896540
transform 1 0 6164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_71
timestamp 1704896540
transform 1 0 7084 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_106
timestamp 1704896540
transform 1 0 10304 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_113
timestamp 1704896540
transform 1 0 10948 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_124
timestamp 1704896540
transform 1 0 11960 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_133
timestamp 1704896540
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1704896540
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_141
timestamp 1704896540
transform 1 0 13524 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_167
timestamp 1704896540
transform 1 0 15916 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_177
timestamp 1704896540
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_186
timestamp 1704896540
transform 1 0 17664 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1704896540
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1704896540
transform 1 0 18676 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_206
timestamp 1704896540
transform 1 0 19504 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_241
timestamp 1704896540
transform 1 0 22724 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 1704896540
transform 1 0 23552 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_256
timestamp 1704896540
transform 1 0 24104 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_266
timestamp 1704896540
transform 1 0 25024 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_290
timestamp 1704896540
transform 1 0 27232 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_302
timestamp 1704896540
transform 1 0 28336 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_317
timestamp 1704896540
transform 1 0 29716 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_332
timestamp 1704896540
transform 1 0 31096 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1704896540
transform 1 0 828 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_27
timestamp 1704896540
transform 1 0 3036 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1704896540
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1704896540
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_101
timestamp 1704896540
transform 1 0 9844 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_122
timestamp 1704896540
transform 1 0 11776 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_132
timestamp 1704896540
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_144
timestamp 1704896540
transform 1 0 13800 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_156
timestamp 1704896540
transform 1 0 14904 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_181
timestamp 1704896540
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_213
timestamp 1704896540
transform 1 0 20148 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1704896540
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1704896540
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_262
timestamp 1704896540
transform 1 0 24656 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_271
timestamp 1704896540
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1704896540
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_289
timestamp 1704896540
transform 1 0 27140 0 -1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_302
timestamp 1704896540
transform 1 0 28336 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_314
timestamp 1704896540
transform 1 0 29440 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_322
timestamp 1704896540
transform 1 0 30176 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_328
timestamp 1704896540
transform 1 0 30728 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_334
timestamp 1704896540
transform 1 0 31280 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 1704896540
transform 1 0 828 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_52
timestamp 1704896540
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_77
timestamp 1704896540
transform 1 0 7636 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_109
timestamp 1704896540
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1704896540
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_144
timestamp 1704896540
transform 1 0 13800 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_158
timestamp 1704896540
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_175
timestamp 1704896540
transform 1 0 16652 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 1704896540
transform 1 0 18124 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1704896540
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1704896540
transform 1 0 18676 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_209
timestamp 1704896540
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_218
timestamp 1704896540
transform 1 0 20608 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_229
timestamp 1704896540
transform 1 0 21620 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_241
timestamp 1704896540
transform 1 0 22724 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_249
timestamp 1704896540
transform 1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_253
timestamp 1704896540
transform 1 0 23828 0 1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1704896540
transform 1 0 24932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_277
timestamp 1704896540
transform 1 0 26036 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_285
timestamp 1704896540
transform 1 0 26772 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_295
timestamp 1704896540
transform 1 0 27692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1704896540
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_322
timestamp 1704896540
transform 1 0 30176 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_330
timestamp 1704896540
transform 1 0 30912 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_334
timestamp 1704896540
transform 1 0 31280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_26
timestamp 1704896540
transform 1 0 2944 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_42
timestamp 1704896540
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_69
timestamp 1704896540
transform 1 0 6900 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_93
timestamp 1704896540
transform 1 0 9108 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_122
timestamp 1704896540
transform 1 0 11776 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_140
timestamp 1704896540
transform 1 0 13432 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_146
timestamp 1704896540
transform 1 0 13984 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_153
timestamp 1704896540
transform 1 0 14628 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_157
timestamp 1704896540
transform 1 0 14996 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1704896540
transform 1 0 15824 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_176
timestamp 1704896540
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_188
timestamp 1704896540
transform 1 0 17848 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_194
timestamp 1704896540
transform 1 0 18400 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_206
timestamp 1704896540
transform 1 0 19504 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_212
timestamp 1704896540
transform 1 0 20056 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_216
timestamp 1704896540
transform 1 0 20424 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_232
timestamp 1704896540
transform 1 0 21896 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_238
timestamp 1704896540
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_253
timestamp 1704896540
transform 1 0 23828 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_257
timestamp 1704896540
transform 1 0 24196 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 1704896540
transform 1 0 25852 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1704896540
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_281
timestamp 1704896540
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_285
timestamp 1704896540
transform 1 0 26772 0 -1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_304
timestamp 1704896540
transform 1 0 28520 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_316
timestamp 1704896540
transform 1 0 29624 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_320
timestamp 1704896540
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_333
timestamp 1704896540
transform 1 0 31188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1704896540
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_109
timestamp 1704896540
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 1704896540
transform 1 0 10948 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_120
timestamp 1704896540
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1704896540
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_157
timestamp 1704896540
transform 1 0 14996 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_165
timestamp 1704896540
transform 1 0 15732 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_169
timestamp 1704896540
transform 1 0 16100 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_180
timestamp 1704896540
transform 1 0 17112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 1704896540
transform 1 0 18216 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_205
timestamp 1704896540
transform 1 0 19412 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_213
timestamp 1704896540
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_220
timestamp 1704896540
transform 1 0 20792 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_225
timestamp 1704896540
transform 1 0 21252 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1704896540
transform 1 0 21896 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1704896540
transform 1 0 23000 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_263
timestamp 1704896540
transform 1 0 24748 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_278
timestamp 1704896540
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_296
timestamp 1704896540
transform 1 0 27784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_302
timestamp 1704896540
transform 1 0 28336 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_321
timestamp 1704896540
transform 1 0 30084 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_326
timestamp 1704896540
transform 1 0 30544 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_334
timestamp 1704896540
transform 1 0 31280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27692 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 18308 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 28888 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 15088 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 19412 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 19780 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 19688 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform 1 0 12144 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform 1 0 10120 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 23552 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 4692 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 11684 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 4692 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 21620 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform 1 0 12880 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform -1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 10672 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 4508 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 6992 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 7360 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform 1 0 6348 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform -1 0 4784 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 10304 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 9936 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 8096 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 4508 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform 1 0 6992 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform -1 0 5888 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform 1 0 8464 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 10856 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 8464 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform -1 0 6532 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform -1 0 13616 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform 1 0 30268 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform 1 0 29808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 29532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform -1 0 28336 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform 1 0 27508 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform 1 0 27232 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform 1 0 26404 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1704896540
transform 1 0 25852 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform 1 0 24472 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  max_cap10
timestamp 1704896540
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap11
timestamp 1704896540
transform -1 0 7084 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1704896540
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1704896540
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1704896540
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1704896540
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1704896540
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1704896540
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1704896540
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1704896540
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1704896540
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1704896540
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1704896540
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1704896540
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1704896540
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1704896540
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1704896540
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1704896540
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1704896540
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1704896540
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1704896540
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1704896540
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1704896540
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1704896540
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1704896540
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1704896540
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1704896540
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1704896540
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1704896540
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1704896540
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1704896540
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1704896540
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1704896540
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1704896540
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1704896540
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1704896540
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1704896540
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1704896540
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1704896540
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1704896540
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1704896540
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1704896540
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1704896540
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1704896540
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1704896540
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1704896540
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1704896540
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1704896540
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1704896540
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1704896540
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1704896540
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1704896540
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1704896540
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1704896540
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1704896540
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1704896540
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1704896540
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1704896540
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1704896540
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1704896540
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1704896540
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1704896540
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1704896540
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1704896540
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1704896540
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1704896540
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1704896540
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1704896540
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1704896540
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1704896540
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1704896540
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1704896540
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1704896540
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1704896540
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1704896540
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1704896540
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1704896540
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1704896540
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1704896540
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1704896540
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1704896540
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1704896540
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1704896540
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1704896540
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1704896540
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1704896540
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1704896540
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1704896540
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1704896540
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1704896540
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1704896540
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1704896540
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1704896540
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1704896540
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1704896540
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1704896540
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1704896540
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1704896540
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1704896540
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1704896540
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1704896540
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1704896540
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1704896540
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1704896540
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1704896540
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1704896540
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1704896540
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1704896540
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1704896540
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1704896540
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1704896540
transform 1 0 28888 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 16180 21216 16180 21216 4 VGND
rlabel metal1 s 16100 21760 16100 21760 4 VPWR
rlabel metal1 s 22080 7276 22080 7276 4 DJ8.ACC\[0\]
rlabel metal2 s 22678 6817 22678 6817 4 DJ8.ACC\[1\]
rlabel metal2 s 21390 5797 21390 5797 4 DJ8.ACC\[2\]
rlabel metal1 s 13984 3706 13984 3706 4 DJ8.ACC\[3\]
rlabel metal3 s 18262 7480 18262 7480 4 DJ8.ACC\[4\]
rlabel metal4 s 6900 6732 6900 6732 4 DJ8.ACC\[5\]
rlabel metal2 s 6670 6936 6670 6936 4 DJ8.ACC\[6\]
rlabel metal2 s 13662 6851 13662 6851 4 DJ8.ACC\[7\]
rlabel metal1 s 20056 7514 20056 7514 4 DJ8.ALU.c_in
rlabel metal1 s 28658 6188 28658 6188 4 DJ8.ALU.opalu\[0\]
rlabel metal1 s 28842 6256 28842 6256 4 DJ8.ALU.opalu\[1\]
rlabel metal1 s 28934 5882 28934 5882 4 DJ8.ALU.opalu\[2\]
rlabel metal1 s 11822 8262 11822 8262 4 DJ8.EF\[0\]
rlabel metal1 s 5290 16116 5290 16116 4 DJ8.EF\[10\]
rlabel metal1 s 7958 16626 7958 16626 4 DJ8.EF\[11\]
rlabel metal1 s 6946 17782 6946 17782 4 DJ8.EF\[12\]
rlabel metal2 s 2898 17017 2898 17017 4 DJ8.EF\[13\]
rlabel metal2 s 3910 15657 3910 15657 4 DJ8.EF\[14\]
rlabel metal1 s 3059 14042 3059 14042 4 DJ8.EF\[15\]
rlabel metal2 s 12742 9010 12742 9010 4 DJ8.EF\[1\]
rlabel metal1 s 14674 11118 14674 11118 4 DJ8.EF\[2\]
rlabel metal1 s 7222 10982 7222 10982 4 DJ8.EF\[3\]
rlabel metal1 s 13800 8262 13800 8262 4 DJ8.EF\[4\]
rlabel metal1 s 3634 9520 3634 9520 4 DJ8.EF\[5\]
rlabel metal1 s 3772 12818 3772 12818 4 DJ8.EF\[6\]
rlabel metal1 s 4945 11866 4945 11866 4 DJ8.EF\[7\]
rlabel metal1 s 7682 13702 7682 13702 4 DJ8.EF\[8\]
rlabel metal2 s 7222 9350 7222 9350 4 DJ8.EF\[9\]
rlabel metal1 s 10764 9622 10764 9622 4 DJ8.GH\[0\]
rlabel metal1 s 2622 15028 2622 15028 4 DJ8.GH\[10\]
rlabel metal2 s 7774 16864 7774 16864 4 DJ8.GH\[11\]
rlabel metal1 s 10258 17748 10258 17748 4 DJ8.GH\[12\]
rlabel metal1 s 4002 17544 4002 17544 4 DJ8.GH\[13\]
rlabel metal2 s 5290 14654 5290 14654 4 DJ8.GH\[14\]
rlabel metal1 s 1932 14450 1932 14450 4 DJ8.GH\[15\]
rlabel metal1 s 15502 10438 15502 10438 4 DJ8.GH\[1\]
rlabel metal1 s 14812 11186 14812 11186 4 DJ8.GH\[2\]
rlabel metal1 s 9016 12410 9016 12410 4 DJ8.GH\[3\]
rlabel metal1 s 12834 10472 12834 10472 4 DJ8.GH\[4\]
rlabel metal1 s 5612 12682 5612 12682 4 DJ8.GH\[5\]
rlabel metal1 s 5878 13294 5878 13294 4 DJ8.GH\[6\]
rlabel metal1 s 2254 13464 2254 13464 4 DJ8.GH\[7\]
rlabel metal1 s 8418 13158 8418 13158 4 DJ8.GH\[8\]
rlabel metal1 s 7084 14586 7084 14586 4 DJ8.GH\[9\]
rlabel metal2 s 10350 5423 10350 5423 4 DJ8.REGS.regs\[1\]\[0\]
rlabel metal2 s 6854 6052 6854 6052 4 DJ8.REGS.regs\[1\]\[1\]
rlabel metal1 s 966 5644 966 5644 4 DJ8.REGS.regs\[1\]\[2\]
rlabel metal1 s 9936 2482 9936 2482 4 DJ8.REGS.regs\[1\]\[3\]
rlabel metal1 s 8418 3366 8418 3366 4 DJ8.REGS.regs\[1\]\[4\]
rlabel metal1 s 3082 4114 3082 4114 4 DJ8.REGS.regs\[1\]\[5\]
rlabel metal1 s 2530 4998 2530 4998 4 DJ8.REGS.regs\[1\]\[6\]
rlabel metal1 s 2162 5814 2162 5814 4 DJ8.REGS.regs\[1\]\[7\]
rlabel metal1 s 7360 6766 7360 6766 4 DJ8.REGS.regs\[2\]\[0\]
rlabel metal1 s 6532 4250 6532 4250 4 DJ8.REGS.regs\[2\]\[1\]
rlabel metal1 s 4232 10030 4232 10030 4 DJ8.REGS.regs\[2\]\[2\]
rlabel metal1 s 10097 3570 10097 3570 4 DJ8.REGS.regs\[2\]\[3\]
rlabel metal1 s 8556 4794 8556 4794 4 DJ8.REGS.regs\[2\]\[4\]
rlabel metal1 s 4140 7310 4140 7310 4 DJ8.REGS.regs\[2\]\[5\]
rlabel metal1 s 2852 11118 2852 11118 4 DJ8.REGS.regs\[2\]\[6\]
rlabel metal1 s 3289 10778 3289 10778 4 DJ8.REGS.regs\[2\]\[7\]
rlabel metal1 s 9614 6766 9614 6766 4 DJ8.REGS.regs\[3\]\[0\]
rlabel metal1 s 5704 6222 5704 6222 4 DJ8.REGS.regs\[3\]\[1\]
rlabel metal1 s 2070 6392 2070 6392 4 DJ8.REGS.regs\[3\]\[2\]
rlabel metal1 s 7498 6426 7498 6426 4 DJ8.REGS.regs\[3\]\[3\]
rlabel metal1 s 7452 8466 7452 8466 4 DJ8.REGS.regs\[3\]\[4\]
rlabel metal1 s 4232 8942 4232 8942 4 DJ8.REGS.regs\[3\]\[5\]
rlabel metal1 s 4048 7854 4048 7854 4 DJ8.REGS.regs\[3\]\[6\]
rlabel metal2 s 3726 7174 3726 7174 4 DJ8.REGS.regs\[3\]\[7\]
rlabel metal1 s 16238 9044 16238 9044 4 DJ8.REGS.write_addr\[0\]
rlabel metal1 s 17020 7310 17020 7310 4 DJ8.REGS.write_addr\[1\]
rlabel metal2 s 19366 13129 19366 13129 4 DJ8.REGS.write_addr\[2\]
rlabel metal2 s 15594 7752 15594 7752 4 DJ8.flag_Z
rlabel metal2 s 21574 10574 21574 10574 4 DJ8.ir\[0\]
rlabel metal1 s 21298 9690 21298 9690 4 DJ8.ir\[14\]
rlabel metal1 s 21298 9520 21298 9520 4 DJ8.ir\[15\]
rlabel metal1 s 22770 8908 22770 8908 4 DJ8.ir\[1\]
rlabel metal1 s 21574 10506 21574 10506 4 DJ8.ir\[2\]
rlabel metal1 s 19688 11118 19688 11118 4 DJ8.ir\[3\]
rlabel metal1 s 19918 10200 19918 10200 4 DJ8.ir\[4\]
rlabel metal1 s 15548 8942 15548 8942 4 DJ8.ir\[5\]
rlabel metal2 s 13662 13503 13662 13503 4 DJ8.ir\[6\]
rlabel metal2 s 12558 14705 12558 14705 4 DJ8.ir\[7\]
rlabel metal1 s 20608 11662 20608 11662 4 DJ8.pc\[0\]
rlabel metal2 s 10350 18564 10350 18564 4 DJ8.pc\[10\]
rlabel metal1 s 10672 18190 10672 18190 4 DJ8.pc\[11\]
rlabel metal1 s 2576 20230 2576 20230 4 DJ8.pc\[12\]
rlabel metal1 s 3818 19346 3818 19346 4 DJ8.pc\[13\]
rlabel metal1 s 2714 18394 2714 18394 4 DJ8.pc\[14\]
rlabel metal1 s 20102 12342 20102 12342 4 DJ8.pc\[1\]
rlabel metal1 s 15134 11866 15134 11866 4 DJ8.pc\[2\]
rlabel metal1 s 13754 11288 13754 11288 4 DJ8.pc\[3\]
rlabel metal1 s 13800 12886 13800 12886 4 DJ8.pc\[4\]
rlabel metal1 s 13616 13430 13616 13430 4 DJ8.pc\[5\]
rlabel metal2 s 8326 14178 8326 14178 4 DJ8.pc\[6\]
rlabel metal2 s 9154 13566 9154 13566 4 DJ8.pc\[7\]
rlabel metal1 s 7866 16150 7866 16150 4 DJ8.pc\[8\]
rlabel metal1 s 10718 17000 10718 17000 4 DJ8.pc\[9\]
rlabel metal1 s 26841 11866 26841 11866 4 DJ8.state\[0\]
rlabel metal1 s 18814 10098 18814 10098 4 DJ8.state\[1\]
rlabel metal1 s 26910 12750 26910 12750 4 DJ8.state\[2\]
rlabel metal1 s 17158 12954 17158 12954 4 DJ8.state\[3\]
rlabel metal1 s 13570 20400 13570 20400 4 DJ8.we
rlabel metal1 s 16054 12648 16054 12648 4 _0000_
rlabel metal2 s 17618 11917 17618 11917 4 _0001_
rlabel metal1 s 11822 9554 11822 9554 4 _0003_
rlabel metal1 s 9798 10200 9798 10200 4 _0004_
rlabel metal2 s 9338 9622 9338 9622 4 _0005_
rlabel metal2 s 7774 12036 7774 12036 4 _0006_
rlabel metal2 s 6026 11900 6026 11900 4 _0007_
rlabel metal1 s 1426 12410 1426 12410 4 _0008_
rlabel metal1 s 3956 12954 3956 12954 4 _0009_
rlabel metal2 s 1242 13668 1242 13668 4 _0010_
rlabel metal1 s 18078 9112 18078 9112 4 _0011_
rlabel metal1 s 16560 7990 16560 7990 4 _0012_
rlabel metal1 s 27600 10234 27600 10234 4 _0013_
rlabel metal1 s 28428 6970 28428 6970 4 _0014_
rlabel metal1 s 28198 6732 28198 6732 4 _0015_
rlabel metal1 s 27094 7208 27094 7208 4 _0016_
rlabel metal2 s 20010 9282 20010 9282 4 _0017_
rlabel metal1 s 23000 8602 23000 8602 4 _0018_
rlabel metal1 s 14076 6426 14076 6426 4 _0019_
rlabel metal1 s 13156 7242 13156 7242 4 _0020_
rlabel metal2 s 12834 6188 12834 6188 4 _0021_
rlabel metal1 s 11306 5338 11306 5338 4 _0022_
rlabel metal1 s 11454 3638 11454 3638 4 _0023_
rlabel metal1 s 10074 3026 10074 3026 4 _0024_
rlabel metal1 s 11362 4590 11362 4590 4 _0025_
rlabel metal2 s 10718 5304 10718 5304 4 _0026_
rlabel metal2 s 13110 5372 13110 5372 4 _0027_
rlabel metal1 s 8556 4250 8556 4250 4 _0028_
rlabel metal2 s 4738 6120 4738 6120 4 _0029_
rlabel metal2 s 2346 3332 2346 3332 4 _0030_
rlabel metal1 s 8464 3162 8464 3162 4 _0031_
rlabel metal1 s 6808 3162 6808 3162 4 _0032_
rlabel metal1 s 1472 3434 1472 3434 4 _0033_
rlabel metal1 s 1104 4250 1104 4250 4 _0034_
rlabel metal1 s 1196 4794 1196 4794 4 _0035_
rlabel metal1 s 7958 3162 7958 3162 4 _0036_
rlabel metal1 s 4728 4250 4728 4250 4 _0037_
rlabel metal1 s 2599 10166 2599 10166 4 _0038_
rlabel metal1 s 10074 4590 10074 4590 4 _0039_
rlabel metal1 s 6440 3366 6440 3366 4 _0040_
rlabel metal1 s 1104 4454 1104 4454 4 _0041_
rlabel metal1 s 1196 11322 1196 11322 4 _0042_
rlabel metal1 s 782 10234 782 10234 4 _0043_
rlabel metal1 s 8096 6902 8096 6902 4 _0044_
rlabel metal1 s 4232 3638 4232 3638 4 _0045_
rlabel metal1 s 2852 4726 2852 4726 4 _0046_
rlabel metal1 s 5612 6154 5612 6154 4 _0047_
rlabel metal1 s 5145 8602 5145 8602 4 _0048_
rlabel metal1 s 2576 8602 2576 8602 4 _0049_
rlabel metal1 s 2024 7990 2024 7990 4 _0050_
rlabel metal2 s 2806 5882 2806 5882 4 _0051_
rlabel metal1 s 5934 13498 5934 13498 4 _0052_
rlabel metal1 s 5152 14586 5152 14586 4 _0053_
rlabel metal1 s 1334 15606 1334 15606 4 _0054_
rlabel metal1 s 6026 16558 6026 16558 4 _0055_
rlabel metal1 s 6302 18122 6302 18122 4 _0056_
rlabel metal1 s 3128 17306 3128 17306 4 _0057_
rlabel metal1 s 3404 15130 3404 15130 4 _0058_
rlabel metal1 s 3910 13906 3910 13906 4 _0059_
rlabel metal1 s 11086 6698 11086 6698 4 _0060_
rlabel metal1 s 13938 9384 13938 9384 4 _0061_
rlabel metal1 s 13110 10200 13110 10200 4 _0062_
rlabel metal2 s 5566 10880 5566 10880 4 _0063_
rlabel metal1 s 11638 8058 11638 8058 4 _0064_
rlabel metal1 s 1932 9350 1932 9350 4 _0065_
rlabel metal1 s 2438 7446 2438 7446 4 _0066_
rlabel metal1 s 3358 11662 3358 11662 4 _0067_
rlabel metal1 s 6670 13294 6670 13294 4 _0068_
rlabel metal1 s 5060 14042 5060 14042 4 _0069_
rlabel metal1 s 3634 15470 3634 15470 4 _0070_
rlabel metal1 s 5881 17306 5881 17306 4 _0071_
rlabel metal2 s 10994 18530 10994 18530 4 _0072_
rlabel metal1 s 1196 17306 1196 17306 4 _0073_
rlabel metal1 s 1196 16218 1196 16218 4 _0074_
rlabel metal1 s 1334 14586 1334 14586 4 _0075_
rlabel metal1 s 18492 7242 18492 7242 4 _0076_
rlabel metal2 s 25714 10336 25714 10336 4 _0077_
rlabel metal1 s 27140 8942 27140 8942 4 _0078_
rlabel metal1 s 28244 8602 28244 8602 4 _0079_
rlabel metal1 s 26128 10234 26128 10234 4 _0080_
rlabel metal1 s 23368 10166 23368 10166 4 _0081_
rlabel metal1 s 24787 8602 24787 8602 4 _0082_
rlabel metal1 s 24932 7990 24932 7990 4 _0083_
rlabel metal1 s 20654 8330 20654 8330 4 _0084_
rlabel metal1 s 1196 18938 1196 18938 4 _0085_
rlabel metal2 s 3082 19652 3082 19652 4 _0086_
rlabel metal1 s 2047 18258 2047 18258 4 _0087_
rlabel metal1 s 14582 13158 14582 13158 4 _0088_
rlabel metal2 s 16146 10863 16146 10863 4 _0089_
rlabel metal1 s 19964 10642 19964 10642 4 _0090_
rlabel metal1 s 13202 11866 13202 11866 4 _0091_
rlabel metal1 s 12098 11866 12098 11866 4 _0092_
rlabel metal1 s 11454 12682 11454 12682 4 _0093_
rlabel metal2 s 11960 13294 11960 13294 4 _0094_
rlabel metal1 s 11723 14042 11723 14042 4 _0095_
rlabel metal2 s 10258 15300 10258 15300 4 _0096_
rlabel metal1 s 7636 15402 7636 15402 4 _0097_
rlabel metal1 s 9775 16082 9775 16082 4 _0098_
rlabel metal2 s 9706 17680 9706 17680 4 _0099_
rlabel metal1 s 8924 17306 8924 17306 4 _0100_
rlabel metal1 s 7268 20434 7268 20434 4 _0101_
rlabel metal1 s 5934 19958 5934 19958 4 _0102_
rlabel metal1 s 8786 21080 8786 21080 4 _0103_
rlabel metal1 s 3726 21114 3726 21114 4 _0104_
rlabel metal1 s 3404 20298 3404 20298 4 _0105_
rlabel metal1 s 1196 19958 1196 19958 4 _0106_
rlabel metal1 s 1196 18598 1196 18598 4 _0107_
rlabel metal2 s 2714 21012 2714 21012 4 _0108_
rlabel metal1 s 3082 6222 3082 6222 4 _0109_
rlabel metal1 s 8050 13838 8050 13838 4 _0110_
rlabel metal1 s 6210 13260 6210 13260 4 _0111_
rlabel metal1 s 5750 14450 5750 14450 4 _0112_
rlabel metal1 s 1012 15538 1012 15538 4 _0113_
rlabel metal1 s 5566 16626 5566 16626 4 _0114_
rlabel metal1 s 6072 17850 6072 17850 4 _0115_
rlabel metal1 s 3266 17102 3266 17102 4 _0116_
rlabel metal1 s 3542 14948 3542 14948 4 _0117_
rlabel metal1 s 2990 13498 2990 13498 4 _0118_
rlabel metal2 s 9476 11322 9476 11322 4 _0119_
rlabel metal1 s 1518 9010 1518 9010 4 _0120_
rlabel metal1 s 10764 6834 10764 6834 4 _0121_
rlabel metal2 s 12374 9316 12374 9316 4 _0122_
rlabel metal1 s 12650 9384 12650 9384 4 _0123_
rlabel metal1 s 5520 10574 5520 10574 4 _0124_
rlabel metal2 s 10994 8619 10994 8619 4 _0125_
rlabel metal1 s 3082 9486 3082 9486 4 _0126_
rlabel metal2 s 2898 7701 2898 7701 4 _0127_
rlabel metal1 s 3082 11322 3082 11322 4 _0128_
rlabel metal1 s 10350 13362 10350 13362 4 _0129_
rlabel metal3 s 10534 13141 10534 13141 4 _0130_
rlabel metal1 s 6762 12954 6762 12954 4 _0131_
rlabel metal1 s 5290 13838 5290 13838 4 _0132_
rlabel metal1 s 3266 15538 3266 15538 4 _0133_
rlabel metal1 s 8556 16150 8556 16150 4 _0134_
rlabel metal1 s 7958 17850 7958 17850 4 _0135_
rlabel metal1 s 1472 17102 1472 17102 4 _0136_
rlabel metal1 s 1472 16014 1472 16014 4 _0137_
rlabel metal1 s 1656 14450 1656 14450 4 _0138_
rlabel metal1 s 15962 5032 15962 5032 4 _0139_
rlabel metal1 s 18124 5814 18124 5814 4 _0140_
rlabel metal1 s 17710 4794 17710 4794 4 _0141_
rlabel metal1 s 18216 5882 18216 5882 4 _0142_
rlabel metal2 s 17894 6902 17894 6902 4 _0143_
rlabel metal1 s 17250 6426 17250 6426 4 _0144_
rlabel metal1 s 18400 6902 18400 6902 4 _0145_
rlabel metal1 s 18492 7310 18492 7310 4 _0146_
rlabel metal1 s 25668 10098 25668 10098 4 _0147_
rlabel metal1 s 26266 9010 26266 9010 4 _0148_
rlabel metal1 s 27600 8398 27600 8398 4 _0149_
rlabel metal1 s 25990 10132 25990 10132 4 _0150_
rlabel metal1 s 24196 10098 24196 10098 4 _0151_
rlabel metal1 s 25116 9010 25116 9010 4 _0152_
rlabel metal1 s 23644 8602 23644 8602 4 _0153_
rlabel metal1 s 20562 9010 20562 9010 4 _0154_
rlabel metal1 s 10028 12274 10028 12274 4 _0155_
rlabel metal1 s 9246 13770 9246 13770 4 _0156_
rlabel metal1 s 8372 17102 8372 17102 4 _0157_
rlabel metal1 s 7406 17510 7406 17510 4 _0158_
rlabel metal2 s 10902 17765 10902 17765 4 _0159_
rlabel metal1 s 3680 18394 3680 18394 4 _0160_
rlabel metal1 s 17388 9690 17388 9690 4 _0161_
rlabel metal2 s 5106 17153 5106 17153 4 _0162_
rlabel metal1 s 2990 18938 2990 18938 4 _0163_
rlabel metal1 s 17756 8602 17756 8602 4 _0164_
rlabel metal2 s 17894 9505 17894 9505 4 _0165_
rlabel metal2 s 2530 18785 2530 18785 4 _0166_
rlabel metal1 s 1518 18802 1518 18802 4 _0167_
rlabel metal1 s 4278 18258 4278 18258 4 _0168_
rlabel metal1 s 5796 18802 5796 18802 4 _0169_
rlabel metal1 s 4554 18938 4554 18938 4 _0170_
rlabel metal1 s 4048 18938 4048 18938 4 _0171_
rlabel metal1 s 3726 19176 3726 19176 4 _0172_
rlabel metal1 s 9384 14926 9384 14926 4 _0173_
rlabel metal2 s 4554 17051 4554 17051 4 _0174_
rlabel metal1 s 4278 17102 4278 17102 4 _0175_
rlabel metal1 s 4186 17306 4186 17306 4 _0176_
rlabel metal1 s 3082 18292 3082 18292 4 _0177_
rlabel metal1 s 18032 10778 18032 10778 4 _0178_
rlabel metal2 s 18262 13889 18262 13889 4 _0179_
rlabel metal2 s 17158 12478 17158 12478 4 _0180_
rlabel metal1 s 16744 10778 16744 10778 4 _0181_
rlabel metal1 s 16882 11220 16882 11220 4 _0182_
rlabel metal1 s 15134 10234 15134 10234 4 _0183_
rlabel metal1 s 16100 10234 16100 10234 4 _0184_
rlabel metal1 s 18630 10778 18630 10778 4 _0185_
rlabel metal1 s 17710 11084 17710 11084 4 _0186_
rlabel metal1 s 9821 14450 9821 14450 4 _0187_
rlabel metal1 s 10442 11696 10442 11696 4 _0188_
rlabel metal2 s 10258 10948 10258 10948 4 _0189_
rlabel metal1 s 9706 11628 9706 11628 4 _0190_
rlabel metal1 s 9246 17680 9246 17680 4 _0191_
rlabel metal1 s 12650 11628 12650 11628 4 _0192_
rlabel metal1 s 10718 10234 10718 10234 4 _0193_
rlabel metal1 s 10259 12240 10259 12240 4 _0194_
rlabel metal1 s 11546 11730 11546 11730 4 _0195_
rlabel metal1 s 9614 12784 9614 12784 4 _0196_
rlabel metal2 s 9504 12750 9504 12750 4 _0197_
rlabel metal1 s 10534 12784 10534 12784 4 _0198_
rlabel metal1 s 10212 13430 10212 13430 4 _0199_
rlabel metal1 s 9752 13294 9752 13294 4 _0200_
rlabel metal1 s 10442 12410 10442 12410 4 _0201_
rlabel metal1 s 9890 13770 9890 13770 4 _0202_
rlabel metal2 s 8694 14960 8694 14960 4 _0203_
rlabel metal1 s 9890 13838 9890 13838 4 _0204_
rlabel metal1 s 10810 14042 10810 14042 4 _0205_
rlabel metal2 s 9062 13906 9062 13906 4 _0206_
rlabel metal1 s 8952 14450 8952 14450 4 _0207_
rlabel metal1 s 9476 14586 9476 14586 4 _0208_
rlabel metal2 s 8786 17510 8786 17510 4 _0209_
rlabel metal1 s 10856 17034 10856 17034 4 _0210_
rlabel metal1 s 12144 16218 12144 16218 4 _0211_
rlabel metal1 s 9890 15572 9890 15572 4 _0212_
rlabel metal2 s 10534 16575 10534 16575 4 _0213_
rlabel metal1 s 6624 15674 6624 15674 4 _0214_
rlabel metal1 s 10074 16660 10074 16660 4 _0215_
rlabel metal2 s 10994 16983 10994 16983 4 _0216_
rlabel metal1 s 12098 17612 12098 17612 4 _0217_
rlabel metal1 s 10442 17136 10442 17136 4 _0218_
rlabel metal1 s 10350 17816 10350 17816 4 _0219_
rlabel metal2 s 10533 17714 10533 17714 4 _0220_
rlabel metal1 s 9614 17136 9614 17136 4 _0221_
rlabel metal2 s 16330 20774 16330 20774 4 _0222_
rlabel metal1 s 16008 20978 16008 20978 4 _0223_
rlabel metal1 s 1886 20400 1886 20400 4 _0224_
rlabel metal1 s 6762 21114 6762 21114 4 _0225_
rlabel metal1 s 6302 19176 6302 19176 4 _0226_
rlabel metal1 s 8694 21454 8694 21454 4 _0227_
rlabel metal1 s 3358 21012 3358 21012 4 _0228_
rlabel metal1 s 3082 20944 3082 20944 4 _0229_
rlabel metal1 s 1104 20366 1104 20366 4 _0230_
rlabel metal1 s 966 18836 966 18836 4 _0231_
rlabel metal1 s 3082 20468 3082 20468 4 _0232_
rlabel metal2 s 15824 17204 15824 17204 4 _0233_
rlabel metal2 s 11730 13362 11730 13362 4 _0234_
rlabel metal1 s 18538 9078 18538 9078 4 _0235_
rlabel metal1 s 16698 11662 16698 11662 4 _0236_
rlabel metal1 s 19550 12172 19550 12172 4 _0237_
rlabel metal1 s 16974 12240 16974 12240 4 _0238_
rlabel metal1 s 18124 12682 18124 12682 4 _0239_
rlabel metal3 s 18446 12971 18446 12971 4 _0240_
rlabel metal2 s 19274 11373 19274 11373 4 _0241_
rlabel metal1 s 9246 14348 9246 14348 4 _0242_
rlabel metal1 s 19136 11322 19136 11322 4 _0243_
rlabel metal1 s 20286 11560 20286 11560 4 _0244_
rlabel metal2 s 21206 11067 21206 11067 4 _0245_
rlabel metal2 s 20378 11781 20378 11781 4 _0246_
rlabel metal1 s 13754 14450 13754 14450 4 _0247_
rlabel metal1 s 9016 14994 9016 14994 4 _0248_
rlabel metal1 s 11868 15674 11868 15674 4 _0249_
rlabel metal1 s 7682 14586 7682 14586 4 _0250_
rlabel metal1 s 8648 15130 8648 15130 4 _0251_
rlabel metal1 s 11546 15946 11546 15946 4 _0252_
rlabel metal1 s 11408 16218 11408 16218 4 _0253_
rlabel metal2 s 8142 17527 8142 17527 4 _0254_
rlabel metal1 s 9982 18938 9982 18938 4 _0255_
rlabel metal1 s 8602 18938 8602 18938 4 _0256_
rlabel metal1 s 9246 19210 9246 19210 4 _0257_
rlabel metal2 s 4830 19040 4830 19040 4 _0258_
rlabel metal1 s 5750 18870 5750 18870 4 _0259_
rlabel metal2 s 5658 18768 5658 18768 4 _0260_
rlabel metal1 s 6118 19346 6118 19346 4 _0261_
rlabel metal1 s 17756 12206 17756 12206 4 _0262_
rlabel metal1 s 10258 3978 10258 3978 4 _0263_
rlabel metal1 s 8326 6766 8326 6766 4 _0264_
rlabel metal4 s 9821 6052 9821 6052 4 _0265_
rlabel metal1 s 10212 6630 10212 6630 4 _0266_
rlabel metal1 s 8119 8330 8119 8330 4 _0267_
rlabel metal1 s 10306 6222 10306 6222 4 _0268_
rlabel metal2 s 6118 6205 6118 6205 4 _0269_
rlabel metal1 s 10258 6120 10258 6120 4 _0270_
rlabel metal2 s 9522 4624 9522 4624 4 _0271_
rlabel metal1 s 8740 10506 8740 10506 4 _0272_
rlabel metal1 s 8050 10574 8050 10574 4 _0273_
rlabel metal1 s 9614 6222 9614 6222 4 _0274_
rlabel metal1 s 10258 6426 10258 6426 4 _0275_
rlabel metal3 s 7613 6052 7613 6052 4 _0276_
rlabel metal1 s 5129 9486 5129 9486 4 _0277_
rlabel metal1 s 4600 8330 4600 8330 4 _0278_
rlabel metal1 s 10396 7922 10396 7922 4 _0279_
rlabel metal2 s 9982 7378 9982 7378 4 _0280_
rlabel metal1 s 20286 7820 20286 7820 4 _0281_
rlabel metal2 s 21850 9282 21850 9282 4 _0282_
rlabel metal1 s 21850 12308 21850 12308 4 _0283_
rlabel metal1 s 21459 11118 21459 11118 4 _0284_
rlabel metal1 s 20608 10982 20608 10982 4 _0285_
rlabel metal1 s 20838 12138 20838 12138 4 _0286_
rlabel metal1 s 21206 12716 21206 12716 4 _0287_
rlabel metal2 s 19458 12920 19458 12920 4 _0288_
rlabel metal1 s 16330 11526 16330 11526 4 _0289_
rlabel metal2 s 14766 12699 14766 12699 4 _0290_
rlabel metal1 s 11408 20366 11408 20366 4 _0291_
rlabel metal1 s 6716 7310 6716 7310 4 _0292_
rlabel metal1 s 6164 7514 6164 7514 4 _0293_
rlabel metal1 s 7130 7888 7130 7888 4 _0294_
rlabel metal1 s 6854 7378 6854 7378 4 _0295_
rlabel metal1 s 6670 19142 6670 19142 4 _0296_
rlabel metal1 s 19412 11594 19412 11594 4 _0297_
rlabel metal2 s 22770 13039 22770 13039 4 _0298_
rlabel metal3 s 23782 12291 23782 12291 4 _0299_
rlabel metal1 s 19826 12274 19826 12274 4 _0300_
rlabel metal1 s 23736 10506 23736 10506 4 _0301_
rlabel metal2 s 24426 11594 24426 11594 4 _0302_
rlabel metal2 s 11454 19652 11454 19652 4 _0303_
rlabel metal1 s 10902 19278 10902 19278 4 _0304_
rlabel metal2 s 4922 10438 4922 10438 4 _0305_
rlabel metal2 s 5290 10659 5290 10659 4 _0306_
rlabel metal1 s 10672 11050 10672 11050 4 _0307_
rlabel metal2 s 1564 5882 1564 5882 4 _0308_
rlabel metal2 s 1058 7123 1058 7123 4 _0309_
rlabel metal3 s 11523 18972 11523 18972 4 _0310_
rlabel metal2 s 19550 11084 19550 11084 4 _0311_
rlabel metal1 s 20792 14042 20792 14042 4 _0312_
rlabel metal2 s 14030 12478 14030 12478 4 _0313_
rlabel metal2 s 20286 12002 20286 12002 4 _0314_
rlabel metal1 s 22724 12274 22724 12274 4 _0315_
rlabel metal1 s 22218 12410 22218 12410 4 _0316_
rlabel metal1 s 20930 13804 20930 13804 4 _0317_
rlabel metal1 s 30360 15538 30360 15538 4 _0318_
rlabel metal1 s 30222 17102 30222 17102 4 _0319_
rlabel metal1 s 10856 19890 10856 19890 4 _0320_
rlabel metal1 s 9062 7378 9062 7378 4 _0321_
rlabel metal1 s 9890 6834 9890 6834 4 _0322_
rlabel metal1 s 8234 7344 8234 7344 4 _0323_
rlabel metal2 s 10074 6902 10074 6902 4 _0324_
rlabel metal1 s 20608 7990 20608 7990 4 _0325_
rlabel metal1 s 15732 12886 15732 12886 4 _0326_
rlabel metal2 s 13662 12223 13662 12223 4 _0327_
rlabel metal2 s 19642 12988 19642 12988 4 _0328_
rlabel metal1 s 15180 16014 15180 16014 4 _0329_
rlabel metal1 s 13018 17714 13018 17714 4 _0330_
rlabel metal1 s 12374 18054 12374 18054 4 _0331_
rlabel metal1 s 9108 20366 9108 20366 4 _0332_
rlabel metal2 s 8050 6681 8050 6681 4 _0333_
rlabel metal1 s 8372 6426 8372 6426 4 _0334_
rlabel metal1 s 7590 9452 7590 9452 4 _0335_
rlabel metal1 s 9292 7922 9292 7922 4 _0336_
rlabel metal2 s 19366 6205 19366 6205 4 _0337_
rlabel metal1 s 16146 14484 16146 14484 4 _0338_
rlabel metal1 s 13386 13838 13386 13838 4 _0339_
rlabel metal1 s 14122 14042 14122 14042 4 _0340_
rlabel metal2 s 14398 14518 14398 14518 4 _0341_
rlabel metal1 s 30222 14450 30222 14450 4 _0342_
rlabel metal1 s 13018 16524 13018 16524 4 _0343_
rlabel metal1 s 18768 18190 18768 18190 4 _0344_
rlabel metal2 s 10534 21012 10534 21012 4 _0345_
rlabel metal1 s 4646 9146 4646 9146 4 _0346_
rlabel metal2 s 5290 8636 5290 8636 4 _0347_
rlabel metal1 s 4278 6256 4278 6256 4 _0348_
rlabel metal1 s 5060 6426 5060 6426 4 _0349_
rlabel metal1 s 1702 20434 1702 20434 4 _0350_
rlabel metal1 s 15962 13906 15962 13906 4 _0351_
rlabel metal2 s 6578 10081 6578 10081 4 _0352_
rlabel metal1 s 15686 13430 15686 13430 4 _0353_
rlabel metal1 s 17618 13770 17618 13770 4 _0354_
rlabel metal1 s 15824 14926 15824 14926 4 _0355_
rlabel metal1 s 26542 17068 26542 17068 4 _0356_
rlabel metal1 s 9706 20230 9706 20230 4 _0357_
rlabel metal1 s 8096 19278 8096 19278 4 _0358_
rlabel metal1 s 4784 11186 4784 11186 4 _0359_
rlabel metal1 s 5980 7922 5980 7922 4 _0360_
rlabel metal1 s 4186 6800 4186 6800 4 _0361_
rlabel metal1 s 4968 6970 4968 6970 4 _0362_
rlabel metal1 s 1978 18666 1978 18666 4 _0363_
rlabel metal3 s 8050 12852 8050 12852 4 _0364_
rlabel metal1 s 12328 14382 12328 14382 4 _0365_
rlabel metal1 s 21620 14382 21620 14382 4 _0366_
rlabel metal2 s 10994 20876 10994 20876 4 _0367_
rlabel metal1 s 10166 21352 10166 21352 4 _0368_
rlabel metal1 s 4278 12614 4278 12614 4 _0369_
rlabel metal1 s 5198 6630 5198 6630 4 _0370_
rlabel metal1 s 1380 5610 1380 5610 4 _0371_
rlabel metal1 s 5382 6868 5382 6868 4 _0372_
rlabel metal3 s 19366 7939 19366 7939 4 _0373_
rlabel metal1 s 5290 12070 5290 12070 4 _0374_
rlabel metal2 s 12466 14212 12466 14212 4 _0375_
rlabel metal2 s 16974 18683 16974 18683 4 _0376_
rlabel metal1 s 9108 20842 9108 20842 4 _0377_
rlabel metal1 s 3634 14586 3634 14586 4 _0378_
rlabel metal1 s 14168 20978 14168 20978 4 _0379_
rlabel metal1 s 14214 20910 14214 20910 4 _0380_
rlabel metal1 s 14260 21658 14260 21658 4 _0381_
rlabel metal1 s 14168 21114 14168 21114 4 _0382_
rlabel metal1 s 14214 21352 14214 21352 4 _0383_
rlabel metal1 s 14260 21454 14260 21454 4 _0384_
rlabel metal2 s 24425 6222 24425 6222 4 _0385_
rlabel metal2 s 24334 9044 24334 9044 4 _0386_
rlabel metal1 s 19090 6732 19090 6732 4 _0387_
rlabel metal1 s 25392 12070 25392 12070 4 _0388_
rlabel metal1 s 23966 12206 23966 12206 4 _0389_
rlabel metal1 s 25116 16694 25116 16694 4 _0390_
rlabel metal2 s 15226 20978 15226 20978 4 _0391_
rlabel metal2 s 20838 13090 20838 13090 4 _0392_
rlabel metal1 s 18906 13362 18906 13362 4 _0393_
rlabel metal2 s 22126 13158 22126 13158 4 _0394_
rlabel metal1 s 22310 16422 22310 16422 4 _0395_
rlabel metal2 s 21022 13464 21022 13464 4 _0396_
rlabel metal1 s 19504 14586 19504 14586 4 _0397_
rlabel metal1 s 20378 20973 20378 20973 4 _0398_
rlabel metal1 s 30912 13362 30912 13362 4 _0399_
rlabel metal1 s 20976 20366 20976 20366 4 _0400_
rlabel metal1 s 27922 21046 27922 21046 4 _0401_
rlabel metal1 s 19458 14484 19458 14484 4 _0402_
rlabel metal2 s 16790 14654 16790 14654 4 _0403_
rlabel metal1 s 30498 17000 30498 17000 4 _0404_
rlabel metal1 s 22448 18802 22448 18802 4 _0405_
rlabel metal1 s 20700 12750 20700 12750 4 _0406_
rlabel metal1 s 18998 12716 18998 12716 4 _0407_
rlabel metal1 s 20194 13736 20194 13736 4 _0408_
rlabel metal1 s 18538 14382 18538 14382 4 _0409_
rlabel metal1 s 26818 14960 26818 14960 4 _0410_
rlabel metal2 s 21850 13923 21850 13923 4 _0411_
rlabel metal1 s 27370 17068 27370 17068 4 _0412_
rlabel metal1 s 27324 16626 27324 16626 4 _0413_
rlabel metal1 s 27922 17306 27922 17306 4 _0414_
rlabel metal1 s 26910 19924 26910 19924 4 _0415_
rlabel metal1 s 26680 15674 26680 15674 4 _0416_
rlabel metal2 s 21022 20332 21022 20332 4 _0417_
rlabel metal1 s 28014 20944 28014 20944 4 _0418_
rlabel metal1 s 27139 20366 27139 20366 4 _0419_
rlabel metal1 s 16238 14926 16238 14926 4 _0420_
rlabel metal2 s 30406 14994 30406 14994 4 _0421_
rlabel metal1 s 28060 19754 28060 19754 4 _0422_
rlabel metal1 s 25990 13362 25990 13362 4 _0423_
rlabel metal1 s 14168 19278 14168 19278 4 _0424_
rlabel metal1 s 20562 13328 20562 13328 4 _0425_
rlabel metal1 s 18722 13464 18722 13464 4 _0426_
rlabel metal1 s 24794 12750 24794 12750 4 _0427_
rlabel metal1 s 24564 12954 24564 12954 4 _0428_
rlabel metal1 s 27646 14484 27646 14484 4 _0429_
rlabel metal1 s 27094 14348 27094 14348 4 _0430_
rlabel metal1 s 27232 12750 27232 12750 4 _0431_
rlabel metal1 s 27922 14416 27922 14416 4 _0432_
rlabel metal1 s 27232 14246 27232 14246 4 _0433_
rlabel metal2 s 20654 14144 20654 14144 4 _0434_
rlabel metal2 s 15962 20417 15962 20417 4 _0435_
rlabel metal1 s 21390 14926 21390 14926 4 _0436_
rlabel metal2 s 11868 19822 11868 19822 4 _0437_
rlabel metal1 s 20424 14586 20424 14586 4 _0438_
rlabel metal1 s 24656 15606 24656 15606 4 _0439_
rlabel metal1 s 30038 12716 30038 12716 4 _0440_
rlabel metal1 s 15916 14314 15916 14314 4 _0441_
rlabel metal1 s 21390 14586 21390 14586 4 _0442_
rlabel metal2 s 26818 14620 26818 14620 4 _0443_
rlabel metal1 s 26680 14586 26680 14586 4 _0444_
rlabel metal3 s 14628 16184 14628 16184 4 _0445_
rlabel metal1 s 22632 19822 22632 19822 4 _0446_
rlabel metal2 s 17434 18428 17434 18428 4 _0447_
rlabel metal1 s 15502 20230 15502 20230 4 _0448_
rlabel metal2 s 21574 20077 21574 20077 4 _0449_
rlabel metal1 s 23598 12954 23598 12954 4 _0450_
rlabel metal1 s 23874 18190 23874 18190 4 _0451_
rlabel metal1 s 25852 16490 25852 16490 4 _0452_
rlabel metal1 s 24610 19856 24610 19856 4 _0453_
rlabel metal2 s 30222 17799 30222 17799 4 _0454_
rlabel metal1 s 23736 19958 23736 19958 4 _0455_
rlabel metal1 s 24104 14994 24104 14994 4 _0456_
rlabel metal1 s 19136 19482 19136 19482 4 _0457_
rlabel metal1 s 20148 19482 20148 19482 4 _0458_
rlabel metal1 s 25024 19754 25024 19754 4 _0459_
rlabel metal1 s 26726 17646 26726 17646 4 _0460_
rlabel metal2 s 14950 14603 14950 14603 4 _0461_
rlabel metal1 s 26864 19210 26864 19210 4 _0462_
rlabel metal1 s 26910 17034 26910 17034 4 _0463_
rlabel metal1 s 30682 15912 30682 15912 4 _0464_
rlabel metal2 s 30222 16592 30222 16592 4 _0465_
rlabel metal1 s 22494 16966 22494 16966 4 _0466_
rlabel metal1 s 27140 17306 27140 17306 4 _0467_
rlabel metal2 s 26910 19108 26910 19108 4 _0468_
rlabel metal1 s 26680 19482 26680 19482 4 _0469_
rlabel metal1 s 27140 20026 27140 20026 4 _0470_
rlabel metal2 s 16974 8687 16974 8687 4 _0471_
rlabel metal1 s 25300 9418 25300 9418 4 _0472_
rlabel metal2 s 23598 7276 23598 7276 4 _0473_
rlabel metal1 s 22218 5780 22218 5780 4 _0474_
rlabel metal1 s 23138 5100 23138 5100 4 _0475_
rlabel metal1 s 23138 14586 23138 14586 4 _0476_
rlabel metal2 s 14766 15725 14766 15725 4 _0477_
rlabel metal1 s 23230 14892 23230 14892 4 _0478_
rlabel metal1 s 25438 14994 25438 14994 4 _0479_
rlabel metal1 s 26542 15470 26542 15470 4 _0480_
rlabel metal1 s 29808 13362 29808 13362 4 _0481_
rlabel metal1 s 30268 13362 30268 13362 4 _0482_
rlabel metal3 s 16974 20349 16974 20349 4 _0483_
rlabel metal1 s 29026 13328 29026 13328 4 _0484_
rlabel metal1 s 28796 14450 28796 14450 4 _0485_
rlabel metal1 s 25622 12206 25622 12206 4 _0486_
rlabel metal1 s 27830 13498 27830 13498 4 _0487_
rlabel metal2 s 25346 14365 25346 14365 4 _0488_
rlabel metal1 s 26082 15606 26082 15606 4 _0489_
rlabel metal1 s 25024 14994 25024 14994 4 _0490_
rlabel metal1 s 26588 15130 26588 15130 4 _0491_
rlabel metal1 s 29762 15674 29762 15674 4 _0492_
rlabel metal1 s 19826 12886 19826 12886 4 _0493_
rlabel metal1 s 24748 13770 24748 13770 4 _0494_
rlabel metal1 s 28934 15130 28934 15130 4 _0495_
rlabel metal1 s 29486 15504 29486 15504 4 _0496_
rlabel metal1 s 28014 15470 28014 15470 4 _0497_
rlabel metal2 s 26864 14926 26864 14926 4 _0498_
rlabel metal1 s 27232 15334 27232 15334 4 _0499_
rlabel metal1 s 24380 15946 24380 15946 4 _0500_
rlabel metal1 s 25806 15470 25806 15470 4 _0501_
rlabel metal1 s 26450 15538 26450 15538 4 _0502_
rlabel metal1 s 27508 15606 27508 15606 4 _0503_
rlabel metal1 s 27784 15674 27784 15674 4 _0504_
rlabel metal2 s 16790 7616 16790 7616 4 _0505_
rlabel metal1 s 24748 7310 24748 7310 4 _0506_
rlabel metal1 s 23966 7276 23966 7276 4 _0507_
rlabel metal2 s 25806 6834 25806 6834 4 _0508_
rlabel metal1 s 25576 8058 25576 8058 4 _0509_
rlabel metal1 s 24058 7344 24058 7344 4 _0510_
rlabel metal1 s 25438 6222 25438 6222 4 _0511_
rlabel metal1 s 24426 5032 24426 5032 4 _0512_
rlabel metal1 s 23644 4658 23644 4658 4 _0513_
rlabel metal2 s 18262 6868 18262 6868 4 _0514_
rlabel metal1 s 18400 6766 18400 6766 4 _0515_
rlabel metal2 s 19734 12908 19734 12908 4 _0516_
rlabel metal2 s 20562 3264 20562 3264 4 _0517_
rlabel metal2 s 25714 4114 25714 4114 4 _0518_
rlabel metal2 s 24242 6086 24242 6086 4 _0519_
rlabel metal1 s 24150 6766 24150 6766 4 _0520_
rlabel metal1 s 25208 6222 25208 6222 4 _0521_
rlabel metal1 s 26174 5542 26174 5542 4 _0522_
rlabel metal1 s 26788 4726 26788 4726 4 _0523_
rlabel metal1 s 26680 4522 26680 4522 4 _0524_
rlabel metal2 s 20562 4590 20562 4590 4 _0525_
rlabel metal1 s 24380 3366 24380 3366 4 _0526_
rlabel metal1 s 29302 5134 29302 5134 4 _0527_
rlabel metal2 s 29670 4726 29670 4726 4 _0528_
rlabel metal1 s 21666 3672 21666 3672 4 _0529_
rlabel metal1 s 29486 5066 29486 5066 4 _0530_
rlabel metal1 s 26634 4080 26634 4080 4 _0531_
rlabel metal1 s 27140 4998 27140 4998 4 _0532_
rlabel metal1 s 27094 5746 27094 5746 4 _0533_
rlabel metal1 s 19550 4012 19550 4012 4 _0534_
rlabel metal2 s 26634 5372 26634 5372 4 _0535_
rlabel metal1 s 26082 5134 26082 5134 4 _0536_
rlabel metal2 s 26909 4046 26909 4046 4 _0537_
rlabel metal1 s 25254 5202 25254 5202 4 _0538_
rlabel metal1 s 25254 5270 25254 5270 4 _0539_
rlabel metal1 s 24288 4658 24288 4658 4 _0540_
rlabel metal1 s 22448 5610 22448 5610 4 _0541_
rlabel metal1 s 23322 4692 23322 4692 4 _0542_
rlabel metal1 s 23138 4590 23138 4590 4 _0543_
rlabel metal1 s 18262 6222 18262 6222 4 _0544_
rlabel metal1 s 23966 4624 23966 4624 4 _0545_
rlabel metal2 s 16606 4641 16606 4641 4 _0546_
rlabel metal1 s 14628 6290 14628 6290 4 _0547_
rlabel metal1 s 14904 5746 14904 5746 4 _0548_
rlabel metal1 s 15502 5780 15502 5780 4 _0549_
rlabel metal2 s 15042 4794 15042 4794 4 _0550_
rlabel metal1 s 21758 4658 21758 4658 4 _0551_
rlabel metal1 s 20194 2618 20194 2618 4 _0552_
rlabel metal1 s 25070 6188 25070 6188 4 _0553_
rlabel metal1 s 24518 6256 24518 6256 4 _0554_
rlabel metal2 s 22126 5712 22126 5712 4 _0555_
rlabel metal1 s 21942 4658 21942 4658 4 _0556_
rlabel metal1 s 22402 4692 22402 4692 4 _0557_
rlabel metal1 s 21804 5134 21804 5134 4 _0558_
rlabel metal1 s 7866 13736 7866 13736 4 _0559_
rlabel metal1 s 16928 8398 16928 8398 4 _0560_
rlabel metal1 s 17250 7174 17250 7174 4 _0561_
rlabel metal1 s 8418 13872 8418 13872 4 _0562_
rlabel metal1 s 8510 9078 8510 9078 4 _0563_
rlabel metal2 s 9798 10914 9798 10914 4 _0564_
rlabel metal1 s 10488 9350 10488 9350 4 _0565_
rlabel metal1 s 12006 16592 12006 16592 4 _0566_
rlabel metal2 s 15410 20723 15410 20723 4 _0567_
rlabel metal1 s 20079 15946 20079 15946 4 _0568_
rlabel metal1 s 19366 16218 19366 16218 4 _0569_
rlabel metal1 s 18722 17306 18722 17306 4 _0570_
rlabel metal1 s 12558 18292 12558 18292 4 _0571_
rlabel metal1 s 12880 17102 12880 17102 4 _0572_
rlabel metal2 s 16974 18020 16974 18020 4 _0573_
rlabel metal1 s 17940 15674 17940 15674 4 _0574_
rlabel metal2 s 12098 16575 12098 16575 4 _0575_
rlabel metal1 s 17020 17306 17020 17306 4 _0576_
rlabel metal1 s 17342 18394 17342 18394 4 _0577_
rlabel metal3 s 17687 19516 17687 19516 4 _0578_
rlabel metal2 s 17802 19074 17802 19074 4 _0579_
rlabel metal1 s 17250 20468 17250 20468 4 _0580_
rlabel metal1 s 17618 20434 17618 20434 4 _0581_
rlabel metal2 s 16974 19754 16974 19754 4 _0582_
rlabel metal1 s 17158 18836 17158 18836 4 _0583_
rlabel metal3 s 19780 18904 19780 18904 4 _0584_
rlabel metal2 s 14766 16303 14766 16303 4 _0585_
rlabel metal1 s 29302 16660 29302 16660 4 _0586_
rlabel metal1 s 29164 18802 29164 18802 4 _0587_
rlabel metal1 s 20102 16660 20102 16660 4 _0588_
rlabel metal2 s 28750 17187 28750 17187 4 _0589_
rlabel metal2 s 28934 18224 28934 18224 4 _0590_
rlabel metal1 s 29026 18836 29026 18836 4 _0591_
rlabel metal1 s 16560 20230 16560 20230 4 _0592_
rlabel metal1 s 29348 18938 29348 18938 4 _0593_
rlabel metal1 s 23046 20230 23046 20230 4 _0594_
rlabel metal1 s 11684 19278 11684 19278 4 _0595_
rlabel metal1 s 30820 20570 30820 20570 4 _0596_
rlabel metal1 s 29670 21114 29670 21114 4 _0597_
rlabel metal2 s 28796 20196 28796 20196 4 _0598_
rlabel metal2 s 29394 20298 29394 20298 4 _0599_
rlabel metal2 s 29072 18972 29072 18972 4 _0600_
rlabel metal2 s 27462 6052 27462 6052 4 _0601_
rlabel metal2 s 25898 5338 25898 5338 4 _0602_
rlabel metal1 s 27738 3502 27738 3502 4 _0603_
rlabel metal1 s 26956 4658 26956 4658 4 _0604_
rlabel metal1 s 25208 4590 25208 4590 4 _0605_
rlabel metal1 s 23092 4046 23092 4046 4 _0606_
rlabel metal1 s 23460 4114 23460 4114 4 _0607_
rlabel metal1 s 24104 3162 24104 3162 4 _0608_
rlabel metal1 s 23506 4012 23506 4012 4 _0609_
rlabel metal1 s 26174 4658 26174 4658 4 _0610_
rlabel metal1 s 27186 4658 27186 4658 4 _0611_
rlabel metal1 s 27646 3978 27646 3978 4 _0612_
rlabel metal1 s 26496 3706 26496 3706 4 _0613_
rlabel metal3 s 27186 4029 27186 4029 4 _0614_
rlabel metal1 s 27830 4182 27830 4182 4 _0615_
rlabel metal1 s 26128 4046 26128 4046 4 _0616_
rlabel metal1 s 28106 4182 28106 4182 4 _0617_
rlabel metal1 s 24012 4046 24012 4046 4 _0618_
rlabel metal3 s 13938 4709 13938 4709 4 _0619_
rlabel metal1 s 5980 14586 5980 14586 4 _0620_
rlabel metal1 s 8648 9622 8648 9622 4 _0621_
rlabel metal1 s 20976 17306 20976 17306 4 _0622_
rlabel metal1 s 14766 18156 14766 18156 4 _0623_
rlabel metal1 s 21482 17748 21482 17748 4 _0624_
rlabel metal1 s 19182 15436 19182 15436 4 _0625_
rlabel metal1 s 18124 15470 18124 15470 4 _0626_
rlabel metal2 s 18998 15521 18998 15521 4 _0627_
rlabel metal1 s 18906 15674 18906 15674 4 _0628_
rlabel metal1 s 14674 16456 14674 16456 4 _0629_
rlabel metal1 s 17388 15674 17388 15674 4 _0630_
rlabel metal1 s 18906 16116 18906 16116 4 _0631_
rlabel metal1 s 20332 16150 20332 16150 4 _0632_
rlabel metal2 s 21390 17068 21390 17068 4 _0633_
rlabel metal1 s 14628 16626 14628 16626 4 _0634_
rlabel metal1 s 13754 16762 13754 16762 4 _0635_
rlabel metal1 s 12926 16524 12926 16524 4 _0636_
rlabel metal2 s 13202 17034 13202 17034 4 _0637_
rlabel metal1 s 12466 16966 12466 16966 4 _0638_
rlabel metal1 s 22264 15606 22264 15606 4 _0639_
rlabel metal1 s 16560 14586 16560 14586 4 _0640_
rlabel metal1 s 13110 15402 13110 15402 4 _0641_
rlabel metal1 s 12834 15572 12834 15572 4 _0642_
rlabel metal1 s 11822 16694 11822 16694 4 _0643_
rlabel metal2 s 13202 15980 13202 15980 4 _0644_
rlabel metal2 s 12558 16388 12558 16388 4 _0645_
rlabel metal3 s 12006 17051 12006 17051 4 _0646_
rlabel metal2 s 22034 19380 22034 19380 4 _0647_
rlabel metal2 s 21114 14727 21114 14727 4 _0648_
rlabel metal1 s 20976 7310 20976 7310 4 _0649_
rlabel metal1 s 21482 1836 21482 1836 4 _0650_
rlabel metal1 s 21114 1870 21114 1870 4 _0651_
rlabel metal1 s 25070 2414 25070 2414 4 _0652_
rlabel metal1 s 24242 2516 24242 2516 4 _0653_
rlabel metal1 s 23414 2890 23414 2890 4 _0654_
rlabel metal1 s 25806 2618 25806 2618 4 _0655_
rlabel metal2 s 26450 2652 26450 2652 4 _0656_
rlabel metal1 s 27324 2346 27324 2346 4 _0657_
rlabel metal1 s 26266 2550 26266 2550 4 _0658_
rlabel metal1 s 26266 2074 26266 2074 4 _0659_
rlabel metal1 s 25116 2346 25116 2346 4 _0660_
rlabel metal1 s 23598 2448 23598 2448 4 _0661_
rlabel metal2 s 23322 3332 23322 3332 4 _0662_
rlabel metal1 s 25484 2074 25484 2074 4 _0663_
rlabel metal1 s 25254 2074 25254 2074 4 _0664_
rlabel metal3 s 21022 3587 21022 3587 4 _0665_
rlabel metal1 s 25254 3060 25254 3060 4 _0666_
rlabel metal1 s 25300 2550 25300 2550 4 _0667_
rlabel metal1 s 25116 2958 25116 2958 4 _0668_
rlabel metal2 s 25714 3298 25714 3298 4 _0669_
rlabel metal1 s 22954 3026 22954 3026 4 _0670_
rlabel metal2 s 14306 2621 14306 2621 4 _0671_
rlabel metal1 s 3036 15878 3036 15878 4 _0672_
rlabel metal1 s 9660 10438 9660 10438 4 _0673_
rlabel metal1 s 14306 19448 14306 19448 4 _0674_
rlabel metal1 s 12052 18258 12052 18258 4 _0675_
rlabel metal1 s 14352 18190 14352 18190 4 _0676_
rlabel metal1 s 13662 18258 13662 18258 4 _0677_
rlabel metal1 s 15916 18190 15916 18190 4 _0678_
rlabel metal1 s 14030 18156 14030 18156 4 _0679_
rlabel metal1 s 14628 16218 14628 16218 4 _0680_
rlabel metal1 s 14030 17136 14030 17136 4 _0681_
rlabel metal1 s 14168 17306 14168 17306 4 _0682_
rlabel metal1 s 14766 18258 14766 18258 4 _0683_
rlabel metal1 s 23414 16660 23414 16660 4 _0684_
rlabel metal1 s 22816 16082 22816 16082 4 _0685_
rlabel metal1 s 23276 15946 23276 15946 4 _0686_
rlabel metal1 s 22586 16082 22586 16082 4 _0687_
rlabel metal1 s 23000 16218 23000 16218 4 _0688_
rlabel metal2 s 22954 19958 22954 19958 4 _0689_
rlabel metal1 s 23644 19142 23644 19142 4 _0690_
rlabel metal1 s 16514 21046 16514 21046 4 _0691_
rlabel metal1 s 23920 19686 23920 19686 4 _0692_
rlabel metal1 s 22908 18190 22908 18190 4 _0693_
rlabel metal1 s 26312 18122 26312 18122 4 _0694_
rlabel metal1 s 21758 6834 21758 6834 4 _0695_
rlabel metal1 s 19067 6834 19067 6834 4 _0696_
rlabel metal1 s 20010 3570 20010 3570 4 _0697_
rlabel metal2 s 19090 5712 19090 5712 4 _0698_
rlabel metal2 s 19734 1632 19734 1632 4 _0699_
rlabel metal2 s 21942 2278 21942 2278 4 _0700_
rlabel metal1 s 22402 2380 22402 2380 4 _0701_
rlabel metal1 s 15686 2448 15686 2448 4 _0702_
rlabel metal1 s 22540 2618 22540 2618 4 _0703_
rlabel metal2 s 22034 2652 22034 2652 4 _0704_
rlabel metal2 s 20838 1802 20838 1802 4 _0705_
rlabel metal1 s 20470 1870 20470 1870 4 _0706_
rlabel metal1 s 20378 2006 20378 2006 4 _0707_
rlabel metal1 s 21206 2074 21206 2074 4 _0708_
rlabel metal2 s 18630 6528 18630 6528 4 _0709_
rlabel metal1 s 21620 2958 21620 2958 4 _0710_
rlabel metal1 s 21714 3570 21714 3570 4 _0711_
rlabel metal1 s 21298 3604 21298 3604 4 _0712_
rlabel metal1 s 21850 3026 21850 3026 4 _0713_
rlabel metal2 s 21620 2550 21620 2550 4 _0714_
rlabel metal1 s 21666 2482 21666 2482 4 _0715_
rlabel metal2 s 14214 1972 14214 1972 4 _0716_
rlabel metal1 s 14996 2890 14996 2890 4 _0717_
rlabel metal1 s 8188 12614 8188 12614 4 _0718_
rlabel metal3 s 25438 20995 25438 20995 4 _0719_
rlabel metal1 s 23276 20774 23276 20774 4 _0720_
rlabel metal2 s 19090 21284 19090 21284 4 _0721_
rlabel metal1 s 23460 20978 23460 20978 4 _0722_
rlabel metal1 s 23000 20570 23000 20570 4 _0723_
rlabel metal1 s 24242 20910 24242 20910 4 _0724_
rlabel metal1 s 24978 20570 24978 20570 4 _0725_
rlabel metal1 s 24794 20978 24794 20978 4 _0726_
rlabel metal1 s 24886 18258 24886 18258 4 _0727_
rlabel metal1 s 27416 12954 27416 12954 4 _0728_
rlabel metal1 s 26312 18190 26312 18190 4 _0729_
rlabel metal1 s 24656 18394 24656 18394 4 _0730_
rlabel metal1 s 24242 21114 24242 21114 4 _0731_
rlabel metal2 s 20286 21284 20286 21284 4 _0732_
rlabel metal2 s 15778 21267 15778 21267 4 _0733_
rlabel metal1 s 17802 21454 17802 21454 4 _0734_
rlabel metal1 s 14490 19482 14490 19482 4 _0735_
rlabel metal1 s 15824 19482 15824 19482 4 _0736_
rlabel metal1 s 14766 20230 14766 20230 4 _0737_
rlabel metal1 s 15226 19278 15226 19278 4 _0738_
rlabel metal1 s 14720 19482 14720 19482 4 _0739_
rlabel metal1 s 14720 20570 14720 20570 4 _0740_
rlabel metal1 s 17066 21556 17066 21556 4 _0741_
rlabel metal1 s 24886 21386 24886 21386 4 _0742_
rlabel metal2 s 25944 21420 25944 21420 4 _0743_
rlabel metal1 s 20884 6698 20884 6698 4 _0744_
rlabel metal1 s 16974 2516 16974 2516 4 _0745_
rlabel metal2 s 19642 2481 19642 2481 4 _0746_
rlabel metal1 s 16422 2414 16422 2414 4 _0747_
rlabel metal1 s 17388 2074 17388 2074 4 _0748_
rlabel metal1 s 15870 2511 15870 2511 4 _0749_
rlabel metal1 s 14950 2074 14950 2074 4 _0750_
rlabel metal1 s 15594 2550 15594 2550 4 _0751_
rlabel metal1 s 19412 1190 19412 1190 4 _0752_
rlabel metal1 s 17342 2006 17342 2006 4 _0753_
rlabel metal1 s 17986 1802 17986 1802 4 _0754_
rlabel metal1 s 19090 1394 19090 1394 4 _0755_
rlabel metal1 s 19136 1530 19136 1530 4 _0756_
rlabel metal1 s 17894 2380 17894 2380 4 _0757_
rlabel metal1 s 18722 2618 18722 2618 4 _0758_
rlabel metal2 s 19090 2652 19090 2652 4 _0759_
rlabel metal1 s 19734 2822 19734 2822 4 _0760_
rlabel metal1 s 20654 3706 20654 3706 4 _0761_
rlabel metal1 s 16882 3026 16882 3026 4 _0762_
rlabel metal2 s 20470 3604 20470 3604 4 _0763_
rlabel metal1 s 19826 3026 19826 3026 4 _0764_
rlabel metal1 s 19320 2822 19320 2822 4 _0765_
rlabel metal1 s 15134 2380 15134 2380 4 _0766_
rlabel metal1 s 15640 2618 15640 2618 4 _0767_
rlabel metal1 s 14490 3502 14490 3502 4 _0768_
rlabel metal1 s 14260 8262 14260 8262 4 _0769_
rlabel metal1 s 6164 12274 6164 12274 4 _0770_
rlabel metal2 s 29946 19924 29946 19924 4 _0771_
rlabel metal1 s 28842 19890 28842 19890 4 _0772_
rlabel metal1 s 24610 19244 24610 19244 4 _0773_
rlabel metal1 s 24564 17782 24564 17782 4 _0774_
rlabel metal1 s 24196 17782 24196 17782 4 _0775_
rlabel metal1 s 24610 17578 24610 17578 4 _0776_
rlabel metal1 s 26128 16762 26128 16762 4 _0777_
rlabel metal1 s 26174 17578 26174 17578 4 _0778_
rlabel metal1 s 25346 17646 25346 17646 4 _0779_
rlabel metal1 s 25116 17850 25116 17850 4 _0780_
rlabel metal1 s 12282 18326 12282 18326 4 _0781_
rlabel metal2 s 11822 18462 11822 18462 4 _0782_
rlabel metal1 s 11454 18394 11454 18394 4 _0783_
rlabel metal1 s 11592 18734 11592 18734 4 _0784_
rlabel metal1 s 12029 19210 12029 19210 4 _0785_
rlabel metal1 s 11546 18904 11546 18904 4 _0786_
rlabel metal3 s 11086 18683 11086 18683 4 _0787_
rlabel metal1 s 30314 17680 30314 17680 4 _0788_
rlabel metal2 s 30314 15266 30314 15266 4 _0789_
rlabel metal1 s 30728 17306 30728 17306 4 _0790_
rlabel metal1 s 30544 17714 30544 17714 4 _0791_
rlabel metal2 s 29946 18292 29946 18292 4 _0792_
rlabel metal1 s 25254 18700 25254 18700 4 _0793_
rlabel metal1 s 24748 18938 24748 18938 4 _0794_
rlabel metal3 s 19826 8483 19826 8483 4 _0795_
rlabel metal2 s 20467 4658 20467 4658 4 _0796_
rlabel metal1 s 16974 4726 16974 4726 4 _0797_
rlabel metal1 s 16974 4080 16974 4080 4 _0798_
rlabel metal1 s 17158 4012 17158 4012 4 _0799_
rlabel metal1 s 17618 3502 17618 3502 4 _0800_
rlabel metal1 s 16698 3434 16698 3434 4 _0801_
rlabel metal1 s 15226 3570 15226 3570 4 _0802_
rlabel metal1 s 15088 3706 15088 3706 4 _0803_
rlabel metal1 s 17756 2618 17756 2618 4 _0804_
rlabel metal1 s 17618 2958 17618 2958 4 _0805_
rlabel metal1 s 17894 4556 17894 4556 4 _0806_
rlabel metal1 s 17572 3570 17572 3570 4 _0807_
rlabel metal1 s 18124 2482 18124 2482 4 _0808_
rlabel metal1 s 18078 4182 18078 4182 4 _0809_
rlabel metal1 s 17572 4046 17572 4046 4 _0810_
rlabel metal1 s 16652 4182 16652 4182 4 _0811_
rlabel metal2 s 19182 4284 19182 4284 4 _0812_
rlabel metal2 s 19458 4250 19458 4250 4 _0813_
rlabel metal1 s 15824 4046 15824 4046 4 _0814_
rlabel metal2 s 15686 4386 15686 4386 4 _0815_
rlabel metal1 s 15502 4590 15502 4590 4 _0816_
rlabel metal1 s 14306 4080 14306 4080 4 _0817_
rlabel metal1 s 2300 16966 2300 16966 4 _0818_
rlabel metal1 s 1886 12274 1886 12274 4 _0819_
rlabel metal1 s 15226 5066 15226 5066 4 _0820_
rlabel metal1 s 22540 18938 22540 18938 4 _0821_
rlabel metal1 s 21574 19176 21574 19176 4 _0822_
rlabel metal1 s 21344 19278 21344 19278 4 _0823_
rlabel metal2 s 21298 20570 21298 20570 4 _0824_
rlabel metal2 s 20102 20060 20102 20060 4 _0825_
rlabel metal1 s 19964 19890 19964 19890 4 _0826_
rlabel metal2 s 19826 20128 19826 20128 4 _0827_
rlabel metal1 s 19136 19754 19136 19754 4 _0828_
rlabel metal2 s 20838 19482 20838 19482 4 _0829_
rlabel metal2 s 20378 19210 20378 19210 4 _0830_
rlabel metal1 s 19456 18258 19456 18258 4 _0831_
rlabel metal2 s 19550 18547 19550 18547 4 _0832_
rlabel metal1 s 20470 18803 20470 18803 4 _0833_
rlabel metal1 s 19274 18768 19274 18768 4 _0834_
rlabel metal1 s 20470 18598 20470 18598 4 _0835_
rlabel metal1 s 19964 16762 19964 16762 4 _0836_
rlabel metal1 s 19642 16626 19642 16626 4 _0837_
rlabel metal1 s 19412 16490 19412 16490 4 _0838_
rlabel metal1 s 19872 17714 19872 17714 4 _0839_
rlabel metal1 s 20378 17578 20378 17578 4 _0840_
rlabel metal1 s 20930 18700 20930 18700 4 _0841_
rlabel metal1 s 20608 19278 20608 19278 4 _0842_
rlabel metal2 s 20654 9469 20654 9469 4 _0843_
rlabel metal1 s 18354 5746 18354 5746 4 _0844_
rlabel metal1 s 17388 6834 17388 6834 4 _0845_
rlabel metal1 s 17618 6256 17618 6256 4 _0846_
rlabel metal1 s 17894 6222 17894 6222 4 _0847_
rlabel metal1 s 16974 5134 16974 5134 4 _0848_
rlabel metal1 s 16514 5678 16514 5678 4 _0849_
rlabel metal1 s 16008 5270 16008 5270 4 _0850_
rlabel metal1 s 15962 5134 15962 5134 4 _0851_
rlabel metal2 s 17158 5202 17158 5202 4 _0852_
rlabel metal1 s 17802 4692 17802 4692 4 _0853_
rlabel metal2 s 18170 4964 18170 4964 4 _0854_
rlabel metal2 s 18078 5440 18078 5440 4 _0855_
rlabel metal1 s 20010 5882 20010 5882 4 _0856_
rlabel metal2 s 19642 5712 19642 5712 4 _0857_
rlabel metal1 s 19826 5168 19826 5168 4 _0858_
rlabel metal1 s 18354 5236 18354 5236 4 _0859_
rlabel metal1 s 17112 5066 17112 5066 4 _0860_
rlabel metal1 s 15157 5338 15157 5338 4 _0861_
rlabel metal1 s 14352 4794 14352 4794 4 _0862_
rlabel metal1 s 14536 4250 14536 4250 4 _0863_
rlabel metal2 s 14214 5780 14214 5780 4 _0864_
rlabel metal1 s 3588 12750 3588 12750 4 _0865_
rlabel metal1 s 14904 4794 14904 4794 4 _0866_
rlabel metal2 s 2162 13872 2162 13872 4 _0867_
rlabel metal1 s 1656 13362 1656 13362 4 _0868_
rlabel metal2 s 17434 9044 17434 9044 4 _0869_
rlabel metal1 s 17664 7446 17664 7446 4 _0870_
rlabel metal1 s 27232 10098 27232 10098 4 _0871_
rlabel metal1 s 28750 6834 28750 6834 4 _0872_
rlabel metal1 s 29118 6834 29118 6834 4 _0873_
rlabel metal2 s 26266 6528 26266 6528 4 _0874_
rlabel metal1 s 20056 9010 20056 9010 4 _0875_
rlabel metal1 s 23000 8398 23000 8398 4 _0876_
rlabel metal1 s 18262 9894 18262 9894 4 _0877_
rlabel metal1 s 15364 8398 15364 8398 4 _0878_
rlabel metal1 s 14858 6358 14858 6358 4 _0879_
rlabel metal1 s 14076 6222 14076 6222 4 _0880_
rlabel metal1 s 11086 7344 11086 7344 4 _0881_
rlabel metal1 s 12190 6868 12190 6868 4 _0882_
rlabel metal2 s 12650 7242 12650 7242 4 _0883_
rlabel metal2 s 12466 7174 12466 7174 4 _0884_
rlabel metal1 s 9798 5780 9798 5780 4 _0885_
rlabel metal1 s 10672 5134 10672 5134 4 _0886_
rlabel metal1 s 11454 3162 11454 3162 4 _0887_
rlabel metal1 s 9154 4046 9154 4046 4 _0888_
rlabel metal1 s 10948 4250 10948 4250 4 _0889_
rlabel metal1 s 10672 4658 10672 4658 4 _0890_
rlabel metal1 s 13294 4726 13294 4726 4 _0891_
rlabel metal1 s 9062 5814 9062 5814 4 _0892_
rlabel metal1 s 7682 3026 7682 3026 4 _0893_
rlabel metal1 s 8050 4080 8050 4080 4 _0894_
rlabel metal1 s 5428 5610 5428 5610 4 _0895_
rlabel metal1 s 3128 2958 3128 2958 4 _0896_
rlabel metal1 s 8740 2958 8740 2958 4 _0897_
rlabel metal1 s 6992 2958 6992 2958 4 _0898_
rlabel metal1 s 1794 3162 1794 3162 4 _0899_
rlabel metal1 s 966 4046 966 4046 4 _0900_
rlabel metal1 s 1012 4658 1012 4658 4 _0901_
rlabel metal2 s 9614 9826 9614 9826 4 _0902_
rlabel metal1 s 7544 5678 7544 5678 4 _0903_
rlabel metal1 s 8096 2958 8096 2958 4 _0904_
rlabel metal1 s 4784 4658 4784 4658 4 _0905_
rlabel metal1 s 3128 10574 3128 10574 4 _0906_
rlabel metal1 s 9936 4182 9936 4182 4 _0907_
rlabel metal1 s 6118 3570 6118 3570 4 _0908_
rlabel metal1 s 1564 4658 1564 4658 4 _0909_
rlabel metal1 s 1564 11186 1564 11186 4 _0910_
rlabel metal1 s 1288 10098 1288 10098 4 _0911_
rlabel metal1 s 10764 6766 10764 6766 4 _0912_
rlabel metal1 s 11868 9010 11868 9010 4 _0913_
rlabel metal2 s 9062 6528 9062 6528 4 _0914_
rlabel metal1 s 7820 6358 7820 6358 4 _0915_
rlabel metal1 s 4462 4012 4462 4012 4 _0916_
rlabel metal1 s 3174 5134 3174 5134 4 _0917_
rlabel metal1 s 6670 5848 6670 5848 4 _0918_
rlabel metal1 s 5704 9010 5704 9010 4 _0919_
rlabel metal1 s 3082 8398 3082 8398 4 _0920_
rlabel metal1 s 506 7616 506 7616 4 _0921_
rlabel metal2 s 20746 15436 20746 15436 4 clk
rlabel metal1 s 21758 11186 21758 11186 4 clknet_0_clk
rlabel metal1 s 2530 4692 2530 4692 4 clknet_3_0__leaf_clk
rlabel metal1 s 9890 3060 9890 3060 4 clknet_3_1__leaf_clk
rlabel metal1 s 2714 17782 2714 17782 4 clknet_3_2__leaf_clk
rlabel metal1 s 12466 19924 12466 19924 4 clknet_3_3__leaf_clk
rlabel metal1 s 15272 7786 15272 7786 4 clknet_3_4__leaf_clk
rlabel metal1 s 15088 10778 15088 10778 4 clknet_3_5__leaf_clk
rlabel metal1 s 29394 10132 29394 10132 4 clknet_3_6__leaf_clk
rlabel metal2 s 19274 9010 19274 9010 4 clknet_3_7__leaf_clk
rlabel metal3 s 30199 20740 30199 20740 4 net1
rlabel metal2 s 2622 5984 2622 5984 4 net10
rlabel metal2 s 4094 16320 4094 16320 4 net11
rlabel metal1 s 6578 4454 6578 4454 4 net12
rlabel metal1 s 7261 6222 7261 6222 4 net13
rlabel metal1 s 7222 7242 7222 7242 4 net14
rlabel metal2 s 9154 6018 9154 6018 4 net15
rlabel metal1 s 16698 10438 16698 10438 4 net16
rlabel metal2 s 12742 11305 12742 11305 4 net17
rlabel metal1 s 4699 16626 4699 16626 4 net18
rlabel metal1 s 8333 16694 8333 16694 4 net19
rlabel metal1 s 28060 20434 28060 20434 4 net2
rlabel metal1 s 2629 18122 2629 18122 4 net20
rlabel metal1 s 6907 20298 6907 20298 4 net21
rlabel metal1 s 12719 20774 12719 20774 4 net22
rlabel metal1 s 28711 10166 28711 10166 4 net23
rlabel metal2 s 25806 9452 25806 9452 4 net24
rlabel metal1 s 20339 10506 20339 10506 4 net25
rlabel metal1 s 17303 12682 17303 12682 4 net26
rlabel metal1 s 12880 20026 12880 20026 4 net27
rlabel metal1 s 27094 11730 27094 11730 4 net28
rlabel metal2 s 17618 12517 17618 12517 4 net29
rlabel metal2 s 27554 18768 27554 18768 4 net3
rlabel metal1 s 29348 10030 29348 10030 4 net30
rlabel metal1 s 14122 7922 14122 7922 4 net31
rlabel metal2 s 18722 14467 18722 14467 4 net32
rlabel metal1 s 18814 10166 18814 10166 4 net33
rlabel metal2 s 18998 11407 18998 11407 4 net34
rlabel metal2 s 12558 11662 12558 11662 4 net35
rlabel metal1 s 10120 14586 10120 14586 4 net36
rlabel metal1 s 10672 14994 10672 14994 4 net37
rlabel metal2 s 19826 11441 19826 11441 4 net38
rlabel metal1 s 3726 8500 3726 8500 4 net39
rlabel metal1 s 29486 19244 29486 19244 4 net4
rlabel metal1 s 9522 16524 9522 16524 4 net40
rlabel metal1 s 3864 10234 3864 10234 4 net41
rlabel metal2 s 20930 10217 20930 10217 4 net42
rlabel metal1 s 13708 11730 13708 11730 4 net43
rlabel metal1 s 3956 5134 3956 5134 4 net44
rlabel metal1 s 11086 5882 11086 5882 4 net45
rlabel metal1 s 2346 11186 2346 11186 4 net46
rlabel metal1 s 9660 3706 9660 3706 4 net47
rlabel metal1 s 3726 7412 3726 7412 4 net48
rlabel metal2 s 6302 6256 6302 6256 4 net49
rlabel metal1 s 27232 21590 27232 21590 4 net5
rlabel metal1 s 6486 8602 6486 8602 4 net50
rlabel metal1 s 7314 3978 7314 3978 4 net51
rlabel metal2 s 2806 7038 2806 7038 4 net52
rlabel metal1 s 9430 2618 9430 2618 4 net53
rlabel metal1 s 9062 6086 9062 6086 4 net54
rlabel metal1 s 7268 5882 7268 5882 4 net55
rlabel metal1 s 3772 3162 3772 3162 4 net56
rlabel metal1 s 7728 5882 7728 5882 4 net57
rlabel metal1 s 5290 5882 5290 5882 4 net58
rlabel metal1 s 9246 15538 9246 15538 4 net59
rlabel metal1 s 27002 18258 27002 18258 4 net6
rlabel metal1 s 9108 17102 9108 17102 4 net60
rlabel metal1 s 7636 2618 7636 2618 4 net61
rlabel metal2 s 5842 3910 5842 3910 4 net62
rlabel metal1 s 12673 7786 12673 7786 4 net63
rlabel metal1 s 25990 21590 25990 21590 4 net7
rlabel metal1 s 25438 19278 25438 19278 4 net8
rlabel metal1 s 23046 21590 23046 21590 4 net9
rlabel metal4 s 30268 22001 30268 22001 4 rst_n
rlabel metal4 s 29532 22001 29532 22001 4 ui_in[0]
rlabel metal4 s 28796 22069 28796 22069 4 ui_in[1]
rlabel metal4 s 28060 22001 28060 22001 4 ui_in[2]
rlabel metal4 s 27324 21865 27324 21865 4 ui_in[3]
rlabel metal4 s 26588 21933 26588 21933 4 ui_in[4]
rlabel metal4 s 25852 22001 25852 22001 4 ui_in[5]
rlabel metal4 s 25116 22069 25116 22069 4 ui_in[6]
rlabel metal4 s 24380 22001 24380 22001 4 ui_in[7]
rlabel metal3 s 6486 21131 6486 21131 4 uio_oe[0]
rlabel metal3 s 6670 19227 6670 19227 4 uio_oe[1]
rlabel metal1 s 5888 21046 5888 21046 4 uio_oe[2]
rlabel metal2 s 5014 21335 5014 21335 4 uio_oe[3]
rlabel metal3 s 4002 21131 4002 21131 4 uio_oe[4]
rlabel metal2 s 1610 20553 1610 20553 4 uio_oe[5]
rlabel metal1 s 2438 21080 2438 21080 4 uio_oe[6]
rlabel metal2 s 1334 21403 1334 21403 4 uio_oe[7]
rlabel metal4 s 11868 21389 11868 21389 4 uio_out[0]
rlabel metal4 s 11132 20709 11132 20709 4 uio_out[1]
rlabel metal4 s 10396 21593 10396 21593 4 uio_out[2]
rlabel metal4 s 9630 22104 9690 22304 4 uio_out[3]
port 33 nsew
rlabel metal2 s 12558 21811 12558 21811 4 uio_out[4]
rlabel metal4 s 8158 22104 8218 22304 4 uio_out[5]
port 35 nsew
rlabel metal4 s 7452 22001 7452 22001 4 uio_out[6]
rlabel metal4 s 6716 22001 6716 22001 4 uio_out[7]
rlabel metal1 s 14168 21046 14168 21046 4 uo_out[0]
rlabel metal2 s 13754 20689 13754 20689 4 uo_out[1]
rlabel metal2 s 13762 21114 13762 21114 4 uo_out[2]
rlabel metal1 s 14858 21386 14858 21386 4 uo_out[3]
rlabel metal1 s 13616 21590 13616 21590 4 uo_out[4]
rlabel metal2 s 13432 18156 13432 18156 4 uo_out[5]
rlabel metal1 s 13110 21318 13110 21318 4 uo_out[6]
rlabel metal1 s 14352 21590 14352 21590 4 uo_out[7]
flabel metal4 s 31488 496 31808 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23714 496 24034 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 15940 496 16260 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8166 496 8486 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 27601 496 27921 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 19827 496 20147 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12053 496 12373 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4279 496 4599 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 30974 22104 31034 22304 0 FreeSans 600 90 0 0 clk
port 3 nsew
flabel metal4 s 31710 22104 31770 22304 0 FreeSans 600 90 0 0 ena
port 4 nsew
flabel metal4 s 30238 22104 30298 22304 0 FreeSans 600 90 0 0 rst_n
port 5 nsew
flabel metal4 s 29502 22104 29562 22304 0 FreeSans 600 90 0 0 ui_in[0]
port 6 nsew
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 600 90 0 0 ui_in[1]
port 7 nsew
flabel metal4 s 28030 22104 28090 22304 0 FreeSans 600 90 0 0 ui_in[2]
port 8 nsew
flabel metal4 s 27294 22104 27354 22304 0 FreeSans 600 90 0 0 ui_in[3]
port 9 nsew
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 600 90 0 0 ui_in[4]
port 10 nsew
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 600 90 0 0 ui_in[5]
port 11 nsew
flabel metal4 s 25086 22104 25146 22304 0 FreeSans 600 90 0 0 ui_in[6]
port 12 nsew
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 600 90 0 0 ui_in[7]
port 13 nsew
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 600 90 0 0 uio_in[0]
port 14 nsew
flabel metal4 s 22878 22104 22938 22304 0 FreeSans 600 90 0 0 uio_in[1]
port 15 nsew
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 600 90 0 0 uio_in[2]
port 16 nsew
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 600 90 0 0 uio_in[3]
port 17 nsew
flabel metal4 s 20670 22104 20730 22304 0 FreeSans 600 90 0 0 uio_in[4]
port 18 nsew
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 600 90 0 0 uio_in[5]
port 19 nsew
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 600 90 0 0 uio_in[6]
port 20 nsew
flabel metal4 s 18462 22104 18522 22304 0 FreeSans 600 90 0 0 uio_in[7]
port 21 nsew
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 600 90 0 0 uio_oe[0]
port 22 nsew
flabel metal4 s 5214 22104 5274 22304 0 FreeSans 600 90 0 0 uio_oe[1]
port 23 nsew
flabel metal4 s 4478 22104 4538 22304 0 FreeSans 600 90 0 0 uio_oe[2]
port 24 nsew
flabel metal4 s 3742 22104 3802 22304 0 FreeSans 600 90 0 0 uio_oe[3]
port 25 nsew
flabel metal4 s 3006 22104 3066 22304 0 FreeSans 600 90 0 0 uio_oe[4]
port 26 nsew
flabel metal4 s 2270 22104 2330 22304 0 FreeSans 600 90 0 0 uio_oe[5]
port 27 nsew
flabel metal4 s 1534 22104 1594 22304 0 FreeSans 600 90 0 0 uio_oe[6]
port 28 nsew
flabel metal4 s 798 22104 858 22304 0 FreeSans 600 90 0 0 uio_oe[7]
port 29 nsew
flabel metal4 s 11838 22104 11898 22304 0 FreeSans 600 90 0 0 uio_out[0]
port 30 nsew
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 600 90 0 0 uio_out[1]
port 31 nsew
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 600 90 0 0 uio_out[2]
port 32 nsew
flabel metal4 s 9660 22204 9660 22204 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 600 90 0 0 uio_out[4]
port 34 nsew
flabel metal4 s 8188 22204 8188 22204 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 7422 22104 7482 22304 0 FreeSans 600 90 0 0 uio_out[6]
port 36 nsew
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 600 90 0 0 uio_out[7]
port 37 nsew
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 600 90 0 0 uo_out[0]
port 38 nsew
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 600 90 0 0 uo_out[1]
port 39 nsew
flabel metal4 s 16254 22104 16314 22304 0 FreeSans 600 90 0 0 uo_out[2]
port 40 nsew
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 600 90 0 0 uo_out[3]
port 41 nsew
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 600 90 0 0 uo_out[4]
port 42 nsew
flabel metal4 s 14046 22104 14106 22304 0 FreeSans 600 90 0 0 uo_out[5]
port 43 nsew
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 600 90 0 0 uo_out[6]
port 44 nsew
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 600 90 0 0 uo_out[7]
port 45 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 22304
string GDS_END 4029328
string GDS_FILE tt_um_dvxf_dj8v.gds
string GDS_START 848424
<< end >>
