magic
tech sky130A
magscale 1 2
timestamp 1717170941
<< metal1 >>
rect 704 21700 904 22564
rect 704 21640 796 21700
rect 856 21640 904 21700
rect 704 19902 904 21640
rect 704 19696 904 19702
rect 1264 21578 1464 22244
rect 1264 21518 1336 21578
rect 1396 21518 1464 21578
rect 1264 19502 1464 21518
rect 2206 22206 2406 22584
rect 2206 22146 2268 22206
rect 2328 22146 2406 22206
rect 1258 19302 1264 19502
rect 1464 19302 1470 19502
rect 2206 19140 2406 22146
rect 2206 18934 2406 18940
rect 3164 22164 3364 22546
rect 3164 22104 3226 22164
rect 3286 22104 3364 22164
rect 3164 18718 3364 22104
rect 3164 18512 3364 18518
rect 3644 22130 3844 22586
rect 3644 22070 3740 22130
rect 3800 22070 3844 22130
rect 3644 18278 3844 22070
rect 4666 22144 4866 22466
rect 4666 22084 4748 22144
rect 4808 22084 4866 22144
rect 4226 18278 4426 18284
rect 3644 18078 4226 18278
rect 4226 18072 4426 18078
rect 4666 17898 4866 22084
rect 4666 17692 4866 17698
rect 5128 22156 5328 22486
rect 5128 22096 5212 22156
rect 5272 22096 5328 22156
rect 5128 17516 5328 22096
rect 5888 22144 6088 22486
rect 5888 22084 5948 22144
rect 6008 22084 6088 22144
rect 5368 17516 5568 17522
rect 5128 17316 5368 17516
rect 5368 17310 5568 17316
rect 5888 17152 6088 22084
rect 26174 19902 26374 19922
rect 6284 19702 6290 19902
rect 6490 19702 26374 19902
rect 6264 19302 6270 19502
rect 6470 19302 25806 19502
rect 6284 18940 6290 19140
rect 6490 18940 25186 19140
rect 6290 18718 6490 18724
rect 6490 18518 24608 18718
rect 6290 18512 6490 18518
rect 6270 18278 6470 18284
rect 6470 18078 23974 18278
rect 6270 18072 6470 18078
rect 6284 17698 6290 17898
rect 6490 17698 23374 17898
rect 6344 17316 6350 17516
rect 6550 17316 22774 17516
rect 5888 16952 22174 17152
rect 22574 16952 22774 17316
rect 23174 16952 23374 17698
rect 23774 16952 23974 18078
rect 24408 16952 24608 18518
rect 24986 16952 25186 18940
rect 25606 16952 25806 19302
rect 26174 16952 26374 19702
rect 20594 15540 20600 15740
rect 20800 15540 20806 15740
rect 20600 2150 20800 15540
rect 27174 7552 27700 7752
rect 27580 7260 27700 7552
rect 27580 7134 27700 7140
<< via1 >>
rect 796 21640 856 21700
rect 704 19702 904 19902
rect 1336 21518 1396 21578
rect 2268 22146 2328 22206
rect 1264 19302 1464 19502
rect 2206 18940 2406 19140
rect 3226 22104 3286 22164
rect 3164 18518 3364 18718
rect 3740 22070 3800 22130
rect 4748 22084 4808 22144
rect 4226 18078 4426 18278
rect 4666 17698 4866 17898
rect 5212 22096 5272 22156
rect 5948 22084 6008 22144
rect 5368 17316 5568 17516
rect 6290 19702 6490 19902
rect 6270 19302 6470 19502
rect 6290 18940 6490 19140
rect 6290 18518 6490 18718
rect 6270 18078 6470 18278
rect 6290 17698 6490 17898
rect 6350 17316 6550 17516
rect 20600 15540 20800 15740
rect 27580 7140 27700 7260
<< metal2 >>
rect 2268 22318 2328 22320
rect 2261 22262 2270 22318
rect 2326 22262 2335 22318
rect 2268 22206 2328 22262
rect 3226 22254 3286 22256
rect 3219 22198 3228 22254
rect 3284 22198 3293 22254
rect 5948 22200 6008 22202
rect 2268 22140 2328 22146
rect 3226 22164 3286 22198
rect 3740 22196 3800 22198
rect 5212 22196 5272 22198
rect 3733 22140 3742 22196
rect 3798 22140 3807 22196
rect 4748 22190 4808 22192
rect 4741 22144 4750 22190
rect 4806 22144 4815 22190
rect 3226 22098 3286 22104
rect 3740 22130 3800 22140
rect 4741 22134 4748 22144
rect 4808 22134 4815 22144
rect 5205 22156 5214 22196
rect 5270 22156 5279 22196
rect 5205 22140 5212 22156
rect 5272 22140 5279 22156
rect 5941 22144 5950 22200
rect 6006 22144 6015 22200
rect 5212 22090 5272 22096
rect 4748 22078 4808 22084
rect 5948 22078 6008 22084
rect 3740 22064 3800 22070
rect 796 21820 856 21822
rect 789 21764 798 21820
rect 854 21764 863 21820
rect 796 21700 856 21764
rect 1336 21698 1396 21700
rect 1329 21642 1338 21698
rect 1394 21642 1403 21698
rect 796 21634 856 21640
rect 1336 21578 1396 21642
rect 1336 21512 1396 21518
rect 6290 19902 6490 19908
rect 698 19702 704 19902
rect 904 19702 6290 19902
rect 6290 19696 6490 19702
rect 1264 19502 1464 19508
rect 6270 19502 6470 19508
rect 1464 19302 6270 19502
rect 1264 19296 1464 19302
rect 6270 19296 6470 19302
rect 6290 19140 6490 19146
rect 2200 18940 2206 19140
rect 2406 18940 6290 19140
rect 6290 18934 6490 18940
rect 3158 18518 3164 18718
rect 3364 18518 6290 18718
rect 6490 18518 6496 18718
rect 4220 18078 4226 18278
rect 4426 18078 6270 18278
rect 6470 18078 6476 18278
rect 6290 17898 6490 17904
rect 4660 17698 4666 17898
rect 4866 17698 6290 17898
rect 6290 17692 6490 17698
rect 6350 17516 6550 17522
rect 5362 17316 5368 17516
rect 5568 17316 6350 17516
rect 6350 17310 6550 17316
rect 20600 16395 20800 16400
rect 20596 16205 20605 16395
rect 20795 16205 20804 16395
rect 20600 15740 20800 16205
rect 20600 15534 20800 15540
rect 27574 7140 27580 7260
rect 27700 7140 27706 7260
rect 27580 5280 27700 7140
rect 29465 5280 29575 5284
rect 27580 5275 29580 5280
rect 27580 5165 29465 5275
rect 29575 5165 29580 5275
rect 27580 5160 29580 5165
rect 29465 5156 29575 5160
<< via2 >>
rect 2270 22262 2326 22318
rect 3228 22198 3284 22254
rect 3742 22140 3798 22196
rect 4750 22144 4806 22190
rect 4750 22134 4806 22144
rect 5214 22156 5270 22196
rect 5214 22140 5270 22156
rect 5950 22144 6006 22200
rect 798 21764 854 21820
rect 1338 21642 1394 21698
rect 20605 16205 20795 16395
rect 29465 5165 29575 5275
<< metal3 >>
rect 2260 22386 2266 22450
rect 2330 22386 2336 22450
rect 3224 22400 3288 22406
rect 2268 22323 2328 22386
rect 3224 22330 3288 22336
rect 2265 22318 2331 22323
rect 2265 22262 2270 22318
rect 2326 22262 2331 22318
rect 2265 22257 2331 22262
rect 3226 22259 3286 22330
rect 3732 22296 3738 22360
rect 3802 22296 3808 22360
rect 3223 22254 3289 22259
rect 3223 22198 3228 22254
rect 3284 22198 3289 22254
rect 3740 22201 3800 22296
rect 4740 22290 4746 22354
rect 4810 22290 4816 22354
rect 5204 22318 5210 22382
rect 5274 22318 5280 22382
rect 3223 22193 3289 22198
rect 3737 22196 3803 22201
rect 3737 22140 3742 22196
rect 3798 22140 3803 22196
rect 4748 22195 4808 22290
rect 5212 22201 5272 22318
rect 5940 22286 5946 22350
rect 6010 22286 6016 22350
rect 5948 22205 6008 22286
rect 5209 22196 5275 22201
rect 3737 22135 3803 22140
rect 4745 22190 4811 22195
rect 4745 22134 4750 22190
rect 4806 22134 4811 22190
rect 5209 22140 5214 22196
rect 5270 22140 5275 22196
rect 5209 22135 5275 22140
rect 5945 22200 6011 22205
rect 5945 22144 5950 22200
rect 6006 22144 6011 22200
rect 5945 22139 6011 22144
rect 4745 22129 4811 22134
rect 2413 22028 2711 22033
rect 8159 22028 8165 22043
rect 2412 22027 8165 22028
rect 788 21910 794 21974
rect 858 21910 864 21974
rect 796 21825 856 21910
rect 793 21820 859 21825
rect 793 21764 798 21820
rect 854 21764 859 21820
rect 1328 21800 1334 21864
rect 1398 21800 1404 21864
rect 793 21759 859 21764
rect 1336 21703 1396 21800
rect 2412 21729 2413 22027
rect 2711 21729 8165 22027
rect 2412 21728 8165 21729
rect 2413 21723 2711 21728
rect 8159 21725 8165 21728
rect 8483 22028 8489 22043
rect 15933 22028 15939 22043
rect 8483 21728 15939 22028
rect 8483 21725 8489 21728
rect 15933 21725 15939 21728
rect 16257 22028 16263 22043
rect 23707 22028 23713 22043
rect 16257 21955 23713 22028
rect 16257 21757 20601 21955
rect 20799 21757 23713 21955
rect 16257 21728 23713 21757
rect 16257 21725 16263 21728
rect 23707 21725 23713 21728
rect 24031 22028 24037 22043
rect 31481 22028 31487 22043
rect 24031 21728 31487 22028
rect 24031 21725 24037 21728
rect 31481 21725 31487 21728
rect 31805 22028 31811 22043
rect 31805 21728 31812 22028
rect 31805 21725 31811 21728
rect 1333 21698 1399 21703
rect 1333 21642 1338 21698
rect 1394 21642 1399 21698
rect 1333 21637 1399 21642
rect 733 21366 1031 21371
rect 4274 21366 4280 21377
rect 732 21365 4280 21366
rect 732 21067 733 21365
rect 1031 21067 4280 21365
rect 732 21066 4280 21067
rect 733 21061 1031 21066
rect 4274 21063 4280 21066
rect 4594 21366 4600 21377
rect 12046 21366 12052 21377
rect 4594 21066 12052 21366
rect 4594 21063 4600 21066
rect 12046 21059 12052 21066
rect 12370 21366 12376 21377
rect 19820 21366 19826 21381
rect 12370 21066 19826 21366
rect 12370 21059 12376 21066
rect 19820 21063 19826 21066
rect 20144 21366 20150 21381
rect 27594 21366 27600 21379
rect 20144 21066 27600 21366
rect 20144 21063 20150 21066
rect 27594 21061 27600 21066
rect 27918 21366 27924 21379
rect 27918 21066 27926 21366
rect 27918 21061 27924 21066
rect 20600 20714 20800 20720
rect 20600 16395 20800 20514
rect 20600 16205 20605 16395
rect 20795 16205 20800 16395
rect 20600 16200 20800 16205
rect 31313 5280 31431 5285
rect 29460 5279 31432 5280
rect 29460 5275 31313 5279
rect 29460 5165 29465 5275
rect 29575 5165 31313 5275
rect 29460 5161 31313 5165
rect 31431 5161 31432 5279
rect 29460 5160 31432 5161
rect 31313 5155 31431 5160
<< via3 >>
rect 2266 22386 2330 22450
rect 3224 22336 3288 22400
rect 3738 22296 3802 22360
rect 4746 22290 4810 22354
rect 5210 22318 5274 22382
rect 5946 22286 6010 22350
rect 794 21910 858 21974
rect 1334 21800 1398 21864
rect 2413 21729 2711 22027
rect 8165 21725 8483 22043
rect 15939 21725 16257 22043
rect 20601 21757 20799 21955
rect 23713 21725 24031 22043
rect 31487 21725 31805 22043
rect 733 21067 1031 21365
rect 4280 21063 4594 21377
rect 12052 21059 12370 21377
rect 19826 21063 20144 21381
rect 27600 21061 27918 21379
rect 20600 20514 20800 20714
rect 31313 5161 31431 5279
<< metal4 >>
rect 798 45070 858 45152
rect 790 44952 858 45070
rect 790 44822 850 44952
rect 1534 44822 1594 45152
rect 2270 44822 2330 45152
rect 3006 44822 3066 45152
rect 3742 44822 3802 45152
rect 4478 44822 4538 45152
rect 5214 44822 5274 45152
rect 5950 44822 6010 45152
rect 6686 44836 6746 45152
rect 790 44820 6010 44822
rect 594 44762 6010 44820
rect 594 44760 850 44762
rect 594 44162 654 44760
rect 790 44758 850 44760
rect 1534 44758 1594 44762
rect 2270 44758 2330 44762
rect 3006 44758 3066 44762
rect 3742 44758 3802 44762
rect 4478 44758 4538 44762
rect 5214 44758 5274 44762
rect 5950 44758 6010 44762
rect 6684 44758 6746 44836
rect 7422 44820 7482 45152
rect 8158 44824 8218 45152
rect 7420 44758 7482 44820
rect 8156 44758 8218 44824
rect 8894 44816 8954 45152
rect 9630 44836 9690 45152
rect 10366 44840 10426 45152
rect 11102 44840 11162 45152
rect 8892 44758 8954 44816
rect 9628 44758 9690 44836
rect 10364 44758 10426 44840
rect 11100 44758 11162 44840
rect 11838 44828 11898 45152
rect 12574 44834 12634 45152
rect 13310 44836 13370 45152
rect 11836 44758 11898 44828
rect 12572 44758 12634 44834
rect 13308 44758 13370 44836
rect 14046 44818 14106 45152
rect 14782 44838 14842 45152
rect 15518 44860 15578 45152
rect 14044 44758 14106 44818
rect 14780 44758 14842 44838
rect 15516 44758 15578 44860
rect 16254 44842 16314 45152
rect 16252 44758 16314 44842
rect 16990 44836 17050 45152
rect 17726 45052 17786 45152
rect 16988 44758 17050 44836
rect 17724 44952 17786 45052
rect 18462 45040 18522 45152
rect 19198 45066 19258 45152
rect 19934 45074 19994 45152
rect 18460 44952 18522 45040
rect 19196 44952 19258 45066
rect 19932 44952 19994 45074
rect 20670 45064 20730 45152
rect 21406 45090 21466 45152
rect 20668 44952 20730 45064
rect 21404 44952 21466 45090
rect 22142 45076 22202 45152
rect 22140 44952 22202 45076
rect 22878 45008 22938 45152
rect 432 44152 654 44162
rect 200 44102 654 44152
rect 200 21366 500 44102
rect 796 21975 856 44570
rect 1532 21994 1592 44570
rect 793 21974 859 21975
rect 793 21910 794 21974
rect 858 21910 859 21974
rect 793 21909 859 21910
rect 1336 21934 1592 21994
rect 1688 22028 1988 44370
rect 2268 22451 2328 44530
rect 2265 22450 2331 22451
rect 2265 22386 2266 22450
rect 2330 22386 2331 22450
rect 2265 22385 2331 22386
rect 3004 22398 3064 44498
rect 3223 22400 3289 22401
rect 3223 22398 3224 22400
rect 3004 22338 3224 22398
rect 3223 22336 3224 22338
rect 3288 22336 3289 22400
rect 3740 22361 3800 44488
rect 4476 44444 4808 44504
rect 3223 22335 3289 22336
rect 3737 22360 3803 22361
rect 3737 22296 3738 22360
rect 3802 22296 3803 22360
rect 3737 22295 3803 22296
rect 1688 22027 2712 22028
rect 1336 21865 1396 21934
rect 1333 21864 1399 21865
rect 1333 21800 1334 21864
rect 1398 21800 1399 21864
rect 1333 21799 1399 21800
rect 1688 21729 2413 22027
rect 2711 21729 2712 22027
rect 1688 21728 2712 21729
rect 200 21365 1032 21366
rect 200 21067 733 21365
rect 1031 21067 1032 21365
rect 200 21066 1032 21067
rect 200 1000 500 21066
rect 1688 1104 1988 21728
rect 4279 21377 4595 23712
rect 4748 22355 4808 44444
rect 5212 22383 5272 44524
rect 5209 22382 5275 22383
rect 4745 22354 4811 22355
rect 4745 22290 4746 22354
rect 4810 22290 4811 22354
rect 5209 22318 5210 22382
rect 5274 22318 5275 22382
rect 5948 22351 6008 44488
rect 6684 44326 6744 44758
rect 7420 44320 7480 44758
rect 8156 44444 8216 44758
rect 8892 44470 8952 44758
rect 9628 44490 9688 44758
rect 10364 44498 10424 44758
rect 11100 44510 11160 44758
rect 11836 44518 11896 44758
rect 12572 44478 12632 44758
rect 13308 44490 13368 44758
rect 14044 44484 14104 44758
rect 14780 44494 14840 44758
rect 15516 44500 15576 44758
rect 16252 44502 16312 44758
rect 16988 44484 17048 44758
rect 17724 44478 17784 44952
rect 18460 44490 18520 44952
rect 19196 44486 19256 44952
rect 19932 44482 19992 44952
rect 20668 44492 20728 44952
rect 21404 44466 21464 44952
rect 22140 44454 22200 44952
rect 22876 44758 22938 45008
rect 23614 44864 23674 45152
rect 24350 45117 24410 45152
rect 23612 44758 23674 44864
rect 24347 44952 24410 45117
rect 24347 44860 24407 44952
rect 24347 44758 24408 44860
rect 25086 44854 25146 45152
rect 25822 44854 25882 45152
rect 26558 45117 26618 45152
rect 22876 44452 22936 44758
rect 23612 44492 23672 44758
rect 24348 44470 24408 44758
rect 25084 44758 25146 44854
rect 25820 44758 25882 44854
rect 26554 44952 26618 45117
rect 26554 44836 26614 44952
rect 27294 44880 27354 45152
rect 28030 45117 28090 45152
rect 26554 44758 26616 44836
rect 25084 44466 25144 44758
rect 25820 44444 25880 44758
rect 26556 44436 26616 44758
rect 27292 44758 27354 44880
rect 28026 44952 28090 45117
rect 28026 44866 28086 44952
rect 28026 44758 28088 44866
rect 28766 44848 28826 45152
rect 29502 45125 29562 45152
rect 27292 44440 27352 44758
rect 28028 44432 28088 44758
rect 28764 44758 28826 44848
rect 29494 44952 29562 45125
rect 29494 44862 29554 44952
rect 30238 44862 30298 45152
rect 30974 45074 31034 45152
rect 30974 44952 31035 45074
rect 31710 45060 31770 45152
rect 30975 44872 31035 44952
rect 29494 44758 29560 44862
rect 28764 44434 28824 44758
rect 29500 44458 29560 44758
rect 30236 44758 30298 44862
rect 30972 44758 31035 44872
rect 31708 44952 31770 45060
rect 30236 44420 30296 44758
rect 30972 44460 31032 44758
rect 31708 44480 31768 44952
rect 5209 22317 5275 22318
rect 5945 22350 6011 22351
rect 5212 22302 5272 22317
rect 4745 22289 4811 22290
rect 5945 22286 5946 22350
rect 6010 22286 6011 22350
rect 5945 22285 6011 22286
rect 8164 22043 8484 23204
rect 8164 21725 8165 22043
rect 8483 21725 8484 22043
rect 8164 21724 8484 21725
rect 4279 21063 4280 21377
rect 4594 21063 4595 21377
rect 4279 21062 4595 21063
rect 12051 21377 12371 23714
rect 15938 22043 16258 23188
rect 15938 21725 15939 22043
rect 16257 21725 16258 22043
rect 15938 21724 16258 21725
rect 12051 21059 12052 21377
rect 12370 21059 12371 21377
rect 19825 21381 20145 23714
rect 23712 22043 24032 23184
rect 19825 21063 19826 21381
rect 20144 21063 20145 21381
rect 19825 21062 20145 21063
rect 20600 21955 20800 21956
rect 20600 21757 20601 21955
rect 20799 21757 20800 21955
rect 12051 21058 12371 21059
rect 20600 20715 20800 21757
rect 23712 21725 23713 22043
rect 24031 21725 24032 22043
rect 23712 21724 24032 21725
rect 27599 21379 27919 23714
rect 31486 22043 31806 23170
rect 31486 21725 31487 22043
rect 31805 21725 31806 22043
rect 31486 21724 31806 21725
rect 27599 21061 27600 21379
rect 27918 21061 27919 21379
rect 27599 21060 27919 21061
rect 20599 20714 20801 20715
rect 20599 20514 20600 20714
rect 20800 20514 20801 20714
rect 20599 20513 20801 20514
rect 31312 5279 31432 5280
rect 31312 5161 31313 5279
rect 31431 5161 31432 5279
rect 31312 354 31432 5161
rect 370 0 550 354
rect 4786 0 4966 354
rect 9202 0 9382 354
rect 13618 0 13798 354
rect 18034 0 18214 354
rect 22450 0 22630 354
rect 26866 0 27046 354
rect 31252 0 31492 354
use r2r  r2r_0
timestamp 1710085389
transform 1 0 23174 0 1 -448
box -2600 2400 4200 17600
use tt_um_dvxf_dj8v  tt_um_dvxf_dj8v_0
timestamp 1717153468
transform 1 0 -2 0 1 22274
box 492 496 31808 22304
<< labels >>
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1688 1104 1988 44256 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
