MACRO tt_um_dvxf_dj8v_dac
  CLASS BLOCK ;
  FOREIGN tt_um_dvxf_dj8v_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 662.271484 ;
    ANTENNADIFFAREA 1022.153198 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 8.440 5.520 9.940 221.280 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 2.560 218.755 158.420 220.360 ;
      LAYER pwell ;
        RECT 2.755 217.555 4.125 218.365 ;
        RECT 4.685 218.355 7.285 218.465 ;
        RECT 4.685 218.235 8.700 218.355 ;
        RECT 13.345 218.235 14.265 218.455 ;
        RECT 4.685 217.555 15.625 218.235 ;
        RECT 15.645 217.640 16.075 218.425 ;
        RECT 16.095 218.235 17.440 218.465 ;
        RECT 22.445 218.235 23.375 218.455 ;
        RECT 26.095 218.235 28.305 218.465 ;
        RECT 16.095 217.555 17.925 218.235 ;
        RECT 17.935 217.555 28.305 218.235 ;
        RECT 28.525 217.640 28.955 218.425 ;
        RECT 28.975 218.235 29.905 218.465 ;
        RECT 28.975 217.555 32.875 218.235 ;
        RECT 33.115 217.555 34.485 218.335 ;
        RECT 40.455 218.235 41.385 218.465 ;
        RECT 34.505 217.555 37.245 218.235 ;
        RECT 37.485 217.555 41.385 218.235 ;
        RECT 41.405 217.640 41.835 218.425 ;
        RECT 41.855 217.555 44.595 218.235 ;
        RECT 44.615 217.555 45.985 218.335 ;
        RECT 49.195 218.235 50.125 218.465 ;
        RECT 46.225 217.555 50.125 218.235 ;
        RECT 50.135 217.555 52.875 218.235 ;
        RECT 52.895 217.555 54.265 218.365 ;
        RECT 54.285 217.640 54.715 218.425 ;
        RECT 64.705 218.235 65.635 218.465 ;
        RECT 55.205 217.555 57.945 218.235 ;
        RECT 58.875 217.555 61.615 218.235 ;
        RECT 61.635 217.555 64.375 218.235 ;
        RECT 64.705 217.555 66.540 218.235 ;
        RECT 67.165 217.640 67.595 218.425 ;
        RECT 69.690 218.235 70.825 218.465 ;
        RECT 67.615 217.555 70.825 218.235 ;
        RECT 70.835 218.235 71.755 218.465 ;
        RECT 73.620 218.235 74.965 218.465 ;
        RECT 70.835 217.555 73.125 218.235 ;
        RECT 73.135 217.555 74.965 218.235 ;
        RECT 74.975 217.555 78.645 218.365 ;
        RECT 78.655 217.555 80.025 218.365 ;
        RECT 80.045 217.640 80.475 218.425 ;
        RECT 80.495 217.555 82.325 218.365 ;
        RECT 82.335 218.265 83.265 218.465 ;
        RECT 84.600 218.265 85.545 218.465 ;
        RECT 82.335 217.785 85.545 218.265 ;
        RECT 82.475 217.585 85.545 217.785 ;
        RECT 2.895 217.345 3.065 217.555 ;
        RECT 4.275 217.505 4.445 217.535 ;
        RECT 4.270 217.395 4.445 217.505 ;
        RECT 14.850 217.395 14.970 217.505 ;
        RECT 4.275 217.345 4.445 217.395 ;
        RECT 15.315 217.345 15.485 217.555 ;
        RECT 16.695 217.345 16.865 217.535 ;
        RECT 17.615 217.365 17.785 217.555 ;
        RECT 18.075 217.365 18.245 217.555 ;
        RECT 18.350 217.345 18.520 217.535 ;
        RECT 22.225 217.390 22.385 217.500 ;
        RECT 23.410 217.345 23.580 217.535 ;
        RECT 27.275 217.345 27.445 217.535 ;
        RECT 29.115 217.345 29.285 217.535 ;
        RECT 29.390 217.365 29.560 217.555 ;
        RECT 33.255 217.365 33.425 217.555 ;
        RECT 33.900 217.345 34.070 217.535 ;
        RECT 34.630 217.395 34.750 217.505 ;
        RECT 36.935 217.365 37.105 217.555 ;
        RECT 40.800 217.365 40.970 217.555 ;
        RECT 41.995 217.365 42.165 217.555 ;
        RECT 45.215 217.345 45.385 217.535 ;
        RECT 45.675 217.505 45.845 217.555 ;
        RECT 45.670 217.395 45.845 217.505 ;
        RECT 45.675 217.365 45.845 217.395 ;
        RECT 46.410 217.345 46.580 217.535 ;
        RECT 49.540 217.365 49.710 217.555 ;
        RECT 50.275 217.365 50.445 217.555 ;
        RECT 50.550 217.345 50.720 217.535 ;
        RECT 53.035 217.365 53.205 217.555 ;
        RECT 54.870 217.395 54.990 217.505 ;
        RECT 55.150 217.345 55.320 217.535 ;
        RECT 57.635 217.365 57.805 217.555 ;
        RECT 58.105 217.400 58.265 217.510 ;
        RECT 59.015 217.345 59.185 217.555 ;
        RECT 60.670 217.345 60.840 217.535 ;
        RECT 61.775 217.365 61.945 217.555 ;
        RECT 66.375 217.535 66.540 217.555 ;
        RECT 66.375 217.365 66.545 217.535 ;
        RECT 66.835 217.505 67.005 217.535 ;
        RECT 66.830 217.395 67.005 217.505 ;
        RECT 67.290 217.395 67.410 217.505 ;
        RECT 66.835 217.345 67.005 217.395 ;
        RECT 67.755 217.345 67.925 217.555 ;
        RECT 70.050 217.395 70.170 217.505 ;
        RECT 70.515 217.345 70.685 217.535 ;
        RECT 72.815 217.365 72.985 217.555 ;
        RECT 73.275 217.345 73.445 217.555 ;
        RECT 75.115 217.505 75.285 217.555 ;
        RECT 75.110 217.395 75.285 217.505 ;
        RECT 75.115 217.365 75.285 217.395 ;
        RECT 75.580 217.345 75.750 217.535 ;
        RECT 78.795 217.365 78.965 217.555 ;
        RECT 79.265 217.390 79.425 217.500 ;
        RECT 80.635 217.365 80.805 217.555 ;
        RECT 82.475 217.365 82.645 217.585 ;
        RECT 84.600 217.555 85.545 217.585 ;
        RECT 85.555 217.555 91.065 218.365 ;
        RECT 91.075 217.555 92.905 218.365 ;
        RECT 92.925 217.640 93.355 218.425 ;
        RECT 93.385 217.555 97.045 218.465 ;
        RECT 97.055 217.555 100.725 218.365 ;
        RECT 101.755 217.555 103.945 218.465 ;
        RECT 103.955 217.555 105.785 218.365 ;
        RECT 105.805 217.640 106.235 218.425 ;
        RECT 106.715 218.235 107.645 218.465 ;
        RECT 106.715 217.555 109.465 218.235 ;
        RECT 109.475 217.555 114.985 218.365 ;
        RECT 114.995 217.555 118.665 218.365 ;
        RECT 118.685 217.640 119.115 218.425 ;
        RECT 119.135 217.555 122.345 218.465 ;
        RECT 122.355 217.555 123.725 218.335 ;
        RECT 123.735 217.555 126.485 218.365 ;
        RECT 126.495 218.235 127.425 218.465 ;
        RECT 126.495 217.555 129.245 218.235 ;
        RECT 129.255 217.555 130.625 218.335 ;
        RECT 131.565 217.640 131.995 218.425 ;
        RECT 132.015 217.555 133.385 218.335 ;
        RECT 133.395 218.235 134.325 218.465 ;
        RECT 133.395 217.555 136.145 218.235 ;
        RECT 136.155 217.555 137.525 218.335 ;
        RECT 137.535 217.555 138.905 218.335 ;
        RECT 138.915 217.555 140.285 218.365 ;
        RECT 140.295 217.555 141.665 218.335 ;
        RECT 141.675 217.555 144.425 218.365 ;
        RECT 144.445 217.640 144.875 218.425 ;
        RECT 144.895 217.555 147.505 218.465 ;
        RECT 147.655 217.555 149.025 218.335 ;
        RECT 149.035 217.555 150.405 218.335 ;
        RECT 151.335 217.555 152.705 218.335 ;
        RECT 152.715 217.555 156.385 218.365 ;
        RECT 156.855 217.555 158.225 218.365 ;
        RECT 83.395 217.345 83.565 217.535 ;
        RECT 83.855 217.345 84.025 217.535 ;
        RECT 85.695 217.365 85.865 217.555 ;
        RECT 89.375 217.345 89.545 217.535 ;
        RECT 91.215 217.365 91.385 217.555 ;
        RECT 92.130 217.395 92.250 217.505 ;
        RECT 92.595 217.345 92.765 217.535 ;
        RECT 93.510 217.365 93.680 217.555 ;
        RECT 97.195 217.345 97.365 217.555 ;
        RECT 97.655 217.345 97.825 217.535 ;
        RECT 100.410 217.395 100.530 217.505 ;
        RECT 100.885 217.400 101.045 217.510 ;
        RECT 101.790 217.345 101.960 217.535 ;
        RECT 102.255 217.345 102.425 217.535 ;
        RECT 103.630 217.365 103.800 217.555 ;
        RECT 104.095 217.365 104.265 217.555 ;
        RECT 106.390 217.395 106.510 217.505 ;
        RECT 109.155 217.345 109.325 217.555 ;
        RECT 109.615 217.345 109.785 217.555 ;
        RECT 112.370 217.395 112.490 217.505 ;
        RECT 115.135 217.365 115.305 217.555 ;
        RECT 119.280 217.535 119.450 217.555 ;
        RECT 116.050 217.345 116.220 217.535 ;
        RECT 2.755 216.535 4.125 217.345 ;
        RECT 4.135 216.665 14.505 217.345 ;
        RECT 8.645 216.445 9.575 216.665 ;
        RECT 12.295 216.435 14.505 216.665 ;
        RECT 15.175 216.565 16.545 217.345 ;
        RECT 16.555 216.565 17.925 217.345 ;
        RECT 17.935 216.665 21.835 217.345 ;
        RECT 22.995 216.665 26.895 217.345 ;
        RECT 17.935 216.435 18.865 216.665 ;
        RECT 22.995 216.435 23.925 216.665 ;
        RECT 27.135 216.565 28.505 217.345 ;
        RECT 28.525 216.475 28.955 217.260 ;
        RECT 28.975 216.565 30.345 217.345 ;
        RECT 30.585 216.665 34.485 217.345 ;
        RECT 33.555 216.435 34.485 216.665 ;
        RECT 35.155 216.665 45.525 217.345 ;
        RECT 45.995 216.665 49.895 217.345 ;
        RECT 50.135 216.665 54.035 217.345 ;
        RECT 35.155 216.435 37.365 216.665 ;
        RECT 40.085 216.445 41.015 216.665 ;
        RECT 45.995 216.435 46.925 216.665 ;
        RECT 50.135 216.435 51.065 216.665 ;
        RECT 54.285 216.475 54.715 217.260 ;
        RECT 54.735 216.665 58.635 217.345 ;
        RECT 54.735 216.435 55.665 216.665 ;
        RECT 58.875 216.535 60.245 217.345 ;
        RECT 60.255 216.665 64.155 217.345 ;
        RECT 64.405 216.665 67.145 217.345 ;
        RECT 67.615 216.665 69.905 217.345 ;
        RECT 70.375 216.665 73.115 217.345 ;
        RECT 60.255 216.435 61.185 216.665 ;
        RECT 68.985 216.435 69.905 216.665 ;
        RECT 73.135 216.535 74.965 217.345 ;
        RECT 75.435 216.435 79.090 217.345 ;
        RECT 80.045 216.475 80.475 217.260 ;
        RECT 80.495 216.665 83.705 217.345 ;
        RECT 80.495 216.435 81.630 216.665 ;
        RECT 83.715 216.535 89.225 217.345 ;
        RECT 89.235 216.535 91.985 217.345 ;
        RECT 92.455 216.435 95.205 217.345 ;
        RECT 95.215 216.665 97.505 217.345 ;
        RECT 95.215 216.435 96.135 216.665 ;
        RECT 97.515 216.535 100.265 217.345 ;
        RECT 100.755 216.435 102.105 217.345 ;
        RECT 102.115 216.535 105.785 217.345 ;
        RECT 105.805 216.475 106.235 217.260 ;
        RECT 106.255 216.665 109.465 217.345 ;
        RECT 106.255 216.435 107.390 216.665 ;
        RECT 109.475 216.535 112.225 217.345 ;
        RECT 112.890 216.435 116.365 217.345 ;
        RECT 116.520 217.315 116.690 217.535 ;
        RECT 119.275 217.365 119.450 217.535 ;
        RECT 121.110 217.395 121.230 217.505 ;
        RECT 119.275 217.345 119.445 217.365 ;
        RECT 121.580 217.345 121.750 217.535 ;
        RECT 123.415 217.365 123.585 217.555 ;
        RECT 123.875 217.365 124.045 217.555 ;
        RECT 124.795 217.345 124.965 217.535 ;
        RECT 127.555 217.345 127.725 217.535 ;
        RECT 128.935 217.365 129.105 217.555 ;
        RECT 129.395 217.345 129.565 217.535 ;
        RECT 130.315 217.365 130.485 217.555 ;
        RECT 130.785 217.400 130.945 217.510 ;
        RECT 131.230 217.395 131.350 217.505 ;
        RECT 132.150 217.395 132.270 217.505 ;
        RECT 132.610 217.345 132.780 217.535 ;
        RECT 133.075 217.365 133.245 217.555 ;
        RECT 133.995 217.345 134.165 217.535 ;
        RECT 135.835 217.365 136.005 217.555 ;
        RECT 137.215 217.365 137.385 217.555 ;
        RECT 138.595 217.365 138.765 217.555 ;
        RECT 139.055 217.365 139.225 217.555 ;
        RECT 139.970 217.345 140.140 217.535 ;
        RECT 140.435 217.365 140.605 217.555 ;
        RECT 141.815 217.365 141.985 217.555 ;
        RECT 118.180 217.315 119.125 217.345 ;
        RECT 116.375 216.635 119.125 217.315 ;
        RECT 118.180 216.435 119.125 216.635 ;
        RECT 119.135 216.535 120.965 217.345 ;
        RECT 121.435 216.435 124.355 217.345 ;
        RECT 124.665 216.435 127.395 217.345 ;
        RECT 127.430 216.435 129.245 217.345 ;
        RECT 129.255 216.535 131.085 217.345 ;
        RECT 131.565 216.475 131.995 217.260 ;
        RECT 132.495 216.435 133.845 217.345 ;
        RECT 133.855 216.535 136.605 217.345 ;
        RECT 136.630 216.435 140.285 217.345 ;
        RECT 140.295 217.315 141.250 217.345 ;
        RECT 142.280 217.315 142.450 217.535 ;
        RECT 142.735 217.345 142.905 217.535 ;
        RECT 145.040 217.365 145.210 217.555 ;
        RECT 148.255 217.345 148.425 217.535 ;
        RECT 148.715 217.365 148.885 217.555 ;
        RECT 150.095 217.505 150.265 217.555 ;
        RECT 150.090 217.395 150.265 217.505 ;
        RECT 150.095 217.365 150.265 217.395 ;
        RECT 150.555 217.345 150.725 217.535 ;
        RECT 152.395 217.365 152.565 217.555 ;
        RECT 152.855 217.365 153.025 217.555 ;
        RECT 153.315 217.345 153.485 217.535 ;
        RECT 156.085 217.390 156.245 217.500 ;
        RECT 156.530 217.395 156.650 217.505 ;
        RECT 157.915 217.345 158.085 217.555 ;
        RECT 140.295 216.635 142.575 217.315 ;
        RECT 140.295 216.435 141.250 216.635 ;
        RECT 142.595 216.535 148.105 217.345 ;
        RECT 148.115 216.535 149.945 217.345 ;
        RECT 150.415 216.435 153.165 217.345 ;
        RECT 153.175 216.665 155.915 217.345 ;
        RECT 156.855 216.535 158.225 217.345 ;
      LAYER nwell ;
        RECT 2.560 213.315 158.420 216.145 ;
      LAYER pwell ;
        RECT 2.755 212.115 4.125 212.925 ;
        RECT 4.595 212.115 5.965 212.895 ;
        RECT 5.975 212.795 6.905 213.025 ;
        RECT 10.115 212.795 11.045 213.025 ;
        RECT 5.975 212.115 9.875 212.795 ;
        RECT 10.115 212.115 14.015 212.795 ;
        RECT 14.255 212.115 15.625 212.895 ;
        RECT 15.645 212.200 16.075 212.985 ;
        RECT 20.605 212.795 21.535 213.015 ;
        RECT 24.255 212.795 26.465 213.025 ;
        RECT 16.095 212.115 26.465 212.795 ;
        RECT 27.795 212.795 30.005 213.025 ;
        RECT 32.725 212.795 33.655 213.015 ;
        RECT 27.795 212.115 38.165 212.795 ;
        RECT 38.645 212.115 41.385 212.795 ;
        RECT 41.405 212.200 41.835 212.985 ;
        RECT 44.615 212.795 45.545 213.025 ;
        RECT 51.955 212.795 52.885 213.025 ;
        RECT 56.945 212.915 57.865 213.025 ;
        RECT 56.945 212.795 59.280 212.915 ;
        RECT 63.945 212.795 64.865 213.015 ;
        RECT 41.865 212.115 44.605 212.795 ;
        RECT 44.615 212.115 48.515 212.795 ;
        RECT 48.985 212.115 52.885 212.795 ;
        RECT 53.825 212.115 56.565 212.795 ;
        RECT 56.945 212.115 66.225 212.795 ;
        RECT 67.165 212.200 67.595 212.985 ;
        RECT 67.625 212.115 68.975 213.025 ;
        RECT 68.995 212.115 70.365 212.925 ;
        RECT 70.375 212.115 74.045 213.025 ;
        RECT 74.055 212.115 75.405 213.025 ;
        RECT 75.435 212.115 77.265 212.925 ;
        RECT 77.275 212.115 78.625 213.025 ;
        RECT 80.730 212.795 81.865 213.025 ;
        RECT 78.655 212.115 81.865 212.795 ;
        RECT 81.895 212.115 83.245 213.025 ;
        RECT 83.715 212.115 85.065 213.025 ;
        RECT 85.095 212.115 88.015 213.025 ;
        RECT 88.315 212.795 89.235 213.025 ;
        RECT 88.315 212.115 90.605 212.795 ;
        RECT 90.615 212.115 92.445 212.925 ;
        RECT 92.925 212.200 93.355 212.985 ;
        RECT 93.375 212.115 98.885 212.925 ;
        RECT 99.895 212.115 102.895 213.025 ;
        RECT 103.035 212.115 104.405 212.925 ;
        RECT 104.415 212.115 107.890 213.025 ;
        RECT 108.095 212.115 110.845 212.925 ;
        RECT 110.855 212.115 113.260 213.025 ;
        RECT 113.615 212.115 117.285 212.925 ;
        RECT 117.295 212.115 118.665 212.925 ;
        RECT 118.685 212.200 119.115 212.985 ;
        RECT 119.135 212.115 122.805 212.925 ;
        RECT 122.815 212.115 124.645 213.025 ;
        RECT 124.655 212.115 130.165 212.925 ;
        RECT 130.175 212.115 133.845 212.925 ;
        RECT 134.315 212.795 135.685 213.025 ;
        RECT 134.315 212.115 138.445 212.795 ;
        RECT 138.455 212.115 143.965 212.925 ;
        RECT 144.445 212.200 144.875 212.985 ;
        RECT 144.895 212.115 147.680 213.025 ;
        RECT 148.115 212.115 150.855 212.795 ;
        RECT 150.875 212.115 152.245 212.925 ;
        RECT 152.335 212.115 154.545 213.025 ;
        RECT 155.015 212.115 156.365 213.025 ;
        RECT 156.855 212.115 158.225 212.925 ;
        RECT 2.895 211.905 3.065 212.115 ;
        RECT 4.270 211.955 4.390 212.065 ;
        RECT 4.735 211.905 4.905 212.115 ;
        RECT 6.390 211.925 6.560 212.115 ;
        RECT 10.530 211.925 10.700 212.115 ;
        RECT 15.315 211.905 15.485 212.115 ;
        RECT 16.235 211.925 16.405 212.115 ;
        RECT 18.075 211.905 18.245 212.095 ;
        RECT 26.825 211.960 26.985 212.070 ;
        RECT 27.745 211.950 27.905 212.060 ;
        RECT 29.110 211.955 29.230 212.065 ;
        RECT 29.575 211.905 29.745 212.095 ;
        RECT 37.855 211.925 38.025 212.115 ;
        RECT 38.310 211.955 38.430 212.065 ;
        RECT 40.155 211.905 40.325 212.095 ;
        RECT 41.075 211.925 41.245 212.115 ;
        RECT 44.295 211.925 44.465 212.115 ;
        RECT 45.030 211.925 45.200 212.115 ;
        RECT 49.350 211.955 49.470 212.065 ;
        RECT 51.195 211.905 51.365 212.095 ;
        RECT 52.300 211.925 52.470 212.115 ;
        RECT 53.045 211.960 53.205 212.070 ;
        RECT 53.955 211.905 54.125 212.095 ;
        RECT 55.150 211.905 55.320 212.095 ;
        RECT 56.255 211.925 56.425 212.115 ;
        RECT 59.010 211.955 59.130 212.065 ;
        RECT 61.775 211.905 61.945 212.095 ;
        RECT 62.235 211.905 62.405 212.095 ;
        RECT 63.615 211.905 63.785 212.095 ;
        RECT 65.915 211.925 66.085 212.115 ;
        RECT 66.385 211.960 66.545 212.070 ;
        RECT 67.755 211.925 67.925 212.115 ;
        RECT 69.135 211.905 69.305 212.115 ;
        RECT 70.520 211.925 70.690 212.115 ;
        RECT 74.655 211.905 74.825 212.095 ;
        RECT 75.120 211.925 75.290 212.115 ;
        RECT 75.575 211.925 75.745 212.115 ;
        RECT 78.340 211.925 78.510 212.115 ;
        RECT 78.795 211.925 78.965 212.115 ;
        RECT 80.635 211.905 80.805 212.095 ;
        RECT 82.930 211.925 83.100 212.115 ;
        RECT 83.390 211.955 83.510 212.065 ;
        RECT 84.780 211.925 84.950 212.115 ;
        RECT 85.240 211.925 85.410 212.115 ;
        RECT 86.155 211.905 86.325 212.095 ;
        RECT 2.755 211.095 4.125 211.905 ;
        RECT 4.595 211.225 14.965 211.905 ;
        RECT 9.105 211.005 10.035 211.225 ;
        RECT 12.755 210.995 14.965 211.225 ;
        RECT 15.175 211.095 17.925 211.905 ;
        RECT 17.935 211.225 27.215 211.905 ;
        RECT 19.295 211.005 20.215 211.225 ;
        RECT 24.880 211.105 27.215 211.225 ;
        RECT 26.295 210.995 27.215 211.105 ;
        RECT 28.525 211.035 28.955 211.820 ;
        RECT 29.435 211.225 39.805 211.905 ;
        RECT 40.015 211.225 49.205 211.905 ;
        RECT 33.945 211.005 34.875 211.225 ;
        RECT 37.595 210.995 39.805 211.225 ;
        RECT 44.525 211.005 45.455 211.225 ;
        RECT 48.285 210.995 49.205 211.225 ;
        RECT 49.675 211.225 51.505 211.905 ;
        RECT 51.525 211.225 54.265 211.905 ;
        RECT 49.675 210.995 51.020 211.225 ;
        RECT 54.285 211.035 54.715 211.820 ;
        RECT 54.735 211.225 58.635 211.905 ;
        RECT 59.345 211.225 62.085 211.905 ;
        RECT 54.735 210.995 55.665 211.225 ;
        RECT 62.105 210.995 63.455 211.905 ;
        RECT 63.475 211.095 68.985 211.905 ;
        RECT 68.995 211.095 74.505 211.905 ;
        RECT 74.515 211.095 80.025 211.905 ;
        RECT 80.045 211.035 80.475 211.820 ;
        RECT 80.495 211.095 86.005 211.905 ;
        RECT 86.015 211.095 87.845 211.905 ;
        RECT 87.990 211.875 88.160 212.095 ;
        RECT 90.295 211.925 90.465 212.115 ;
        RECT 90.755 211.925 90.925 212.115 ;
        RECT 92.595 212.065 92.765 212.095 ;
        RECT 92.590 211.955 92.765 212.065 ;
        RECT 92.595 211.905 92.765 211.955 ;
        RECT 93.515 211.925 93.685 212.115 ;
        RECT 96.270 211.905 96.440 212.095 ;
        RECT 96.735 211.905 96.905 212.095 ;
        RECT 99.045 211.960 99.205 212.070 ;
        RECT 99.955 211.925 100.125 212.115 ;
        RECT 100.875 211.905 101.045 212.095 ;
        RECT 103.175 211.925 103.345 212.115 ;
        RECT 104.560 212.095 104.730 212.115 ;
        RECT 104.555 211.925 104.730 212.095 ;
        RECT 104.555 211.905 104.725 211.925 ;
        RECT 106.395 211.905 106.565 212.095 ;
        RECT 108.235 211.925 108.405 212.115 ;
        RECT 110.995 211.925 111.165 212.115 ;
        RECT 112.830 211.905 113.000 212.095 ;
        RECT 113.295 211.905 113.465 212.095 ;
        RECT 113.755 211.925 113.925 212.115 ;
        RECT 89.190 211.875 90.145 211.905 ;
        RECT 87.865 211.195 90.145 211.875 ;
        RECT 89.190 210.995 90.145 211.195 ;
        RECT 90.155 210.995 92.905 211.905 ;
        RECT 93.110 210.995 96.585 211.905 ;
        RECT 96.595 210.995 100.655 211.905 ;
        RECT 100.735 211.095 104.405 211.905 ;
        RECT 104.415 211.095 105.785 211.905 ;
        RECT 105.805 211.035 106.235 211.820 ;
        RECT 106.255 211.095 109.925 211.905 ;
        RECT 110.225 210.995 113.145 211.905 ;
        RECT 113.155 211.225 116.825 211.905 ;
        RECT 116.980 211.875 117.150 212.095 ;
        RECT 117.435 211.925 117.605 212.115 ;
        RECT 119.275 211.925 119.445 212.115 ;
        RECT 120.655 211.905 120.825 212.095 ;
        RECT 122.960 211.925 123.130 212.115 ;
        RECT 124.795 212.095 124.965 212.115 ;
        RECT 123.410 211.955 123.530 212.065 ;
        RECT 124.795 211.925 124.970 212.095 ;
        RECT 124.800 211.905 124.970 211.925 ;
        RECT 127.090 211.905 127.260 212.095 ;
        RECT 127.555 211.905 127.725 212.095 ;
        RECT 130.315 211.925 130.485 212.115 ;
        RECT 131.230 211.955 131.350 212.065 ;
        RECT 133.990 211.955 134.110 212.065 ;
        RECT 134.445 211.925 134.615 212.115 ;
        RECT 135.380 211.905 135.550 212.095 ;
        RECT 135.835 211.905 136.005 212.095 ;
        RECT 138.595 211.905 138.765 212.115 ;
        RECT 141.815 211.905 141.985 212.095 ;
        RECT 144.110 211.955 144.230 212.065 ;
        RECT 145.045 211.925 145.215 212.115 ;
        RECT 147.335 211.905 147.505 212.095 ;
        RECT 148.255 211.925 148.425 212.115 ;
        RECT 151.015 212.065 151.185 212.115 ;
        RECT 151.010 211.955 151.185 212.065 ;
        RECT 151.015 211.925 151.185 211.955 ;
        RECT 151.480 211.905 151.650 212.095 ;
        RECT 153.775 211.905 153.945 212.095 ;
        RECT 154.230 211.925 154.400 212.115 ;
        RECT 154.690 211.955 154.810 212.065 ;
        RECT 156.080 211.925 156.250 212.115 ;
        RECT 156.530 211.955 156.650 212.065 ;
        RECT 157.915 211.905 158.085 212.115 ;
        RECT 119.555 211.875 120.505 211.905 ;
        RECT 115.895 210.995 116.825 211.225 ;
        RECT 116.835 211.195 120.505 211.875 ;
        RECT 119.555 210.995 120.505 211.195 ;
        RECT 120.525 210.995 123.255 211.905 ;
        RECT 123.735 210.995 125.085 211.905 ;
        RECT 125.195 210.995 127.405 211.905 ;
        RECT 127.415 211.095 131.085 211.905 ;
        RECT 131.565 211.035 131.995 211.820 ;
        RECT 132.015 210.995 135.675 211.905 ;
        RECT 135.695 211.095 138.445 211.905 ;
        RECT 138.535 210.995 141.535 211.905 ;
        RECT 141.675 211.095 147.185 211.905 ;
        RECT 147.195 211.095 150.865 211.905 ;
        RECT 151.335 210.995 153.525 211.905 ;
        RECT 153.635 211.095 156.385 211.905 ;
        RECT 156.855 211.095 158.225 211.905 ;
      LAYER nwell ;
        RECT 2.560 207.875 158.420 210.705 ;
      LAYER pwell ;
        RECT 2.755 206.675 4.125 207.485 ;
        RECT 8.645 207.355 9.575 207.575 ;
        RECT 12.405 207.355 13.325 207.585 ;
        RECT 4.135 206.675 13.325 207.355 ;
        RECT 14.255 206.675 15.625 207.455 ;
        RECT 15.645 206.760 16.075 207.545 ;
        RECT 17.465 207.355 18.385 207.585 ;
        RECT 16.095 206.675 18.385 207.355 ;
        RECT 18.395 207.355 19.325 207.585 ;
        RECT 25.735 207.355 26.665 207.585 ;
        RECT 29.875 207.355 30.805 207.585 ;
        RECT 18.395 206.675 22.295 207.355 ;
        RECT 22.765 206.675 26.665 207.355 ;
        RECT 26.905 206.675 30.805 207.355 ;
        RECT 31.275 207.355 32.205 207.585 ;
        RECT 31.275 206.675 35.175 207.355 ;
        RECT 35.885 206.675 38.625 207.355 ;
        RECT 38.645 206.675 41.385 207.355 ;
        RECT 41.405 206.760 41.835 207.545 ;
        RECT 45.055 207.355 45.985 207.585 ;
        RECT 42.085 206.675 45.985 207.355 ;
        RECT 45.995 206.675 48.735 207.355 ;
        RECT 48.755 206.675 51.495 207.355 ;
        RECT 51.985 206.675 54.725 207.355 ;
        RECT 54.735 206.675 56.105 207.485 ;
        RECT 56.115 206.675 59.785 207.585 ;
        RECT 59.795 206.675 61.165 207.485 ;
        RECT 61.185 206.675 63.915 207.585 ;
        RECT 64.875 206.675 66.225 207.585 ;
        RECT 67.165 206.760 67.595 207.545 ;
        RECT 67.615 206.675 68.985 207.485 ;
        RECT 69.030 207.355 70.405 207.585 ;
        RECT 72.175 207.355 73.125 207.585 ;
        RECT 69.030 206.905 73.125 207.355 ;
        RECT 2.895 206.465 3.065 206.675 ;
        RECT 4.275 206.625 4.445 206.675 ;
        RECT 4.270 206.515 4.445 206.625 ;
        RECT 4.275 206.485 4.445 206.515 ;
        RECT 4.735 206.465 4.905 206.655 ;
        RECT 7.035 206.465 7.205 206.655 ;
        RECT 7.770 206.465 7.940 206.655 ;
        RECT 13.485 206.520 13.645 206.630 ;
        RECT 14.395 206.485 14.565 206.675 ;
        RECT 15.040 206.465 15.210 206.655 ;
        RECT 16.050 206.465 16.220 206.655 ;
        RECT 16.235 206.485 16.405 206.675 ;
        RECT 18.810 206.485 18.980 206.675 ;
        RECT 20.190 206.465 20.360 206.655 ;
        RECT 24.330 206.465 24.500 206.655 ;
        RECT 26.080 206.485 26.250 206.675 ;
        RECT 28.190 206.515 28.310 206.625 ;
        RECT 29.120 206.465 29.290 206.655 ;
        RECT 30.220 206.485 30.390 206.675 ;
        RECT 30.495 206.465 30.665 206.655 ;
        RECT 30.950 206.515 31.070 206.625 ;
        RECT 31.690 206.485 31.860 206.675 ;
        RECT 35.550 206.515 35.670 206.625 ;
        RECT 38.315 206.485 38.485 206.675 ;
        RECT 41.075 206.485 41.245 206.675 ;
        RECT 41.995 206.465 42.165 206.655 ;
        RECT 42.730 206.465 42.900 206.655 ;
        RECT 45.400 206.485 45.570 206.675 ;
        RECT 46.135 206.485 46.305 206.675 ;
        RECT 48.895 206.485 49.065 206.675 ;
        RECT 50.000 206.465 50.170 206.655 ;
        RECT 51.650 206.515 51.770 206.625 ;
        RECT 53.955 206.465 54.125 206.655 ;
        RECT 54.415 206.485 54.585 206.675 ;
        RECT 54.875 206.485 55.045 206.675 ;
        RECT 56.260 206.485 56.430 206.675 ;
        RECT 2.755 205.655 4.125 206.465 ;
        RECT 4.595 205.685 5.965 206.465 ;
        RECT 5.975 205.685 7.345 206.465 ;
        RECT 7.355 205.785 11.255 206.465 ;
        RECT 11.725 205.785 15.625 206.465 ;
        RECT 7.355 205.555 8.285 205.785 ;
        RECT 14.695 205.555 15.625 205.785 ;
        RECT 15.635 205.785 19.535 206.465 ;
        RECT 19.775 205.785 23.675 206.465 ;
        RECT 23.915 205.785 27.815 206.465 ;
        RECT 15.635 205.555 16.565 205.785 ;
        RECT 19.775 205.555 20.705 205.785 ;
        RECT 23.915 205.555 24.845 205.785 ;
        RECT 28.525 205.595 28.955 206.380 ;
        RECT 28.975 205.555 30.325 206.465 ;
        RECT 30.355 205.785 33.095 206.465 ;
        RECT 33.115 205.785 42.305 206.465 ;
        RECT 42.315 205.785 46.215 206.465 ;
        RECT 46.685 205.785 50.585 206.465 ;
        RECT 33.115 205.555 34.035 205.785 ;
        RECT 36.865 205.565 37.795 205.785 ;
        RECT 42.315 205.555 43.245 205.785 ;
        RECT 49.655 205.555 50.585 205.785 ;
        RECT 50.690 205.785 54.155 206.465 ;
        RECT 54.740 206.435 56.140 206.465 ;
        RECT 57.630 206.435 57.800 206.655 ;
        RECT 58.100 206.465 58.270 206.655 ;
        RECT 59.475 206.465 59.645 206.655 ;
        RECT 59.935 206.485 60.105 206.675 ;
        RECT 61.315 206.485 61.485 206.675 ;
        RECT 64.085 206.520 64.245 206.630 ;
        RECT 64.995 206.465 65.165 206.655 ;
        RECT 65.910 206.485 66.080 206.675 ;
        RECT 67.755 206.655 67.925 206.675 ;
        RECT 66.385 206.520 66.545 206.630 ;
        RECT 67.755 206.485 67.930 206.655 ;
        RECT 69.135 206.485 69.305 206.905 ;
        RECT 70.415 206.675 73.125 206.905 ;
        RECT 73.135 206.675 76.055 207.585 ;
        RECT 76.355 206.675 79.275 207.585 ;
        RECT 79.575 206.675 80.945 207.485 ;
        RECT 80.955 206.675 83.875 207.585 ;
        RECT 84.635 206.675 88.305 207.585 ;
        RECT 88.315 206.675 91.985 207.485 ;
        RECT 92.925 206.760 93.355 207.545 ;
        RECT 95.205 207.355 96.125 207.585 ;
        RECT 93.835 206.675 96.125 207.355 ;
        RECT 96.155 206.675 97.505 207.585 ;
        RECT 97.515 206.675 100.265 207.485 ;
        RECT 100.275 206.675 103.195 207.585 ;
        RECT 103.495 206.675 107.165 207.585 ;
        RECT 107.175 206.675 110.095 207.585 ;
        RECT 110.395 206.675 113.315 207.585 ;
        RECT 114.075 206.675 117.745 207.585 ;
        RECT 118.685 206.760 119.115 207.545 ;
        RECT 119.135 206.675 120.485 207.585 ;
        RECT 120.515 206.675 121.885 207.485 ;
        RECT 121.895 206.675 125.105 207.585 ;
        RECT 125.115 206.675 130.625 207.485 ;
        RECT 132.440 207.385 133.385 207.585 ;
        RECT 130.635 206.705 133.385 207.385 ;
        RECT 67.760 206.465 67.930 206.485 ;
        RECT 70.055 206.465 70.225 206.655 ;
        RECT 73.280 206.485 73.450 206.675 ;
        RECT 75.575 206.465 75.745 206.655 ;
        RECT 76.500 206.485 76.670 206.675 ;
        RECT 79.265 206.510 79.425 206.620 ;
        RECT 79.715 206.485 79.885 206.675 ;
        RECT 80.635 206.465 80.805 206.655 ;
        RECT 81.100 206.485 81.270 206.675 ;
        RECT 87.995 206.655 88.165 206.675 ;
        RECT 84.310 206.515 84.430 206.625 ;
        RECT 87.990 206.485 88.165 206.655 ;
        RECT 88.455 206.625 88.625 206.675 ;
        RECT 88.450 206.515 88.625 206.625 ;
        RECT 88.455 206.485 88.625 206.515 ;
        RECT 87.990 206.465 88.160 206.485 ;
        RECT 88.920 206.465 89.090 206.655 ;
        RECT 92.135 206.465 92.305 206.655 ;
        RECT 93.510 206.515 93.630 206.625 ;
        RECT 93.975 206.485 94.145 206.675 ;
        RECT 94.890 206.515 95.010 206.625 ;
        RECT 96.270 206.485 96.440 206.675 ;
        RECT 97.655 206.485 97.825 206.675 ;
        RECT 98.570 206.465 98.740 206.655 ;
        RECT 99.030 206.485 99.200 206.655 ;
        RECT 100.420 206.485 100.590 206.675 ;
        RECT 99.065 206.465 99.200 206.485 ;
        RECT 50.690 205.555 51.610 205.785 ;
        RECT 54.285 205.595 54.715 206.380 ;
        RECT 54.740 205.755 57.945 206.435 ;
        RECT 54.740 205.555 56.140 205.755 ;
        RECT 57.955 205.555 59.305 206.465 ;
        RECT 59.335 205.655 64.845 206.465 ;
        RECT 64.855 205.655 67.605 206.465 ;
        RECT 67.615 205.555 69.805 206.465 ;
        RECT 69.915 205.655 75.425 206.465 ;
        RECT 75.435 205.655 79.105 206.465 ;
        RECT 80.045 205.595 80.475 206.380 ;
        RECT 80.495 205.655 84.165 206.465 ;
        RECT 84.830 205.555 88.305 206.465 ;
        RECT 88.775 205.555 91.695 206.465 ;
        RECT 91.995 205.655 94.745 206.465 ;
        RECT 95.410 205.555 98.885 206.465 ;
        RECT 99.065 205.555 102.565 206.465 ;
        RECT 102.710 206.435 102.880 206.655 ;
        RECT 105.025 206.510 105.185 206.620 ;
        RECT 106.395 206.465 106.565 206.655 ;
        RECT 106.855 206.485 107.025 206.675 ;
        RECT 107.320 206.485 107.490 206.675 ;
        RECT 108.240 206.465 108.410 206.655 ;
        RECT 110.540 206.485 110.710 206.675 ;
        RECT 112.370 206.465 112.540 206.655 ;
        RECT 112.835 206.485 113.005 206.655 ;
        RECT 113.750 206.515 113.870 206.625 ;
        RECT 114.220 206.485 114.390 206.675 ;
        RECT 112.855 206.465 113.005 206.485 ;
        RECT 115.135 206.465 115.305 206.655 ;
        RECT 117.905 206.520 118.065 206.630 ;
        RECT 120.200 206.485 120.370 206.675 ;
        RECT 120.655 206.465 120.825 206.675 ;
        RECT 122.035 206.485 122.205 206.675 ;
        RECT 123.410 206.515 123.530 206.625 ;
        RECT 123.880 206.465 124.050 206.655 ;
        RECT 125.255 206.485 125.425 206.675 ;
        RECT 127.095 206.465 127.265 206.655 ;
        RECT 130.780 206.485 130.950 206.705 ;
        RECT 132.440 206.675 133.385 206.705 ;
        RECT 133.405 206.675 136.135 207.585 ;
        RECT 136.155 206.675 141.665 207.485 ;
        RECT 141.675 206.675 144.425 207.485 ;
        RECT 144.445 206.760 144.875 207.545 ;
        RECT 145.065 206.675 148.565 207.585 ;
        RECT 149.575 206.675 153.025 207.585 ;
        RECT 153.175 207.355 154.095 207.585 ;
        RECT 153.175 206.675 155.465 207.355 ;
        RECT 155.475 206.675 156.845 207.485 ;
        RECT 156.855 206.675 158.225 207.485 ;
        RECT 133.535 206.655 133.705 206.675 ;
        RECT 132.155 206.465 132.325 206.655 ;
        RECT 133.530 206.485 133.705 206.655 ;
        RECT 133.530 206.465 133.700 206.485 ;
        RECT 134.920 206.465 135.090 206.655 ;
        RECT 136.295 206.485 136.465 206.675 ;
        RECT 136.755 206.465 136.925 206.655 ;
        RECT 141.815 206.485 141.985 206.675 ;
        RECT 145.065 206.655 145.200 206.675 ;
        RECT 142.275 206.465 142.445 206.655 ;
        RECT 145.030 206.485 145.200 206.655 ;
        RECT 146.875 206.465 147.045 206.655 ;
        RECT 147.335 206.465 147.505 206.655 ;
        RECT 148.725 206.520 148.885 206.630 ;
        RECT 149.635 206.485 149.805 206.675 ;
        RECT 152.855 206.465 153.025 206.655 ;
        RECT 155.155 206.485 155.325 206.675 ;
        RECT 155.615 206.485 155.785 206.675 ;
        RECT 156.530 206.515 156.650 206.625 ;
        RECT 157.915 206.465 158.085 206.675 ;
        RECT 103.910 206.435 104.865 206.465 ;
        RECT 102.585 205.755 104.865 206.435 ;
        RECT 103.910 205.555 104.865 205.755 ;
        RECT 105.805 205.595 106.235 206.380 ;
        RECT 106.255 205.655 108.085 206.465 ;
        RECT 108.095 205.555 109.445 206.465 ;
        RECT 109.765 205.555 112.685 206.465 ;
        RECT 112.855 205.645 114.785 206.465 ;
        RECT 114.995 205.655 120.505 206.465 ;
        RECT 120.515 205.655 123.265 206.465 ;
        RECT 113.835 205.555 114.785 205.645 ;
        RECT 123.735 205.555 126.655 206.465 ;
        RECT 126.955 205.655 130.625 206.465 ;
        RECT 131.565 205.595 131.995 206.380 ;
        RECT 132.015 205.655 133.385 206.465 ;
        RECT 133.415 205.555 134.765 206.465 ;
        RECT 134.775 205.555 136.605 206.465 ;
        RECT 136.615 205.655 142.125 206.465 ;
        RECT 142.135 205.655 143.965 206.465 ;
        RECT 144.105 205.555 147.105 206.465 ;
        RECT 147.195 205.655 152.705 206.465 ;
        RECT 152.715 205.655 156.385 206.465 ;
        RECT 156.855 205.655 158.225 206.465 ;
      LAYER nwell ;
        RECT 2.560 202.435 158.420 205.265 ;
      LAYER pwell ;
        RECT 2.755 201.235 4.125 202.045 ;
        RECT 9.565 201.915 10.495 202.135 ;
        RECT 13.325 201.915 14.245 202.145 ;
        RECT 5.055 201.235 14.245 201.915 ;
        RECT 14.255 201.235 15.625 202.015 ;
        RECT 15.645 201.320 16.075 202.105 ;
        RECT 16.135 201.235 19.305 202.145 ;
        RECT 19.315 201.235 21.130 202.145 ;
        RECT 22.205 201.915 23.135 202.145 ;
        RECT 27.575 201.915 28.505 202.145 ;
        RECT 21.300 201.235 23.135 201.915 ;
        RECT 24.605 201.235 28.505 201.915 ;
        RECT 28.530 201.235 30.345 202.145 ;
        RECT 35.325 201.915 36.255 202.135 ;
        RECT 39.085 201.915 40.005 202.145 ;
        RECT 30.815 201.235 40.005 201.915 ;
        RECT 40.035 201.235 41.385 202.145 ;
        RECT 41.405 201.320 41.835 202.105 ;
        RECT 47.285 201.915 48.215 202.135 ;
        RECT 51.045 201.915 51.965 202.145 ;
        RECT 42.775 201.235 51.965 201.915 ;
        RECT 51.985 201.235 54.715 202.145 ;
        RECT 54.735 201.235 56.105 202.015 ;
        RECT 56.115 201.235 58.865 202.145 ;
        RECT 58.875 201.235 61.625 202.145 ;
        RECT 62.555 201.235 66.225 202.145 ;
        RECT 67.165 201.320 67.595 202.105 ;
        RECT 67.615 201.235 68.985 202.045 ;
        RECT 69.125 201.235 72.125 202.145 ;
        RECT 72.295 201.235 75.295 202.145 ;
        RECT 76.090 201.235 79.565 202.145 ;
        RECT 79.575 201.235 81.345 202.145 ;
        RECT 81.415 201.235 84.165 202.045 ;
        RECT 84.175 201.945 85.105 202.145 ;
        RECT 86.440 201.945 87.385 202.145 ;
        RECT 84.175 201.465 87.385 201.945 ;
        RECT 84.315 201.265 87.385 201.465 ;
        RECT 2.895 201.025 3.065 201.235 ;
        RECT 4.275 201.025 4.445 201.215 ;
        RECT 5.195 201.045 5.365 201.235 ;
        RECT 13.475 201.025 13.645 201.215 ;
        RECT 15.315 201.045 15.485 201.235 ;
        RECT 16.235 201.045 16.405 201.235 ;
        RECT 20.835 201.045 21.005 201.235 ;
        RECT 21.300 201.215 21.465 201.235 ;
        RECT 21.295 201.045 21.465 201.215 ;
        RECT 22.680 201.025 22.850 201.215 ;
        RECT 23.605 201.080 23.765 201.190 ;
        RECT 27.920 201.045 28.090 201.235 ;
        RECT 28.190 201.075 28.310 201.185 ;
        RECT 28.655 201.045 28.825 201.235 ;
        RECT 30.495 201.185 30.665 201.215 ;
        RECT 30.955 201.185 31.125 201.235 ;
        RECT 29.110 201.075 29.230 201.185 ;
        RECT 30.490 201.075 30.665 201.185 ;
        RECT 30.950 201.075 31.125 201.185 ;
        RECT 30.495 201.025 30.665 201.075 ;
        RECT 30.955 201.045 31.125 201.075 ;
        RECT 31.690 201.025 31.860 201.215 ;
        RECT 38.960 201.025 39.130 201.215 ;
        RECT 39.690 201.075 39.810 201.185 ;
        RECT 41.070 201.045 41.240 201.235 ;
        RECT 41.995 201.025 42.165 201.215 ;
        RECT 42.460 201.025 42.630 201.215 ;
        RECT 42.915 201.045 43.085 201.235 ;
        RECT 46.140 201.025 46.310 201.215 ;
        RECT 52.115 201.045 52.285 201.235 ;
        RECT 53.030 201.025 53.200 201.215 ;
        RECT 53.505 201.070 53.665 201.180 ;
        RECT 55.795 201.045 55.965 201.235 ;
        RECT 56.255 201.045 56.425 201.235 ;
        RECT 56.715 201.025 56.885 201.215 ;
        RECT 58.555 201.025 58.725 201.215 ;
        RECT 59.015 201.045 59.185 201.235 ;
        RECT 60.395 201.025 60.565 201.215 ;
        RECT 61.785 201.080 61.945 201.190 ;
        RECT 62.235 201.025 62.405 201.215 ;
        RECT 62.695 201.025 62.865 201.215 ;
        RECT 65.910 201.045 66.080 201.235 ;
        RECT 66.385 201.080 66.545 201.190 ;
        RECT 67.755 201.045 67.925 201.235 ;
        RECT 68.215 201.025 68.385 201.215 ;
        RECT 71.895 201.045 72.065 201.235 ;
        RECT 72.355 201.045 72.525 201.235 ;
        RECT 73.735 201.025 73.905 201.215 ;
        RECT 75.570 201.075 75.690 201.185 ;
        RECT 79.250 201.180 79.420 201.235 ;
        RECT 79.250 201.070 79.425 201.180 ;
        RECT 79.250 201.045 79.420 201.070 ;
        RECT 79.720 201.045 79.890 201.235 ;
        RECT 80.635 201.025 80.805 201.215 ;
        RECT 81.555 201.045 81.725 201.235 ;
        RECT 84.315 201.185 84.485 201.265 ;
        RECT 86.440 201.235 87.385 201.265 ;
        RECT 87.395 201.235 92.905 202.045 ;
        RECT 92.925 201.320 93.355 202.105 ;
        RECT 93.835 201.235 97.045 202.145 ;
        RECT 97.055 201.235 98.885 202.145 ;
        RECT 98.895 201.235 101.645 202.045 ;
        RECT 103.460 201.945 104.405 202.145 ;
        RECT 101.655 201.265 104.405 201.945 ;
        RECT 84.310 201.075 84.485 201.185 ;
        RECT 84.315 201.045 84.485 201.075 ;
        RECT 84.775 201.025 84.945 201.215 ;
        RECT 87.535 201.045 87.705 201.235 ;
        RECT 90.750 201.025 90.920 201.215 ;
        RECT 91.215 201.025 91.385 201.215 ;
        RECT 93.510 201.075 93.630 201.185 ;
        RECT 94.905 201.070 95.065 201.180 ;
        RECT 96.745 201.045 96.915 201.235 ;
        RECT 98.570 201.045 98.740 201.235 ;
        RECT 99.035 201.025 99.205 201.235 ;
        RECT 100.875 201.025 101.045 201.215 ;
        RECT 101.335 201.025 101.505 201.215 ;
        RECT 101.800 201.045 101.970 201.265 ;
        RECT 103.460 201.235 104.405 201.265 ;
        RECT 104.415 201.235 109.925 202.045 ;
        RECT 109.935 201.235 112.685 202.045 ;
        RECT 113.155 201.235 116.365 202.145 ;
        RECT 116.375 201.235 118.205 202.045 ;
        RECT 118.685 201.320 119.115 202.105 ;
        RECT 119.595 201.235 123.725 202.145 ;
        RECT 123.735 201.945 124.680 202.145 ;
        RECT 123.735 201.265 126.485 201.945 ;
        RECT 123.735 201.235 124.680 201.265 ;
        RECT 104.555 201.045 104.725 201.235 ;
        RECT 105.025 201.070 105.185 201.180 ;
        RECT 106.395 201.025 106.565 201.215 ;
        RECT 110.075 201.025 110.245 201.235 ;
        RECT 112.830 201.075 112.950 201.185 ;
        RECT 115.595 201.025 115.765 201.215 ;
        RECT 116.055 201.045 116.225 201.235 ;
        RECT 116.515 201.045 116.685 201.235 ;
        RECT 118.350 201.075 118.470 201.185 ;
        RECT 118.815 201.025 118.985 201.215 ;
        RECT 119.270 201.075 119.390 201.185 ;
        RECT 121.115 201.025 121.285 201.215 ;
        RECT 122.955 201.025 123.125 201.215 ;
        RECT 123.415 201.045 123.585 201.235 ;
        RECT 126.170 201.215 126.340 201.265 ;
        RECT 126.495 201.235 130.165 202.045 ;
        RECT 130.635 201.915 131.975 202.145 ;
        RECT 130.635 201.235 134.765 201.915 ;
        RECT 134.775 201.235 136.605 202.045 ;
        RECT 136.615 201.915 137.535 202.145 ;
        RECT 136.615 201.235 138.905 201.915 ;
        RECT 138.915 201.235 144.425 202.045 ;
        RECT 144.445 201.320 144.875 202.105 ;
        RECT 144.895 201.235 147.635 201.915 ;
        RECT 147.655 201.235 150.405 202.045 ;
        RECT 150.875 201.235 153.795 202.145 ;
        RECT 154.095 201.235 156.845 202.045 ;
        RECT 156.855 201.235 158.225 202.045 ;
        RECT 124.340 201.025 124.510 201.215 ;
        RECT 126.170 201.045 126.345 201.215 ;
        RECT 126.635 201.045 126.805 201.235 ;
        RECT 126.175 201.025 126.345 201.045 ;
        RECT 127.555 201.025 127.725 201.215 ;
        RECT 130.310 201.075 130.430 201.185 ;
        RECT 130.780 201.045 130.950 201.235 ;
        RECT 132.155 201.025 132.325 201.215 ;
        RECT 134.915 201.025 135.085 201.235 ;
        RECT 138.595 201.045 138.765 201.235 ;
        RECT 139.055 201.045 139.225 201.235 ;
        RECT 140.435 201.025 140.605 201.215 ;
        RECT 141.815 201.025 141.985 201.215 ;
        RECT 145.035 201.045 145.205 201.235 ;
        RECT 146.415 201.025 146.585 201.215 ;
        RECT 146.875 201.025 147.045 201.215 ;
        RECT 147.795 201.045 147.965 201.235 ;
        RECT 149.640 201.025 149.810 201.215 ;
        RECT 150.550 201.075 150.670 201.185 ;
        RECT 151.020 201.045 151.190 201.235 ;
        RECT 153.315 201.025 153.485 201.215 ;
        RECT 154.235 201.045 154.405 201.235 ;
        RECT 157.915 201.025 158.085 201.235 ;
        RECT 2.755 200.215 4.125 201.025 ;
        RECT 4.135 200.345 13.325 201.025 ;
        RECT 13.335 200.345 22.525 201.025 ;
        RECT 8.645 200.125 9.575 200.345 ;
        RECT 12.405 200.115 13.325 200.345 ;
        RECT 17.845 200.125 18.775 200.345 ;
        RECT 21.605 200.115 22.525 200.345 ;
        RECT 22.535 200.115 28.045 201.025 ;
        RECT 28.525 200.155 28.955 200.940 ;
        RECT 29.435 200.245 30.805 201.025 ;
        RECT 31.275 200.345 35.175 201.025 ;
        RECT 35.645 200.345 39.545 201.025 ;
        RECT 31.275 200.115 32.205 200.345 ;
        RECT 38.615 200.115 39.545 200.345 ;
        RECT 40.015 200.345 42.305 201.025 ;
        RECT 40.015 200.115 40.935 200.345 ;
        RECT 42.315 200.115 45.970 201.025 ;
        RECT 45.995 200.115 49.650 201.025 ;
        RECT 49.690 200.115 53.345 201.025 ;
        RECT 54.285 200.155 54.715 200.940 ;
        RECT 54.735 200.345 57.025 201.025 ;
        RECT 57.035 200.345 58.865 201.025 ;
        RECT 54.735 200.115 55.655 200.345 ;
        RECT 57.035 200.115 58.380 200.345 ;
        RECT 58.875 200.115 60.690 201.025 ;
        RECT 60.715 200.115 62.530 201.025 ;
        RECT 62.555 200.215 68.065 201.025 ;
        RECT 68.075 200.215 73.585 201.025 ;
        RECT 73.595 200.215 79.105 201.025 ;
        RECT 80.045 200.155 80.475 200.940 ;
        RECT 80.495 200.215 84.165 201.025 ;
        RECT 84.635 200.115 88.765 201.025 ;
        RECT 88.855 200.115 91.065 201.025 ;
        RECT 91.075 200.215 94.745 201.025 ;
        RECT 95.675 200.115 99.345 201.025 ;
        RECT 99.355 200.115 101.170 201.025 ;
        RECT 101.195 200.215 104.865 201.025 ;
        RECT 105.805 200.155 106.235 200.940 ;
        RECT 106.255 200.115 109.925 201.025 ;
        RECT 109.935 200.215 115.445 201.025 ;
        RECT 115.455 200.215 118.205 201.025 ;
        RECT 118.675 200.345 120.965 201.025 ;
        RECT 120.045 200.115 120.965 200.345 ;
        RECT 120.990 200.115 122.805 201.025 ;
        RECT 122.825 200.115 124.175 201.025 ;
        RECT 124.195 200.115 126.025 201.025 ;
        RECT 126.035 200.215 127.405 201.025 ;
        RECT 127.495 200.115 130.495 201.025 ;
        RECT 131.565 200.155 131.995 200.940 ;
        RECT 132.015 200.115 134.765 201.025 ;
        RECT 134.775 200.215 140.285 201.025 ;
        RECT 140.295 200.215 141.665 201.025 ;
        RECT 141.675 200.345 144.885 201.025 ;
        RECT 143.750 200.115 144.885 200.345 ;
        RECT 144.895 200.115 146.710 201.025 ;
        RECT 146.735 200.215 149.485 201.025 ;
        RECT 149.495 200.115 152.970 201.025 ;
        RECT 153.175 200.215 156.845 201.025 ;
        RECT 156.855 200.215 158.225 201.025 ;
      LAYER nwell ;
        RECT 2.560 196.995 158.420 199.825 ;
      LAYER pwell ;
        RECT 2.755 195.795 4.125 196.605 ;
        RECT 4.135 195.795 5.965 196.605 ;
        RECT 5.975 195.795 7.345 196.575 ;
        RECT 7.355 196.475 8.285 196.705 ;
        RECT 14.695 196.475 15.625 196.705 ;
        RECT 7.355 195.795 11.255 196.475 ;
        RECT 11.725 195.795 15.625 196.475 ;
        RECT 15.645 195.880 16.075 196.665 ;
        RECT 16.095 195.795 17.465 196.575 ;
        RECT 17.475 196.475 18.405 196.705 ;
        RECT 17.475 195.795 21.375 196.475 ;
        RECT 21.615 195.795 24.825 196.705 ;
        RECT 32.105 196.475 33.035 196.695 ;
        RECT 35.865 196.475 36.785 196.705 ;
        RECT 39.995 196.475 40.925 196.705 ;
        RECT 24.835 195.795 27.575 196.475 ;
        RECT 27.595 195.795 36.785 196.475 ;
        RECT 37.025 195.795 40.925 196.475 ;
        RECT 41.405 195.880 41.835 196.665 ;
        RECT 42.905 196.475 43.835 196.705 ;
        RECT 42.000 195.795 43.835 196.475 ;
        RECT 44.480 195.795 48.135 196.705 ;
        RECT 48.620 195.795 52.275 196.705 ;
        RECT 52.745 196.475 53.675 196.705 ;
        RECT 55.045 196.475 55.975 196.705 ;
        RECT 57.035 196.475 58.380 196.705 ;
        RECT 52.745 195.795 54.580 196.475 ;
        RECT 55.045 195.795 56.880 196.475 ;
        RECT 57.035 195.795 58.865 196.475 ;
        RECT 59.805 195.795 62.535 196.705 ;
        RECT 62.555 195.795 66.225 196.705 ;
        RECT 67.165 195.880 67.595 196.665 ;
        RECT 68.535 195.795 72.190 196.705 ;
        RECT 72.225 195.795 74.955 196.705 ;
        RECT 74.975 195.795 76.805 196.605 ;
        RECT 77.470 195.795 80.945 196.705 ;
        RECT 80.955 195.795 84.625 196.605 ;
        RECT 85.095 195.795 88.015 196.705 ;
        RECT 88.315 195.795 89.685 196.605 ;
        RECT 89.695 195.795 91.905 196.705 ;
        RECT 92.925 195.880 93.355 196.665 ;
        RECT 93.395 195.795 94.745 196.705 ;
        RECT 95.215 196.475 96.135 196.705 ;
        RECT 95.215 195.795 97.505 196.475 ;
        RECT 97.515 195.795 103.025 196.605 ;
        RECT 103.495 195.795 105.325 196.705 ;
        RECT 105.335 195.795 108.545 196.705 ;
        RECT 109.555 195.795 112.555 196.705 ;
        RECT 112.695 195.795 118.205 196.605 ;
        RECT 118.685 195.880 119.115 196.665 ;
        RECT 119.135 195.795 124.645 196.605 ;
        RECT 125.115 195.795 127.855 196.475 ;
        RECT 127.875 195.795 131.545 196.605 ;
        RECT 132.015 195.795 135.685 196.705 ;
        RECT 136.155 195.795 139.365 196.705 ;
        RECT 139.395 195.795 140.745 196.705 ;
        RECT 140.755 195.795 144.425 196.605 ;
        RECT 144.445 195.880 144.875 196.665 ;
        RECT 144.895 195.795 150.405 196.605 ;
        RECT 150.415 195.795 154.070 196.705 ;
        RECT 154.095 195.795 156.845 196.605 ;
        RECT 156.855 195.795 158.225 196.605 ;
        RECT 2.895 195.585 3.065 195.795 ;
        RECT 4.275 195.585 4.445 195.795 ;
        RECT 7.035 195.605 7.205 195.795 ;
        RECT 7.770 195.605 7.940 195.795 ;
        RECT 13.475 195.585 13.645 195.775 ;
        RECT 15.040 195.605 15.210 195.795 ;
        RECT 15.315 195.585 15.485 195.775 ;
        RECT 17.155 195.605 17.325 195.795 ;
        RECT 17.890 195.605 18.060 195.795 ;
        RECT 21.755 195.605 21.925 195.795 ;
        RECT 24.975 195.605 25.145 195.795 ;
        RECT 26.815 195.585 26.985 195.775 ;
        RECT 27.275 195.585 27.445 195.775 ;
        RECT 27.735 195.605 27.905 195.795 ;
        RECT 29.115 195.585 29.285 195.775 ;
        RECT 38.590 195.585 38.760 195.775 ;
        RECT 40.340 195.605 40.510 195.795 ;
        RECT 42.000 195.775 42.165 195.795 ;
        RECT 47.975 195.775 48.135 195.795 ;
        RECT 52.115 195.775 52.275 195.795 ;
        RECT 54.415 195.775 54.580 195.795 ;
        RECT 56.715 195.775 56.880 195.795 ;
        RECT 41.070 195.635 41.190 195.745 ;
        RECT 41.995 195.605 42.165 195.775 ;
        RECT 42.455 195.585 42.625 195.775 ;
        RECT 46.130 195.635 46.250 195.745 ;
        RECT 47.975 195.605 48.145 195.775 ;
        RECT 50.275 195.605 50.445 195.775 ;
        RECT 52.115 195.605 52.285 195.775 ;
        RECT 50.275 195.585 50.435 195.605 ;
        RECT 53.950 195.585 54.120 195.775 ;
        RECT 54.415 195.605 54.585 195.775 ;
        RECT 56.715 195.605 56.885 195.775 ;
        RECT 58.095 195.585 58.265 195.775 ;
        RECT 58.555 195.605 58.725 195.795 ;
        RECT 59.025 195.640 59.185 195.750 ;
        RECT 59.935 195.605 60.105 195.795 ;
        RECT 61.325 195.585 61.495 195.775 ;
        RECT 61.770 195.585 61.940 195.775 ;
        RECT 62.695 195.605 62.865 195.795 ;
        RECT 63.150 195.635 63.270 195.745 ;
        RECT 63.620 195.585 63.790 195.775 ;
        RECT 66.385 195.640 66.545 195.750 ;
        RECT 66.835 195.585 67.005 195.775 ;
        RECT 67.765 195.640 67.925 195.750 ;
        RECT 68.680 195.605 68.850 195.795 ;
        RECT 71.430 195.585 71.600 195.775 ;
        RECT 71.895 195.585 72.065 195.775 ;
        RECT 72.355 195.605 72.525 195.795 ;
        RECT 75.115 195.585 75.285 195.795 ;
        RECT 80.630 195.775 80.800 195.795 ;
        RECT 76.950 195.635 77.070 195.745 ;
        RECT 78.795 195.585 78.965 195.775 ;
        RECT 80.630 195.605 80.805 195.775 ;
        RECT 81.095 195.605 81.265 195.795 ;
        RECT 84.780 195.745 84.950 195.775 ;
        RECT 84.770 195.635 84.950 195.745 ;
        RECT 80.635 195.585 80.805 195.605 ;
        RECT 84.780 195.585 84.950 195.635 ;
        RECT 85.240 195.605 85.410 195.795 ;
        RECT 87.070 195.585 87.240 195.775 ;
        RECT 87.535 195.585 87.705 195.775 ;
        RECT 88.455 195.605 88.625 195.795 ;
        RECT 89.840 195.605 90.010 195.795 ;
        RECT 92.145 195.640 92.305 195.750 ;
        RECT 93.055 195.585 93.225 195.775 ;
        RECT 93.510 195.605 93.680 195.795 ;
        RECT 94.890 195.635 95.010 195.745 ;
        RECT 96.735 195.585 96.905 195.775 ;
        RECT 97.195 195.605 97.365 195.795 ;
        RECT 97.655 195.605 97.825 195.795 ;
        RECT 100.420 195.585 100.590 195.775 ;
        RECT 101.800 195.585 101.970 195.775 ;
        RECT 102.255 195.585 102.425 195.775 ;
        RECT 103.170 195.635 103.290 195.745 ;
        RECT 103.640 195.605 103.810 195.795 ;
        RECT 105.480 195.605 105.650 195.795 ;
        RECT 106.395 195.585 106.565 195.775 ;
        RECT 108.705 195.640 108.865 195.750 ;
        RECT 109.615 195.605 109.785 195.795 ;
        RECT 2.755 194.775 4.125 195.585 ;
        RECT 4.135 194.905 13.325 195.585 ;
        RECT 8.645 194.685 9.575 194.905 ;
        RECT 12.405 194.675 13.325 194.905 ;
        RECT 13.335 194.775 15.165 195.585 ;
        RECT 15.175 194.905 24.365 195.585 ;
        RECT 24.385 194.905 27.125 195.585 ;
        RECT 19.685 194.685 20.615 194.905 ;
        RECT 23.445 194.675 24.365 194.905 ;
        RECT 27.135 194.805 28.505 195.585 ;
        RECT 28.525 194.715 28.955 195.500 ;
        RECT 28.975 194.905 38.165 195.585 ;
        RECT 33.485 194.685 34.415 194.905 ;
        RECT 37.245 194.675 38.165 194.905 ;
        RECT 38.175 194.905 42.075 195.585 ;
        RECT 42.425 194.905 45.890 195.585 ;
        RECT 38.175 194.675 39.105 194.905 ;
        RECT 44.970 194.675 45.890 194.905 ;
        RECT 46.780 194.675 50.435 195.585 ;
        RECT 50.610 194.675 54.265 195.585 ;
        RECT 54.285 194.715 54.715 195.500 ;
        RECT 54.830 194.905 58.295 195.585 ;
        RECT 54.830 194.675 55.750 194.905 ;
        RECT 58.415 194.675 61.625 195.585 ;
        RECT 61.655 194.675 63.005 195.585 ;
        RECT 63.475 194.675 66.395 195.585 ;
        RECT 66.695 194.775 70.365 195.585 ;
        RECT 70.395 194.675 71.745 195.585 ;
        RECT 71.835 194.675 74.835 195.585 ;
        RECT 74.975 194.775 78.645 195.585 ;
        RECT 78.655 194.775 80.025 195.585 ;
        RECT 80.045 194.715 80.475 195.500 ;
        RECT 80.495 194.675 83.705 195.585 ;
        RECT 83.715 194.675 85.065 195.585 ;
        RECT 86.035 194.675 87.385 195.585 ;
        RECT 87.395 194.775 92.905 195.585 ;
        RECT 92.915 194.775 96.585 195.585 ;
        RECT 96.605 194.675 99.335 195.585 ;
        RECT 99.355 194.675 100.705 195.585 ;
        RECT 100.735 194.675 102.085 195.585 ;
        RECT 102.115 194.775 105.785 195.585 ;
        RECT 105.805 194.715 106.235 195.500 ;
        RECT 106.255 194.775 109.925 195.585 ;
        RECT 110.080 195.555 110.250 195.775 ;
        RECT 112.835 195.605 113.005 195.795 ;
        RECT 113.305 195.630 113.465 195.740 ;
        RECT 114.215 195.585 114.385 195.775 ;
        RECT 117.895 195.585 118.065 195.775 ;
        RECT 118.350 195.635 118.470 195.745 ;
        RECT 119.275 195.605 119.445 195.795 ;
        RECT 121.570 195.585 121.740 195.775 ;
        RECT 124.790 195.635 124.910 195.745 ;
        RECT 125.255 195.585 125.425 195.795 ;
        RECT 112.210 195.555 113.145 195.585 ;
        RECT 110.080 195.355 113.145 195.555 ;
        RECT 109.935 194.875 113.145 195.355 ;
        RECT 109.935 194.675 110.865 194.875 ;
        RECT 112.195 194.675 113.145 194.875 ;
        RECT 114.075 194.675 117.745 195.585 ;
        RECT 117.755 194.775 121.425 195.585 ;
        RECT 121.455 194.675 122.805 195.585 ;
        RECT 122.825 194.905 125.565 195.585 ;
        RECT 125.715 195.555 125.885 195.775 ;
        RECT 128.015 195.605 128.185 195.795 ;
        RECT 129.850 195.585 130.020 195.775 ;
        RECT 130.315 195.585 130.485 195.775 ;
        RECT 131.690 195.635 131.810 195.745 ;
        RECT 132.160 195.585 132.330 195.775 ;
        RECT 135.375 195.605 135.545 195.795 ;
        RECT 135.830 195.635 135.950 195.745 ;
        RECT 136.760 195.585 136.930 195.775 ;
        RECT 137.215 195.585 137.385 195.775 ;
        RECT 139.065 195.605 139.235 195.795 ;
        RECT 139.510 195.605 139.680 195.795 ;
        RECT 139.975 195.585 140.145 195.775 ;
        RECT 140.895 195.605 141.065 195.795 ;
        RECT 141.815 195.585 141.985 195.775 ;
        RECT 144.110 195.585 144.280 195.775 ;
        RECT 144.570 195.585 144.740 195.775 ;
        RECT 145.035 195.605 145.205 195.795 ;
        RECT 148.255 195.585 148.425 195.775 ;
        RECT 150.560 195.605 150.730 195.795 ;
        RECT 153.775 195.585 153.945 195.775 ;
        RECT 154.235 195.605 154.405 195.795 ;
        RECT 156.530 195.635 156.650 195.745 ;
        RECT 157.915 195.585 158.085 195.795 ;
        RECT 126.930 195.555 128.325 195.585 ;
        RECT 125.590 194.875 128.325 195.555 ;
        RECT 126.915 194.675 128.325 194.875 ;
        RECT 128.335 194.675 130.165 195.585 ;
        RECT 130.175 194.775 131.545 195.585 ;
        RECT 131.565 194.715 131.995 195.500 ;
        RECT 132.015 194.675 135.490 195.585 ;
        RECT 135.695 194.675 137.045 195.585 ;
        RECT 137.075 194.775 139.825 195.585 ;
        RECT 139.835 194.905 141.665 195.585 ;
        RECT 140.320 194.675 141.665 194.905 ;
        RECT 141.675 194.775 143.045 195.585 ;
        RECT 143.075 194.675 144.425 195.585 ;
        RECT 144.445 194.675 148.105 195.585 ;
        RECT 148.115 194.775 153.625 195.585 ;
        RECT 153.635 194.775 156.385 195.585 ;
        RECT 156.855 194.775 158.225 195.585 ;
      LAYER nwell ;
        RECT 2.560 191.555 158.420 194.385 ;
      LAYER pwell ;
        RECT 2.755 190.355 4.125 191.165 ;
        RECT 4.135 190.355 5.965 191.165 ;
        RECT 5.975 190.355 7.345 191.135 ;
        RECT 7.355 191.035 8.285 191.265 ;
        RECT 11.495 191.035 12.425 191.265 ;
        RECT 7.355 190.355 11.255 191.035 ;
        RECT 11.495 190.355 15.395 191.035 ;
        RECT 15.645 190.440 16.075 191.225 ;
        RECT 16.555 191.035 17.485 191.265 ;
        RECT 23.895 191.035 24.825 191.265 ;
        RECT 28.035 191.035 28.965 191.265 ;
        RECT 33.485 191.035 34.415 191.255 ;
        RECT 37.245 191.035 38.165 191.265 ;
        RECT 40.235 191.175 41.185 191.265 ;
        RECT 16.555 190.355 20.455 191.035 ;
        RECT 20.925 190.355 24.825 191.035 ;
        RECT 25.065 190.355 28.965 191.035 ;
        RECT 28.975 190.355 38.165 191.035 ;
        RECT 39.255 190.355 41.185 191.175 ;
        RECT 41.405 190.440 41.835 191.225 ;
        RECT 41.855 191.035 42.785 191.265 ;
        RECT 52.345 191.035 53.275 191.255 ;
        RECT 56.105 191.035 57.025 191.265 ;
        RECT 41.855 190.355 45.755 191.035 ;
        RECT 45.995 190.355 47.825 191.035 ;
        RECT 47.835 190.355 57.025 191.035 ;
        RECT 57.035 191.035 57.965 191.265 ;
        RECT 57.035 190.355 60.935 191.035 ;
        RECT 61.175 190.355 62.525 191.265 ;
        RECT 63.475 191.035 64.405 191.265 ;
        RECT 63.475 190.355 67.145 191.035 ;
        RECT 67.165 190.440 67.595 191.225 ;
        RECT 67.615 190.355 71.285 191.165 ;
        RECT 71.295 190.355 72.665 191.165 ;
        RECT 72.675 190.355 74.025 191.265 ;
        RECT 74.055 190.355 75.405 191.265 ;
        RECT 75.435 190.355 80.945 191.165 ;
        RECT 80.955 190.355 84.625 191.165 ;
        RECT 84.635 190.355 86.005 191.165 ;
        RECT 86.015 190.355 89.515 191.265 ;
        RECT 89.695 190.355 92.445 191.165 ;
        RECT 92.925 190.440 93.355 191.225 ;
        RECT 93.570 190.355 97.045 191.265 ;
        RECT 97.055 190.355 100.725 191.265 ;
        RECT 100.735 190.355 102.105 191.165 ;
        RECT 102.115 190.355 104.305 191.265 ;
        RECT 104.415 190.355 105.785 191.165 ;
        RECT 107.600 191.065 108.545 191.265 ;
        RECT 105.795 190.385 108.545 191.065 ;
        RECT 2.895 190.145 3.065 190.355 ;
        RECT 4.275 190.305 4.445 190.355 ;
        RECT 4.270 190.195 4.445 190.305 ;
        RECT 4.275 190.165 4.445 190.195 ;
        RECT 4.735 190.145 4.905 190.335 ;
        RECT 6.115 190.145 6.285 190.335 ;
        RECT 7.035 190.165 7.205 190.355 ;
        RECT 7.770 190.165 7.940 190.355 ;
        RECT 11.910 190.165 12.080 190.355 ;
        RECT 15.310 190.195 15.430 190.305 ;
        RECT 15.775 190.145 15.945 190.335 ;
        RECT 16.230 190.195 16.350 190.305 ;
        RECT 16.970 190.165 17.140 190.355 ;
        RECT 17.155 190.145 17.325 190.335 ;
        RECT 24.240 190.165 24.410 190.355 ;
        RECT 26.815 190.145 26.985 190.335 ;
        RECT 28.380 190.165 28.550 190.355 ;
        RECT 29.115 190.145 29.285 190.355 ;
        RECT 39.255 190.335 39.405 190.355 ;
        RECT 31.870 190.195 31.990 190.305 ;
        RECT 33.250 190.145 33.420 190.335 ;
        RECT 35.095 190.145 35.265 190.335 ;
        RECT 35.565 190.190 35.725 190.300 ;
        RECT 38.325 190.200 38.485 190.310 ;
        RECT 39.235 190.165 39.405 190.335 ;
        RECT 42.270 190.165 42.440 190.355 ;
        RECT 45.215 190.145 45.385 190.335 ;
        RECT 47.515 190.165 47.685 190.355 ;
        RECT 47.975 190.165 48.145 190.355 ;
        RECT 49.355 190.165 49.525 190.335 ;
        RECT 49.825 190.190 49.985 190.300 ;
        RECT 49.355 190.145 49.515 190.165 ;
        RECT 50.735 190.145 50.905 190.335 ;
        RECT 54.880 190.145 55.050 190.335 ;
        RECT 57.450 190.165 57.620 190.355 ;
        RECT 59.660 190.145 59.830 190.335 ;
        RECT 61.320 190.165 61.490 190.355 ;
        RECT 62.235 190.145 62.405 190.335 ;
        RECT 62.705 190.200 62.865 190.310 ;
        RECT 2.755 189.335 4.125 190.145 ;
        RECT 4.595 189.365 5.965 190.145 ;
        RECT 5.975 189.465 15.165 190.145 ;
        RECT 10.485 189.245 11.415 189.465 ;
        RECT 14.245 189.235 15.165 189.465 ;
        RECT 15.635 189.365 17.005 190.145 ;
        RECT 17.015 189.465 26.625 190.145 ;
        RECT 21.525 189.245 22.455 189.465 ;
        RECT 25.285 189.235 26.625 189.465 ;
        RECT 26.675 189.335 28.505 190.145 ;
        RECT 28.525 189.275 28.955 190.060 ;
        RECT 28.975 189.335 31.725 190.145 ;
        RECT 32.215 189.235 33.565 190.145 ;
        RECT 33.575 189.465 35.405 190.145 ;
        RECT 36.420 189.465 45.525 190.145 ;
        RECT 45.860 189.235 49.515 190.145 ;
        RECT 50.705 189.465 54.170 190.145 ;
        RECT 53.250 189.235 54.170 189.465 ;
        RECT 54.285 189.275 54.715 190.060 ;
        RECT 54.735 189.235 56.085 190.145 ;
        RECT 56.345 189.465 60.245 190.145 ;
        RECT 59.315 189.235 60.245 189.465 ;
        RECT 60.255 189.465 62.545 190.145 ;
        RECT 62.555 190.115 63.505 190.145 ;
        RECT 65.910 190.115 66.080 190.335 ;
        RECT 66.375 190.145 66.545 190.335 ;
        RECT 66.835 190.165 67.005 190.355 ;
        RECT 67.755 190.165 67.925 190.355 ;
        RECT 69.135 190.145 69.305 190.335 ;
        RECT 70.975 190.145 71.145 190.335 ;
        RECT 71.435 190.165 71.605 190.355 ;
        RECT 73.740 190.335 73.910 190.355 ;
        RECT 72.825 190.190 72.985 190.300 ;
        RECT 73.735 190.165 73.910 190.335 ;
        RECT 74.200 190.165 74.370 190.355 ;
        RECT 75.575 190.165 75.745 190.355 ;
        RECT 73.740 190.145 73.905 190.165 ;
        RECT 77.870 190.145 78.040 190.335 ;
        RECT 78.335 190.145 78.505 190.335 ;
        RECT 80.630 190.145 80.800 190.335 ;
        RECT 81.095 190.165 81.265 190.355 ;
        RECT 84.315 190.145 84.485 190.335 ;
        RECT 84.775 190.165 84.945 190.355 ;
        RECT 89.380 190.335 89.515 190.355 ;
        RECT 86.615 190.145 86.785 190.335 ;
        RECT 89.380 190.165 89.550 190.335 ;
        RECT 89.835 190.165 90.005 190.355 ;
        RECT 90.290 190.195 90.410 190.305 ;
        RECT 92.590 190.195 92.710 190.305 ;
        RECT 93.970 190.145 94.140 190.335 ;
        RECT 94.440 190.145 94.610 190.335 ;
        RECT 96.730 190.165 96.900 190.355 ;
        RECT 97.200 190.165 97.370 190.355 ;
        RECT 98.120 190.145 98.290 190.335 ;
        RECT 98.575 190.145 98.745 190.335 ;
        RECT 100.875 190.165 101.045 190.355 ;
        RECT 102.260 190.165 102.430 190.355 ;
        RECT 104.555 190.165 104.725 190.355 ;
        RECT 105.010 190.145 105.180 190.335 ;
        RECT 105.470 190.195 105.590 190.305 ;
        RECT 105.940 190.165 106.110 190.385 ;
        RECT 107.600 190.355 108.545 190.385 ;
        RECT 108.555 190.355 112.225 191.165 ;
        RECT 112.695 190.355 114.985 191.265 ;
        RECT 114.995 190.355 118.665 191.165 ;
        RECT 118.685 190.440 119.115 191.225 ;
        RECT 119.135 191.065 120.080 191.265 ;
        RECT 119.135 190.385 121.885 191.065 ;
        RECT 119.135 190.355 120.080 190.385 ;
        RECT 106.395 190.145 106.565 190.335 ;
        RECT 108.695 190.165 108.865 190.355 ;
        RECT 110.085 190.190 110.245 190.300 ;
        RECT 60.255 189.235 61.175 189.465 ;
        RECT 62.555 189.435 66.225 190.115 ;
        RECT 66.235 189.465 68.975 190.145 ;
        RECT 62.555 189.235 63.505 189.435 ;
        RECT 68.995 189.335 70.825 190.145 ;
        RECT 70.835 189.465 72.665 190.145 ;
        RECT 73.740 189.465 75.575 190.145 ;
        RECT 71.320 189.235 72.665 189.465 ;
        RECT 74.645 189.235 75.575 189.465 ;
        RECT 75.975 189.235 78.185 190.145 ;
        RECT 78.195 189.335 80.025 190.145 ;
        RECT 80.045 189.275 80.475 190.060 ;
        RECT 80.505 189.235 84.165 190.145 ;
        RECT 84.175 189.465 86.465 190.145 ;
        RECT 85.545 189.235 86.465 189.465 ;
        RECT 86.475 189.335 90.145 190.145 ;
        RECT 90.615 189.235 94.285 190.145 ;
        RECT 94.295 189.235 97.045 190.145 ;
        RECT 97.055 189.235 98.405 190.145 ;
        RECT 98.435 189.335 102.105 190.145 ;
        RECT 103.135 189.235 105.325 190.145 ;
        RECT 105.805 189.275 106.235 190.060 ;
        RECT 106.255 189.335 109.925 190.145 ;
        RECT 110.995 190.115 111.165 190.335 ;
        RECT 112.370 190.195 112.490 190.305 ;
        RECT 112.840 190.165 113.010 190.355 ;
        RECT 113.760 190.145 113.930 190.335 ;
        RECT 115.135 190.145 115.305 190.355 ;
        RECT 118.810 190.195 118.930 190.305 ;
        RECT 119.280 190.145 119.450 190.335 ;
        RECT 121.570 190.165 121.740 190.385 ;
        RECT 121.895 190.355 127.405 191.165 ;
        RECT 127.415 190.355 132.925 191.165 ;
        RECT 132.935 190.355 134.765 191.165 ;
        RECT 134.775 191.035 136.115 191.265 ;
        RECT 134.775 190.355 138.905 191.035 ;
        RECT 138.915 190.355 144.425 191.165 ;
        RECT 144.445 190.440 144.875 191.225 ;
        RECT 144.895 190.355 150.405 191.165 ;
        RECT 150.875 191.065 151.820 191.265 ;
        RECT 150.875 190.385 153.625 191.065 ;
        RECT 150.875 190.355 151.820 190.385 ;
        RECT 122.035 190.165 122.205 190.355 ;
        RECT 122.955 190.145 123.125 190.335 ;
        RECT 126.635 190.145 126.805 190.335 ;
        RECT 127.100 190.145 127.270 190.335 ;
        RECT 127.555 190.165 127.725 190.355 ;
        RECT 131.235 190.145 131.405 190.335 ;
        RECT 132.165 190.190 132.325 190.300 ;
        RECT 133.075 190.165 133.245 190.355 ;
        RECT 134.920 190.165 135.090 190.355 ;
        RECT 133.085 190.145 133.245 190.165 ;
        RECT 137.215 190.145 137.385 190.335 ;
        RECT 139.055 190.165 139.225 190.355 ;
        RECT 145.035 190.335 145.205 190.355 ;
        RECT 142.735 190.145 142.905 190.335 ;
        RECT 143.195 190.145 143.365 190.335 ;
        RECT 145.035 190.165 145.210 190.335 ;
        RECT 148.725 190.190 148.885 190.300 ;
        RECT 145.040 190.145 145.210 190.165 ;
        RECT 149.640 190.145 149.810 190.335 ;
        RECT 150.550 190.195 150.670 190.305 ;
        RECT 152.855 190.145 153.025 190.335 ;
        RECT 153.310 190.165 153.480 190.385 ;
        RECT 153.635 190.355 156.385 191.165 ;
        RECT 156.855 190.355 158.225 191.165 ;
        RECT 153.775 190.165 153.945 190.355 ;
        RECT 156.530 190.195 156.650 190.305 ;
        RECT 157.915 190.145 158.085 190.355 ;
        RECT 112.195 190.115 113.575 190.145 ;
        RECT 110.870 189.435 113.575 190.115 ;
        RECT 112.195 189.235 113.575 189.435 ;
        RECT 113.615 189.235 114.965 190.145 ;
        RECT 114.995 189.335 118.665 190.145 ;
        RECT 119.135 189.235 122.790 190.145 ;
        RECT 122.815 189.335 124.185 190.145 ;
        RECT 124.205 189.465 126.945 190.145 ;
        RECT 126.955 189.235 128.785 190.145 ;
        RECT 128.805 189.235 131.535 190.145 ;
        RECT 131.565 189.275 131.995 190.060 ;
        RECT 133.085 189.235 136.740 190.145 ;
        RECT 137.075 189.235 140.285 190.145 ;
        RECT 140.305 189.235 143.035 190.145 ;
        RECT 143.055 189.335 144.885 190.145 ;
        RECT 144.895 189.235 148.370 190.145 ;
        RECT 149.495 189.235 152.415 190.145 ;
        RECT 152.715 189.335 156.385 190.145 ;
        RECT 156.855 189.335 158.225 190.145 ;
      LAYER nwell ;
        RECT 2.560 186.115 158.420 188.945 ;
      LAYER pwell ;
        RECT 2.755 184.915 4.125 185.725 ;
        RECT 5.495 185.595 6.415 185.815 ;
        RECT 12.495 185.715 13.415 185.825 ;
        RECT 11.080 185.595 13.415 185.715 ;
        RECT 4.135 184.915 13.415 185.595 ;
        RECT 13.795 184.915 15.625 185.725 ;
        RECT 15.645 185.000 16.075 185.785 ;
        RECT 16.555 184.915 17.925 185.695 ;
        RECT 18.395 185.595 19.325 185.825 ;
        RECT 27.045 185.595 27.975 185.815 ;
        RECT 30.805 185.595 31.725 185.825 ;
        RECT 18.395 184.915 22.295 185.595 ;
        RECT 22.535 184.915 31.725 185.595 ;
        RECT 31.820 184.915 40.925 185.595 ;
        RECT 41.405 185.000 41.835 185.785 ;
        RECT 41.855 185.595 42.785 185.825 ;
        RECT 41.855 184.915 45.755 185.595 ;
        RECT 45.995 184.915 47.345 185.825 ;
        RECT 47.525 184.915 51.180 185.825 ;
        RECT 56.025 185.595 56.955 185.815 ;
        RECT 59.785 185.595 60.705 185.825 ;
        RECT 51.515 184.915 60.705 185.595 ;
        RECT 61.390 184.915 67.120 185.825 ;
        RECT 67.165 185.000 67.595 185.785 ;
        RECT 67.635 184.915 73.125 185.825 ;
        RECT 73.135 184.915 75.745 185.825 ;
        RECT 75.905 185.735 77.495 185.825 ;
        RECT 75.905 184.915 78.475 185.735 ;
        RECT 78.655 184.915 81.395 185.595 ;
        RECT 81.415 184.915 84.155 185.595 ;
        RECT 84.175 184.915 89.685 185.725 ;
        RECT 89.695 184.915 92.445 185.725 ;
        RECT 92.925 185.000 93.355 185.785 ;
        RECT 93.385 184.915 96.125 185.595 ;
        RECT 96.135 184.915 97.505 185.725 ;
        RECT 98.885 185.595 99.805 185.825 ;
        RECT 97.515 184.915 99.805 185.595 ;
        RECT 99.825 184.915 102.555 185.825 ;
        RECT 102.575 184.915 104.405 185.725 ;
        RECT 104.875 184.915 106.690 185.825 ;
        RECT 106.715 184.915 110.385 185.725 ;
        RECT 110.395 184.915 111.765 185.725 ;
        RECT 113.580 185.625 114.525 185.825 ;
        RECT 111.775 184.945 114.525 185.625 ;
        RECT 2.895 184.705 3.065 184.915 ;
        RECT 4.275 184.705 4.445 184.915 ;
        RECT 7.955 184.705 8.125 184.895 ;
        RECT 8.690 184.705 8.860 184.895 ;
        RECT 13.935 184.725 14.105 184.915 ;
        RECT 15.960 184.705 16.130 184.895 ;
        RECT 16.230 184.755 16.350 184.865 ;
        RECT 17.615 184.725 17.785 184.915 ;
        RECT 18.070 184.755 18.190 184.865 ;
        RECT 18.810 184.725 18.980 184.915 ;
        RECT 22.675 184.725 22.845 184.915 ;
        RECT 25.895 184.705 26.065 184.895 ;
        RECT 26.365 184.750 26.525 184.860 ;
        RECT 28.195 184.705 28.365 184.895 ;
        RECT 29.390 184.705 29.560 184.895 ;
        RECT 36.660 184.705 36.830 184.895 ;
        RECT 40.615 184.725 40.785 184.915 ;
        RECT 40.800 184.705 40.970 184.895 ;
        RECT 41.070 184.755 41.190 184.865 ;
        RECT 41.535 184.725 41.705 184.895 ;
        RECT 42.270 184.725 42.440 184.915 ;
        RECT 41.555 184.705 41.705 184.725 ;
        RECT 43.840 184.705 44.010 184.895 ;
        RECT 46.140 184.725 46.310 184.915 ;
        RECT 47.525 184.895 47.685 184.915 ;
        RECT 47.515 184.725 47.690 184.895 ;
        RECT 51.655 184.725 51.825 184.915 ;
        RECT 2.755 183.895 4.125 184.705 ;
        RECT 4.135 183.895 6.885 184.705 ;
        RECT 6.895 183.925 8.265 184.705 ;
        RECT 8.275 184.025 12.175 184.705 ;
        RECT 12.645 184.025 16.545 184.705 ;
        RECT 8.275 183.795 9.205 184.025 ;
        RECT 15.615 183.795 16.545 184.025 ;
        RECT 16.595 184.025 26.205 184.705 ;
        RECT 16.595 183.795 17.935 184.025 ;
        RECT 20.765 183.805 21.695 184.025 ;
        RECT 27.135 183.925 28.505 184.705 ;
        RECT 28.525 183.835 28.955 184.620 ;
        RECT 28.975 184.025 32.875 184.705 ;
        RECT 33.345 184.025 37.245 184.705 ;
        RECT 37.485 184.025 41.385 184.705 ;
        RECT 28.975 183.795 29.905 184.025 ;
        RECT 36.315 183.795 37.245 184.025 ;
        RECT 40.455 183.795 41.385 184.025 ;
        RECT 41.555 183.885 43.485 184.705 ;
        RECT 42.535 183.795 43.485 183.885 ;
        RECT 43.695 183.795 47.350 184.705 ;
        RECT 47.520 184.675 47.690 184.725 ;
        RECT 53.955 184.705 54.125 184.895 ;
        RECT 54.885 184.750 55.045 184.860 ;
        RECT 55.795 184.725 55.965 184.895 ;
        RECT 59.945 184.750 60.105 184.860 ;
        RECT 60.850 184.755 60.970 184.865 ;
        RECT 55.805 184.705 55.965 184.725 ;
        RECT 63.610 184.705 63.780 184.895 ;
        RECT 66.835 184.725 67.005 184.915 ;
        RECT 69.595 184.705 69.765 184.895 ;
        RECT 70.055 184.725 70.225 184.895 ;
        RECT 72.810 184.725 72.980 184.915 ;
        RECT 73.280 184.725 73.450 184.915 ;
        RECT 78.335 184.895 78.475 184.915 ;
        RECT 78.335 184.725 78.505 184.895 ;
        RECT 78.795 184.725 78.965 184.915 ;
        RECT 81.555 184.895 81.725 184.915 ;
        RECT 79.710 184.705 79.880 184.895 ;
        RECT 81.555 184.725 81.730 184.895 ;
        RECT 82.010 184.755 82.130 184.865 ;
        RECT 81.560 184.705 81.730 184.725 ;
        RECT 82.480 184.705 82.650 184.895 ;
        RECT 84.315 184.725 84.485 184.915 ;
        RECT 86.155 184.725 86.325 184.895 ;
        RECT 88.910 184.755 89.030 184.865 ;
        RECT 86.185 184.705 86.325 184.725 ;
        RECT 89.370 184.705 89.540 184.895 ;
        RECT 89.835 184.725 90.005 184.915 ;
        RECT 90.760 184.705 90.930 184.895 ;
        RECT 92.590 184.755 92.710 184.865 ;
        RECT 94.445 184.750 94.605 184.860 ;
        RECT 95.815 184.725 95.985 184.915 ;
        RECT 96.275 184.725 96.445 184.915 ;
        RECT 97.655 184.725 97.825 184.915 ;
        RECT 99.035 184.705 99.205 184.895 ;
        RECT 99.495 184.705 99.665 184.895 ;
        RECT 99.955 184.725 100.125 184.915 ;
        RECT 102.715 184.895 102.885 184.915 ;
        RECT 102.250 184.755 102.370 184.865 ;
        RECT 102.710 184.725 102.885 184.895 ;
        RECT 104.550 184.755 104.670 184.865 ;
        RECT 105.025 184.750 105.185 184.860 ;
        RECT 106.395 184.725 106.565 184.915 ;
        RECT 106.855 184.725 107.025 184.915 ;
        RECT 49.650 184.675 50.585 184.705 ;
        RECT 47.520 184.475 50.585 184.675 ;
        RECT 47.375 183.995 50.585 184.475 ;
        RECT 47.375 183.795 48.305 183.995 ;
        RECT 49.635 183.795 50.585 183.995 ;
        RECT 50.690 184.025 54.155 184.705 ;
        RECT 50.690 183.795 51.610 184.025 ;
        RECT 54.285 183.835 54.715 184.620 ;
        RECT 55.805 183.795 59.460 184.705 ;
        RECT 60.715 183.795 63.925 184.705 ;
        RECT 64.150 183.795 69.880 184.705 ;
        RECT 70.305 183.795 76.345 184.705 ;
        RECT 76.370 183.795 80.025 184.705 ;
        RECT 80.045 183.835 80.475 184.620 ;
        RECT 80.495 183.795 81.845 184.705 ;
        RECT 82.335 183.795 86.005 184.705 ;
        RECT 86.185 183.885 88.755 184.705 ;
        RECT 87.165 183.795 88.755 183.885 ;
        RECT 89.255 183.795 90.605 184.705 ;
        RECT 90.615 183.795 94.285 184.705 ;
        RECT 95.215 183.795 99.345 184.705 ;
        RECT 99.355 183.895 102.105 184.705 ;
        RECT 102.710 184.675 102.880 184.725 ;
        RECT 107.320 184.705 107.490 184.895 ;
        RECT 110.535 184.725 110.705 184.915 ;
        RECT 110.995 184.705 111.165 184.895 ;
        RECT 111.920 184.725 112.090 184.945 ;
        RECT 113.580 184.915 114.525 184.945 ;
        RECT 114.550 184.915 116.365 185.825 ;
        RECT 116.375 184.915 117.725 185.825 ;
        RECT 118.685 185.000 119.115 185.785 ;
        RECT 119.135 184.915 120.965 185.725 ;
        RECT 123.050 185.595 124.185 185.825 ;
        RECT 120.975 184.915 124.185 185.595 ;
        RECT 125.245 184.915 128.245 185.825 ;
        RECT 128.335 184.915 133.845 185.725 ;
        RECT 133.855 184.915 135.205 185.825 ;
        RECT 135.235 184.915 138.905 185.725 ;
        RECT 138.915 184.915 140.285 185.725 ;
        RECT 141.665 185.595 142.585 185.825 ;
        RECT 140.295 184.915 142.585 185.595 ;
        RECT 142.595 184.915 144.425 185.725 ;
        RECT 144.445 185.000 144.875 185.785 ;
        RECT 144.895 184.915 150.405 185.725 ;
        RECT 150.415 184.915 152.245 185.725 ;
        RECT 152.255 184.915 154.995 185.595 ;
        RECT 155.015 184.915 156.845 185.725 ;
        RECT 156.855 184.915 158.225 185.725 ;
        RECT 114.675 184.725 114.845 184.915 ;
        RECT 116.515 184.705 116.685 184.895 ;
        RECT 117.440 184.725 117.610 184.915 ;
        RECT 117.905 184.760 118.065 184.870 ;
        RECT 118.350 184.755 118.470 184.865 ;
        RECT 119.275 184.725 119.445 184.915 ;
        RECT 121.115 184.725 121.285 184.915 ;
        RECT 121.575 184.705 121.745 184.895 ;
        RECT 122.030 184.755 122.150 184.865 ;
        RECT 124.345 184.760 124.505 184.870 ;
        RECT 125.250 184.725 125.420 184.895 ;
        RECT 125.250 184.705 125.395 184.725 ;
        RECT 127.095 184.705 127.265 184.895 ;
        RECT 127.555 184.705 127.725 184.895 ;
        RECT 128.015 184.725 128.185 184.915 ;
        RECT 128.475 184.725 128.645 184.915 ;
        RECT 129.400 184.705 129.570 184.895 ;
        RECT 132.165 184.750 132.325 184.860 ;
        RECT 133.075 184.705 133.245 184.895 ;
        RECT 134.000 184.725 134.170 184.915 ;
        RECT 135.375 184.725 135.545 184.915 ;
        RECT 135.835 184.705 136.005 184.895 ;
        RECT 137.205 184.705 137.375 184.895 ;
        RECT 139.055 184.725 139.225 184.915 ;
        RECT 140.435 184.705 140.605 184.915 ;
        RECT 142.280 184.705 142.450 184.895 ;
        RECT 142.735 184.725 142.905 184.915 ;
        RECT 144.575 184.705 144.745 184.895 ;
        RECT 145.035 184.725 145.205 184.915 ;
        RECT 148.250 184.755 148.370 184.865 ;
        RECT 148.710 184.705 148.880 184.895 ;
        RECT 150.100 184.705 150.270 184.895 ;
        RECT 150.555 184.725 150.725 184.915 ;
        RECT 152.395 184.725 152.565 184.915 ;
        RECT 153.315 184.705 153.485 184.895 ;
        RECT 155.155 184.725 155.325 184.915 ;
        RECT 156.085 184.750 156.245 184.860 ;
        RECT 157.915 184.705 158.085 184.915 ;
        RECT 103.910 184.675 104.865 184.705 ;
        RECT 102.585 183.995 104.865 184.675 ;
        RECT 103.910 183.795 104.865 183.995 ;
        RECT 105.805 183.835 106.235 184.620 ;
        RECT 107.175 183.795 110.845 184.705 ;
        RECT 110.855 183.895 116.365 184.705 ;
        RECT 116.375 183.895 118.205 184.705 ;
        RECT 118.675 183.795 121.885 184.705 ;
        RECT 122.355 183.795 125.395 184.705 ;
        RECT 125.575 183.795 127.390 184.705 ;
        RECT 127.415 183.895 129.245 184.705 ;
        RECT 129.255 183.795 131.545 184.705 ;
        RECT 131.565 183.835 131.995 184.620 ;
        RECT 132.935 183.795 135.685 184.705 ;
        RECT 135.695 183.895 137.065 184.705 ;
        RECT 137.075 183.795 140.285 184.705 ;
        RECT 140.295 183.895 142.125 184.705 ;
        RECT 142.135 183.795 144.325 184.705 ;
        RECT 144.435 183.895 148.105 184.705 ;
        RECT 148.595 183.795 149.945 184.705 ;
        RECT 149.955 183.795 152.875 184.705 ;
        RECT 153.175 184.025 155.915 184.705 ;
        RECT 156.855 183.895 158.225 184.705 ;
      LAYER nwell ;
        RECT 2.560 180.675 158.420 183.505 ;
      LAYER pwell ;
        RECT 2.755 179.475 4.125 180.285 ;
        RECT 5.495 180.155 6.415 180.375 ;
        RECT 12.495 180.275 13.415 180.385 ;
        RECT 11.080 180.155 13.415 180.275 ;
        RECT 4.135 179.475 13.415 180.155 ;
        RECT 14.255 179.475 15.625 180.255 ;
        RECT 15.645 179.560 16.075 180.345 ;
        RECT 16.465 180.275 17.385 180.385 ;
        RECT 16.465 180.155 18.800 180.275 ;
        RECT 23.465 180.155 24.385 180.375 ;
        RECT 16.465 179.475 25.745 180.155 ;
        RECT 25.755 179.475 27.125 180.255 ;
        RECT 32.105 180.155 33.035 180.375 ;
        RECT 35.865 180.155 36.785 180.385 ;
        RECT 27.595 179.475 36.785 180.155 ;
        RECT 36.795 180.155 37.725 180.385 ;
        RECT 36.795 179.475 40.695 180.155 ;
        RECT 41.405 179.560 41.835 180.345 ;
        RECT 41.855 179.705 46.445 180.385 ;
        RECT 47.505 180.155 48.435 180.385 ;
        RECT 42.815 179.475 46.445 179.705 ;
        RECT 46.600 179.475 48.435 180.155 ;
        RECT 48.755 179.475 52.410 180.385 ;
        RECT 52.445 179.475 55.175 180.385 ;
        RECT 60.625 180.155 61.555 180.375 ;
        RECT 64.275 180.155 66.485 180.385 ;
        RECT 56.115 179.475 66.485 180.155 ;
        RECT 67.165 179.560 67.595 180.345 ;
        RECT 69.420 180.185 70.365 180.385 ;
        RECT 67.615 179.505 70.365 180.185 ;
        RECT 2.895 179.265 3.065 179.475 ;
        RECT 4.275 179.265 4.445 179.475 ;
        RECT 7.035 179.265 7.205 179.455 ;
        RECT 7.495 179.265 7.665 179.455 ;
        RECT 9.610 179.265 9.780 179.455 ;
        RECT 13.475 179.265 13.645 179.455 ;
        RECT 13.930 179.315 14.050 179.425 ;
        RECT 14.395 179.285 14.565 179.475 ;
        RECT 15.590 179.265 15.760 179.455 ;
        RECT 19.455 179.265 19.625 179.455 ;
        RECT 25.435 179.285 25.605 179.475 ;
        RECT 26.815 179.285 26.985 179.475 ;
        RECT 27.270 179.315 27.390 179.425 ;
        RECT 27.735 179.285 27.905 179.475 ;
        RECT 29.125 179.310 29.285 179.420 ;
        RECT 30.955 179.265 31.125 179.455 ;
        RECT 31.415 179.265 31.585 179.455 ;
        RECT 32.795 179.265 32.965 179.455 ;
        RECT 37.210 179.285 37.380 179.475 ;
        RECT 41.070 179.315 41.190 179.425 ;
        RECT 42.910 179.265 43.080 179.455 ;
        RECT 43.375 179.285 43.545 179.455 ;
        RECT 46.130 179.285 46.300 179.475 ;
        RECT 46.600 179.455 46.765 179.475 ;
        RECT 46.595 179.285 46.765 179.455 ;
        RECT 43.380 179.265 43.545 179.285 ;
        RECT 47.515 179.265 47.685 179.455 ;
        RECT 47.980 179.265 48.150 179.455 ;
        RECT 48.900 179.285 49.070 179.475 ;
        RECT 51.655 179.265 51.825 179.455 ;
        RECT 52.575 179.285 52.745 179.475 ;
        RECT 54.870 179.315 54.990 179.425 ;
        RECT 2.755 178.455 4.125 179.265 ;
        RECT 4.135 178.455 5.965 179.265 ;
        RECT 5.975 178.485 7.345 179.265 ;
        RECT 7.355 178.455 9.185 179.265 ;
        RECT 9.195 178.585 13.095 179.265 ;
        RECT 9.195 178.355 10.125 178.585 ;
        RECT 13.335 178.455 15.165 179.265 ;
        RECT 15.175 178.585 19.075 179.265 ;
        RECT 19.315 178.585 28.505 179.265 ;
        RECT 15.175 178.355 16.105 178.585 ;
        RECT 23.825 178.365 24.755 178.585 ;
        RECT 27.585 178.355 28.505 178.585 ;
        RECT 28.525 178.395 28.955 179.180 ;
        RECT 29.895 178.485 31.265 179.265 ;
        RECT 31.275 178.485 32.645 179.265 ;
        RECT 32.655 178.585 41.845 179.265 ;
        RECT 37.165 178.365 38.095 178.585 ;
        RECT 40.925 178.355 41.845 178.585 ;
        RECT 41.875 178.355 43.225 179.265 ;
        RECT 43.380 178.585 45.215 179.265 ;
        RECT 44.285 178.355 45.215 178.585 ;
        RECT 45.535 178.585 47.825 179.265 ;
        RECT 45.535 178.355 46.455 178.585 ;
        RECT 47.835 178.355 51.490 179.265 ;
        RECT 51.515 178.585 54.255 179.265 ;
        RECT 55.340 179.235 55.510 179.455 ;
        RECT 56.255 179.285 56.425 179.475 ;
        RECT 58.555 179.265 58.725 179.455 ;
        RECT 66.830 179.315 66.950 179.425 ;
        RECT 67.760 179.285 67.930 179.505 ;
        RECT 69.420 179.475 70.365 179.505 ;
        RECT 70.375 180.155 71.745 180.385 ;
        RECT 70.375 179.475 74.505 180.155 ;
        RECT 74.515 179.475 75.885 180.285 ;
        RECT 75.980 179.475 85.085 180.155 ;
        RECT 85.095 179.475 88.985 180.385 ;
        RECT 89.245 179.475 91.985 180.155 ;
        RECT 92.925 179.560 93.355 180.345 ;
        RECT 93.470 180.155 94.390 180.385 ;
        RECT 103.035 180.155 103.955 180.385 ;
        RECT 93.470 179.475 96.935 180.155 ;
        RECT 97.055 179.475 99.795 180.155 ;
        RECT 100.275 179.475 103.015 180.155 ;
        RECT 103.035 179.475 105.325 180.155 ;
        RECT 105.335 179.475 109.005 180.285 ;
        RECT 109.015 179.475 110.385 180.285 ;
        RECT 110.395 179.475 114.060 180.385 ;
        RECT 114.075 180.185 115.485 180.385 ;
        RECT 114.075 179.505 116.810 180.185 ;
        RECT 114.075 179.475 115.470 179.505 ;
        RECT 69.135 179.265 69.305 179.455 ;
        RECT 70.505 179.285 70.675 179.475 ;
        RECT 74.655 179.285 74.825 179.475 ;
        RECT 79.250 179.265 79.420 179.455 ;
        RECT 79.710 179.315 79.830 179.425 ;
        RECT 80.640 179.265 80.810 179.455 ;
        RECT 84.310 179.315 84.430 179.425 ;
        RECT 84.775 179.285 84.945 179.475 ;
        RECT 85.240 179.285 85.410 179.475 ;
        RECT 87.990 179.265 88.160 179.455 ;
        RECT 88.460 179.285 88.630 179.455 ;
        RECT 88.485 179.265 88.630 179.285 ;
        RECT 91.675 179.265 91.845 179.475 ;
        RECT 92.145 179.320 92.305 179.430 ;
        RECT 93.515 179.265 93.685 179.455 ;
        RECT 96.735 179.285 96.905 179.475 ;
        RECT 97.195 179.285 97.365 179.475 ;
        RECT 99.960 179.425 100.130 179.455 ;
        RECT 99.950 179.315 100.130 179.425 ;
        RECT 99.960 179.265 100.130 179.315 ;
        RECT 100.415 179.285 100.585 179.475 ;
        RECT 104.095 179.265 104.265 179.455 ;
        RECT 105.015 179.285 105.185 179.475 ;
        RECT 105.475 179.285 105.645 179.475 ;
        RECT 109.155 179.285 109.325 179.475 ;
        RECT 109.610 179.265 109.780 179.455 ;
        RECT 110.075 179.265 110.245 179.455 ;
        RECT 110.540 179.285 110.710 179.475 ;
        RECT 116.515 179.285 116.685 179.505 ;
        RECT 116.835 179.475 118.665 180.285 ;
        RECT 118.685 179.560 119.115 180.345 ;
        RECT 121.210 180.155 122.345 180.385 ;
        RECT 119.135 179.475 122.345 180.155 ;
        RECT 122.815 179.475 125.855 180.385 ;
        RECT 126.955 179.475 129.145 180.385 ;
        RECT 129.255 179.475 134.765 180.285 ;
        RECT 134.775 179.475 136.605 180.285 ;
        RECT 137.075 180.155 138.005 180.385 ;
        RECT 137.075 179.475 140.975 180.155 ;
        RECT 141.215 179.475 143.965 180.285 ;
        RECT 144.445 179.560 144.875 180.345 ;
        RECT 144.895 179.475 150.405 180.285 ;
        RECT 150.875 179.475 153.485 180.385 ;
        RECT 153.635 179.475 156.385 180.285 ;
        RECT 156.855 179.475 158.225 180.285 ;
        RECT 116.975 179.285 117.145 179.475 ;
        RECT 117.895 179.265 118.065 179.455 ;
        RECT 118.355 179.265 118.525 179.455 ;
        RECT 119.275 179.285 119.445 179.475 ;
        RECT 125.710 179.455 125.855 179.475 ;
        RECT 120.190 179.265 120.360 179.455 ;
        RECT 121.575 179.265 121.745 179.455 ;
        RECT 122.490 179.315 122.610 179.425 ;
        RECT 125.250 179.265 125.420 179.455 ;
        RECT 125.710 179.285 125.885 179.455 ;
        RECT 126.185 179.320 126.345 179.430 ;
        RECT 127.100 179.285 127.270 179.475 ;
        RECT 128.470 179.315 128.590 179.425 ;
        RECT 129.395 179.285 129.565 179.475 ;
        RECT 125.715 179.265 125.885 179.285 ;
        RECT 131.235 179.265 131.405 179.455 ;
        RECT 134.915 179.285 135.085 179.475 ;
        RECT 135.375 179.265 135.545 179.455 ;
        RECT 135.835 179.265 136.005 179.455 ;
        RECT 136.750 179.315 136.870 179.425 ;
        RECT 137.490 179.285 137.660 179.475 ;
        RECT 140.900 179.285 141.070 179.455 ;
        RECT 140.900 179.265 141.035 179.285 ;
        RECT 141.355 179.265 141.525 179.475 ;
        RECT 142.740 179.265 142.910 179.455 ;
        RECT 144.110 179.315 144.230 179.425 ;
        RECT 145.035 179.285 145.205 179.475 ;
        RECT 150.550 179.315 150.670 179.425 ;
        RECT 151.020 179.285 151.190 179.475 ;
        RECT 152.385 179.265 152.555 179.455 ;
        RECT 153.775 179.285 153.945 179.475 ;
        RECT 155.615 179.265 155.785 179.455 ;
        RECT 156.530 179.315 156.650 179.425 ;
        RECT 157.915 179.265 158.085 179.475 ;
        RECT 57.000 179.235 58.400 179.265 ;
        RECT 54.285 178.395 54.715 179.180 ;
        RECT 55.195 178.555 58.400 179.235 ;
        RECT 58.415 178.585 68.785 179.265 ;
        RECT 57.000 178.355 58.400 178.555 ;
        RECT 62.925 178.365 63.855 178.585 ;
        RECT 66.575 178.355 68.785 178.585 ;
        RECT 68.995 178.455 71.745 179.265 ;
        RECT 72.005 178.355 79.565 179.265 ;
        RECT 80.045 178.395 80.475 179.180 ;
        RECT 80.495 178.585 84.080 179.265 ;
        RECT 80.495 178.355 81.415 178.585 ;
        RECT 84.635 178.355 88.305 179.265 ;
        RECT 88.485 178.355 91.525 179.265 ;
        RECT 91.535 178.585 93.365 179.265 ;
        RECT 92.020 178.355 93.365 178.585 ;
        RECT 93.375 178.355 99.805 179.265 ;
        RECT 99.815 178.355 103.850 179.265 ;
        RECT 103.955 178.455 105.785 179.265 ;
        RECT 105.805 178.395 106.235 179.180 ;
        RECT 106.255 178.355 109.925 179.265 ;
        RECT 109.935 178.585 112.675 179.265 ;
        RECT 112.895 178.355 118.205 179.265 ;
        RECT 118.215 178.585 120.045 179.265 ;
        RECT 118.700 178.355 120.045 178.585 ;
        RECT 120.075 178.355 121.425 179.265 ;
        RECT 121.435 178.455 123.265 179.265 ;
        RECT 123.375 178.355 125.565 179.265 ;
        RECT 125.575 178.455 128.325 179.265 ;
        RECT 128.805 178.585 131.545 179.265 ;
        RECT 131.565 178.395 131.995 179.180 ;
        RECT 132.015 178.355 135.685 179.265 ;
        RECT 135.695 178.455 137.525 179.265 ;
        RECT 137.535 178.355 141.035 179.265 ;
        RECT 141.215 178.455 142.585 179.265 ;
        RECT 142.595 178.355 152.125 179.265 ;
        RECT 152.255 178.355 155.465 179.265 ;
        RECT 155.475 178.455 156.845 179.265 ;
        RECT 156.855 178.455 158.225 179.265 ;
      LAYER nwell ;
        RECT 2.560 175.235 158.420 178.065 ;
      LAYER pwell ;
        RECT 2.755 174.035 4.125 174.845 ;
        RECT 9.565 174.715 10.495 174.935 ;
        RECT 13.325 174.715 14.245 174.945 ;
        RECT 5.055 174.035 14.245 174.715 ;
        RECT 14.255 174.035 15.625 174.845 ;
        RECT 15.645 174.120 16.075 174.905 ;
        RECT 16.095 174.035 17.465 174.845 ;
        RECT 17.475 174.035 18.845 174.815 ;
        RECT 18.855 174.035 22.065 174.945 ;
        RECT 25.275 174.715 26.205 174.945 ;
        RECT 22.305 174.035 26.205 174.715 ;
        RECT 26.215 174.035 31.725 174.845 ;
        RECT 31.735 174.035 33.105 174.845 ;
        RECT 35.875 174.715 36.805 174.945 ;
        RECT 33.125 174.035 35.865 174.715 ;
        RECT 35.875 174.035 39.775 174.715 ;
        RECT 40.015 174.035 41.385 174.845 ;
        RECT 41.405 174.120 41.835 174.905 ;
        RECT 41.855 174.715 42.785 174.945 ;
        RECT 41.855 174.035 45.755 174.715 ;
        RECT 46.455 174.035 50.110 174.945 ;
        RECT 50.445 174.715 51.375 174.945 ;
        RECT 50.445 174.035 52.280 174.715 ;
        RECT 2.895 173.825 3.065 174.035 ;
        RECT 4.275 173.825 4.445 174.015 ;
        RECT 5.195 173.845 5.365 174.035 ;
        RECT 7.030 173.875 7.150 173.985 ;
        RECT 8.415 173.825 8.585 174.015 ;
        RECT 8.875 173.825 9.045 174.015 ;
        RECT 10.530 173.825 10.700 174.015 ;
        RECT 14.395 173.825 14.565 174.035 ;
        RECT 16.235 173.845 16.405 174.035 ;
        RECT 17.615 173.845 17.785 174.035 ;
        RECT 18.085 173.870 18.245 173.980 ;
        RECT 18.995 173.825 19.165 174.035 ;
        RECT 25.620 173.825 25.790 174.035 ;
        RECT 26.355 173.825 26.525 174.035 ;
        RECT 28.190 173.875 28.310 173.985 ;
        RECT 29.110 173.875 29.230 173.985 ;
        RECT 30.495 173.825 30.665 174.015 ;
        RECT 31.230 173.825 31.400 174.015 ;
        RECT 31.875 173.845 32.045 174.035 ;
        RECT 35.095 173.825 35.265 174.015 ;
        RECT 35.555 173.845 35.725 174.035 ;
        RECT 36.290 173.845 36.460 174.035 ;
        RECT 36.930 173.875 37.050 173.985 ;
        RECT 37.395 173.825 37.565 174.015 ;
        RECT 40.155 173.845 40.325 174.035 ;
        RECT 42.270 173.845 42.440 174.035 ;
        RECT 46.600 174.015 46.770 174.035 ;
        RECT 52.115 174.015 52.280 174.035 ;
        RECT 52.585 174.035 56.240 174.945 ;
        RECT 61.085 174.715 62.015 174.935 ;
        RECT 64.845 174.715 66.185 174.945 ;
        RECT 56.575 174.035 66.185 174.715 ;
        RECT 67.165 174.120 67.595 174.905 ;
        RECT 67.615 174.035 68.985 174.845 ;
        RECT 69.150 174.035 75.310 174.945 ;
        RECT 75.435 174.035 78.645 174.945 ;
        RECT 83.165 174.715 84.095 174.935 ;
        RECT 86.925 174.715 87.845 174.945 ;
        RECT 78.655 174.035 87.845 174.715 ;
        RECT 87.950 174.715 88.870 174.945 ;
        RECT 87.950 174.035 91.415 174.715 ;
        RECT 91.555 174.035 92.905 174.945 ;
        RECT 92.925 174.120 93.355 174.905 ;
        RECT 93.375 174.035 97.030 174.945 ;
        RECT 98.395 174.745 99.805 174.945 ;
        RECT 97.070 174.065 99.805 174.745 ;
        RECT 52.585 174.015 52.745 174.035 ;
        RECT 46.130 173.875 46.250 173.985 ;
        RECT 46.595 173.845 46.770 174.015 ;
        RECT 46.595 173.825 46.765 173.845 ;
        RECT 50.270 173.825 50.440 174.015 ;
        RECT 50.740 173.825 50.910 174.015 ;
        RECT 52.115 173.845 52.285 174.015 ;
        RECT 52.575 173.845 52.745 174.015 ;
        RECT 54.885 173.870 55.045 173.980 ;
        RECT 55.795 173.845 55.965 174.015 ;
        RECT 56.715 173.845 56.885 174.035 ;
        RECT 59.945 173.870 60.105 173.980 ;
        RECT 55.805 173.825 55.965 173.845 ;
        RECT 60.855 173.825 61.025 174.015 ;
        RECT 64.535 173.825 64.705 174.015 ;
        RECT 66.385 173.880 66.545 173.990 ;
        RECT 67.755 173.845 67.925 174.035 ;
        RECT 68.210 173.825 68.380 174.015 ;
        RECT 72.365 173.870 72.525 173.980 ;
        RECT 73.280 173.825 73.450 174.015 ;
        RECT 75.135 173.845 75.305 174.035 ;
        RECT 77.410 173.875 77.530 173.985 ;
        RECT 77.875 173.825 78.045 174.015 ;
        RECT 78.330 173.845 78.500 174.035 ;
        RECT 78.795 173.845 78.965 174.035 ;
        RECT 91.215 174.015 91.385 174.035 ;
        RECT 83.390 173.825 83.560 174.015 ;
        RECT 84.775 173.825 84.945 174.015 ;
        RECT 85.230 173.875 85.350 173.985 ;
        RECT 87.995 173.825 88.165 174.015 ;
        RECT 90.755 173.825 90.925 174.015 ;
        RECT 91.210 173.845 91.385 174.015 ;
        RECT 91.670 173.845 91.840 174.035 ;
        RECT 91.210 173.825 91.380 173.845 ;
        RECT 92.595 173.825 92.765 174.015 ;
        RECT 93.520 173.845 93.690 174.035 ;
        RECT 95.825 173.870 95.985 173.980 ;
        RECT 97.195 173.845 97.365 174.065 ;
        RECT 98.410 174.035 99.805 174.065 ;
        RECT 99.845 174.745 101.225 174.945 ;
        RECT 104.380 174.745 105.325 174.945 ;
        RECT 106.670 174.745 107.625 174.945 ;
        RECT 99.845 174.065 102.550 174.745 ;
        RECT 102.575 174.065 105.325 174.745 ;
        RECT 105.345 174.065 107.625 174.745 ;
        RECT 99.845 174.035 101.225 174.065 ;
        RECT 99.490 173.825 99.660 174.015 ;
        RECT 102.255 173.845 102.425 174.065 ;
        RECT 102.720 174.015 102.890 174.065 ;
        RECT 104.380 174.035 105.325 174.065 ;
        RECT 105.470 174.015 105.640 174.065 ;
        RECT 106.670 174.035 107.625 174.065 ;
        RECT 107.655 174.035 109.005 174.945 ;
        RECT 109.935 174.715 111.280 174.945 ;
        RECT 116.825 174.715 117.745 174.945 ;
        RECT 109.935 174.035 111.765 174.715 ;
        RECT 112.695 174.035 115.435 174.715 ;
        RECT 115.455 174.035 117.745 174.715 ;
        RECT 118.685 174.120 119.115 174.905 ;
        RECT 121.895 174.715 123.240 174.945 ;
        RECT 125.075 174.745 126.485 174.945 ;
        RECT 119.135 174.035 121.875 174.715 ;
        RECT 121.895 174.035 123.725 174.715 ;
        RECT 123.750 174.065 126.485 174.745 ;
        RECT 102.715 173.845 102.890 174.015 ;
        RECT 102.715 173.825 102.885 173.845 ;
        RECT 103.175 173.825 103.345 174.015 ;
        RECT 105.470 173.845 105.645 174.015 ;
        RECT 106.390 173.875 106.510 173.985 ;
        RECT 105.475 173.825 105.645 173.845 ;
        RECT 2.755 173.015 4.125 173.825 ;
        RECT 4.135 173.015 6.885 173.825 ;
        RECT 7.355 173.045 8.725 173.825 ;
        RECT 8.735 173.015 10.105 173.825 ;
        RECT 10.115 173.145 14.015 173.825 ;
        RECT 10.115 172.915 11.045 173.145 ;
        RECT 14.255 173.015 17.925 173.825 ;
        RECT 18.855 172.915 22.065 173.825 ;
        RECT 22.305 173.145 26.205 173.825 ;
        RECT 25.275 172.915 26.205 173.145 ;
        RECT 26.215 173.015 28.045 173.825 ;
        RECT 28.525 172.955 28.955 173.740 ;
        RECT 29.435 173.045 30.805 173.825 ;
        RECT 30.815 173.145 34.715 173.825 ;
        RECT 30.815 172.915 31.745 173.145 ;
        RECT 34.955 173.015 36.785 173.825 ;
        RECT 37.255 173.145 46.445 173.825 ;
        RECT 46.455 173.145 49.195 173.825 ;
        RECT 41.765 172.925 42.695 173.145 ;
        RECT 45.525 172.915 46.445 173.145 ;
        RECT 49.235 172.915 50.585 173.825 ;
        RECT 50.595 172.915 54.250 173.825 ;
        RECT 54.285 172.955 54.715 173.740 ;
        RECT 55.805 172.915 59.460 173.825 ;
        RECT 60.825 173.145 64.290 173.825 ;
        RECT 64.505 173.145 67.970 173.825 ;
        RECT 63.370 172.915 64.290 173.145 ;
        RECT 67.050 172.915 67.970 173.145 ;
        RECT 68.100 172.915 72.205 173.825 ;
        RECT 73.135 172.915 77.005 173.825 ;
        RECT 77.735 173.145 80.025 173.825 ;
        RECT 79.105 172.915 80.025 173.145 ;
        RECT 80.045 172.955 80.475 173.740 ;
        RECT 80.495 172.915 83.705 173.825 ;
        RECT 83.715 173.045 85.085 173.825 ;
        RECT 85.565 172.915 88.295 173.825 ;
        RECT 88.325 173.145 91.065 173.825 ;
        RECT 91.095 172.915 92.445 173.825 ;
        RECT 92.455 173.145 95.665 173.825 ;
        RECT 94.530 172.915 95.665 173.145 ;
        RECT 96.885 172.915 99.805 173.825 ;
        RECT 99.945 172.915 102.945 173.825 ;
        RECT 103.035 173.015 104.405 173.825 ;
        RECT 104.425 172.915 105.775 173.825 ;
        RECT 106.860 173.795 107.030 174.015 ;
        RECT 108.690 173.845 108.860 174.035 ;
        RECT 109.165 173.880 109.325 173.990 ;
        RECT 111.455 173.845 111.625 174.035 ;
        RECT 111.925 173.880 112.085 173.990 ;
        RECT 112.835 173.845 113.005 174.035 ;
        RECT 109.435 173.795 110.385 173.825 ;
        RECT 105.805 172.955 106.235 173.740 ;
        RECT 106.715 173.115 110.385 173.795 ;
        RECT 109.435 172.915 110.385 173.115 ;
        RECT 110.395 173.795 111.345 173.825 ;
        RECT 113.750 173.795 113.920 174.015 ;
        RECT 115.595 173.845 115.765 174.035 ;
        RECT 117.435 173.825 117.605 174.015 ;
        RECT 110.395 173.115 114.065 173.795 ;
        RECT 114.170 173.145 117.635 173.825 ;
        RECT 117.900 173.795 118.070 174.015 ;
        RECT 119.275 173.845 119.445 174.035 ;
        RECT 123.415 173.845 123.585 174.035 ;
        RECT 123.875 174.015 124.045 174.065 ;
        RECT 125.090 174.035 126.485 174.065 ;
        RECT 126.505 174.035 129.235 174.945 ;
        RECT 129.255 174.035 131.085 174.845 ;
        RECT 131.650 174.035 134.765 174.945 ;
        RECT 134.775 174.035 136.145 174.845 ;
        RECT 136.155 174.035 137.985 174.945 ;
        RECT 138.470 174.035 140.285 174.945 ;
        RECT 140.295 174.035 143.965 174.845 ;
        RECT 144.445 174.120 144.875 174.905 ;
        RECT 144.895 174.035 148.565 174.845 ;
        RECT 150.830 174.745 151.785 174.945 ;
        RECT 149.505 174.065 151.785 174.745 ;
        RECT 123.870 173.845 124.045 174.015 ;
        RECT 123.870 173.825 124.040 173.845 ;
        RECT 119.560 173.795 120.505 173.825 ;
        RECT 110.395 172.915 111.345 173.115 ;
        RECT 114.170 172.915 115.090 173.145 ;
        RECT 117.755 173.115 120.505 173.795 ;
        RECT 119.560 172.915 120.505 173.115 ;
        RECT 120.515 172.915 124.185 173.825 ;
        RECT 124.195 173.795 125.590 173.825 ;
        RECT 126.635 173.795 126.805 174.015 ;
        RECT 128.935 173.825 129.105 174.035 ;
        RECT 129.395 173.825 129.565 174.035 ;
        RECT 131.230 173.875 131.350 173.985 ;
        RECT 132.155 173.825 132.325 174.015 ;
        RECT 134.450 173.845 134.620 174.035 ;
        RECT 134.915 173.845 135.085 174.035 ;
        RECT 136.300 173.845 136.470 174.035 ;
        RECT 138.135 173.985 138.305 174.015 ;
        RECT 138.130 173.875 138.305 173.985 ;
        RECT 138.135 173.825 138.305 173.875 ;
        RECT 138.595 173.825 138.765 174.035 ;
        RECT 140.435 173.845 140.605 174.035 ;
        RECT 144.115 173.985 144.285 174.015 ;
        RECT 144.110 173.875 144.285 173.985 ;
        RECT 144.115 173.825 144.285 173.875 ;
        RECT 145.035 173.845 145.205 174.035 ;
        RECT 149.630 174.015 149.800 174.065 ;
        RECT 150.830 174.035 151.785 174.065 ;
        RECT 151.795 174.035 155.465 174.845 ;
        RECT 155.475 174.035 156.845 174.845 ;
        RECT 156.855 174.035 158.225 174.845 ;
        RECT 148.725 173.880 148.885 173.990 ;
        RECT 149.630 173.845 149.805 174.015 ;
        RECT 151.935 173.845 152.105 174.035 ;
        RECT 149.635 173.825 149.805 173.845 ;
        RECT 155.155 173.825 155.325 174.015 ;
        RECT 155.615 173.845 155.785 174.035 ;
        RECT 157.915 173.825 158.085 174.035 ;
        RECT 124.195 173.115 126.930 173.795 ;
        RECT 126.955 173.145 129.245 173.825 ;
        RECT 124.195 172.915 125.605 173.115 ;
        RECT 126.955 172.915 127.875 173.145 ;
        RECT 129.255 173.015 131.085 173.825 ;
        RECT 131.565 172.955 131.995 173.740 ;
        RECT 132.015 173.015 134.765 173.825 ;
        RECT 134.870 173.145 138.335 173.825 ;
        RECT 134.870 172.915 135.790 173.145 ;
        RECT 138.455 173.015 143.965 173.825 ;
        RECT 143.975 173.015 149.485 173.825 ;
        RECT 149.495 173.015 155.005 173.825 ;
        RECT 155.015 173.015 156.845 173.825 ;
        RECT 156.855 173.015 158.225 173.825 ;
      LAYER nwell ;
        RECT 2.560 169.795 158.420 172.625 ;
      LAYER pwell ;
        RECT 2.755 168.595 4.125 169.405 ;
        RECT 8.645 169.275 9.575 169.495 ;
        RECT 12.405 169.275 13.325 169.505 ;
        RECT 4.135 168.595 13.325 169.275 ;
        RECT 14.255 168.595 15.625 169.375 ;
        RECT 15.645 168.680 16.075 169.465 ;
        RECT 17.455 169.275 18.375 169.495 ;
        RECT 24.455 169.395 25.375 169.505 ;
        RECT 23.040 169.275 25.375 169.395 ;
        RECT 16.095 168.595 25.375 169.275 ;
        RECT 25.755 168.595 28.505 169.405 ;
        RECT 33.025 169.275 33.955 169.495 ;
        RECT 36.785 169.275 37.705 169.505 ;
        RECT 28.515 168.595 37.705 169.275 ;
        RECT 38.635 168.595 40.005 169.375 ;
        RECT 40.015 168.595 41.385 169.375 ;
        RECT 41.405 168.680 41.835 169.465 ;
        RECT 45.055 169.275 45.985 169.505 ;
        RECT 42.085 168.595 45.985 169.275 ;
        RECT 45.995 168.595 47.810 169.505 ;
        RECT 47.835 168.595 51.045 169.505 ;
        RECT 51.055 168.595 52.405 169.505 ;
        RECT 52.450 168.595 54.265 169.505 ;
        RECT 56.080 169.305 57.480 169.505 ;
        RECT 54.275 168.625 57.480 169.305 ;
        RECT 2.895 168.385 3.065 168.595 ;
        RECT 4.275 168.385 4.445 168.595 ;
        RECT 7.035 168.385 7.205 168.575 ;
        RECT 7.505 168.430 7.665 168.540 ;
        RECT 8.690 168.385 8.860 168.575 ;
        RECT 13.485 168.440 13.645 168.550 ;
        RECT 14.395 168.405 14.565 168.595 ;
        RECT 15.775 168.385 15.945 168.575 ;
        RECT 16.235 168.405 16.405 168.595 ;
        RECT 16.510 168.385 16.680 168.575 ;
        RECT 20.375 168.385 20.545 168.575 ;
        RECT 24.060 168.385 24.230 168.575 ;
        RECT 25.895 168.405 26.065 168.595 ;
        RECT 27.745 168.430 27.905 168.540 ;
        RECT 28.655 168.405 28.825 168.595 ;
        RECT 29.115 168.385 29.285 168.575 ;
        RECT 37.865 168.440 38.025 168.550 ;
        RECT 38.320 168.385 38.490 168.575 ;
        RECT 39.695 168.405 39.865 168.595 ;
        RECT 40.155 168.405 40.325 168.595 ;
        RECT 41.990 168.435 42.110 168.545 ;
        RECT 44.295 168.385 44.465 168.575 ;
        RECT 2.755 167.575 4.125 168.385 ;
        RECT 4.135 167.575 5.965 168.385 ;
        RECT 5.975 167.605 7.345 168.385 ;
        RECT 8.275 167.705 12.175 168.385 ;
        RECT 12.510 167.705 15.975 168.385 ;
        RECT 16.095 167.705 19.995 168.385 ;
        RECT 8.275 167.475 9.205 167.705 ;
        RECT 12.510 167.475 13.430 167.705 ;
        RECT 16.095 167.475 17.025 167.705 ;
        RECT 20.235 167.575 23.905 168.385 ;
        RECT 23.915 167.475 27.570 168.385 ;
        RECT 28.525 167.515 28.955 168.300 ;
        RECT 28.975 167.705 38.165 168.385 ;
        RECT 33.485 167.485 34.415 167.705 ;
        RECT 37.245 167.475 38.165 167.705 ;
        RECT 38.175 167.475 41.830 168.385 ;
        RECT 42.315 167.705 44.605 168.385 ;
        RECT 44.760 168.355 44.930 168.575 ;
        RECT 45.400 168.405 45.570 168.595 ;
        RECT 47.515 168.405 47.685 168.595 ;
        RECT 49.815 168.405 49.985 168.575 ;
        RECT 49.815 168.385 49.965 168.405 ;
        RECT 50.280 168.385 50.450 168.575 ;
        RECT 50.745 168.405 50.915 168.595 ;
        RECT 51.200 168.405 51.370 168.595 ;
        RECT 52.575 168.405 52.745 168.595 ;
        RECT 53.950 168.435 54.070 168.545 ;
        RECT 54.420 168.405 54.590 168.625 ;
        RECT 56.080 168.595 57.480 168.625 ;
        RECT 57.645 168.595 61.300 169.505 ;
        RECT 61.635 168.595 63.005 169.405 ;
        RECT 63.165 168.595 66.820 169.505 ;
        RECT 67.165 168.680 67.595 169.465 ;
        RECT 72.125 169.275 73.055 169.495 ;
        RECT 75.885 169.275 77.225 169.505 ;
        RECT 67.615 168.595 77.225 169.275 ;
        RECT 77.275 169.275 78.410 169.505 ;
        RECT 80.695 169.415 81.645 169.505 ;
        RECT 77.275 168.595 80.485 169.275 ;
        RECT 80.695 168.595 82.625 169.415 ;
        RECT 83.280 169.275 84.625 169.505 ;
        RECT 87.175 169.275 88.765 169.505 ;
        RECT 82.795 168.595 84.625 169.275 ;
        RECT 85.095 168.595 88.765 169.275 ;
        RECT 88.795 168.595 90.145 169.505 ;
        RECT 91.075 169.275 92.420 169.505 ;
        RECT 91.075 168.595 92.905 169.275 ;
        RECT 92.925 168.680 93.355 169.465 ;
        RECT 93.375 168.595 99.565 169.505 ;
        RECT 99.815 168.595 103.025 169.505 ;
        RECT 103.165 168.595 106.165 169.505 ;
        RECT 106.715 168.595 116.685 169.505 ;
        RECT 116.835 168.595 118.665 169.405 ;
        RECT 118.685 168.680 119.115 169.465 ;
        RECT 126.015 169.275 126.935 169.495 ;
        RECT 133.015 169.395 133.935 169.505 ;
        RECT 131.600 169.275 133.935 169.395 ;
        RECT 138.825 169.275 139.755 169.495 ;
        RECT 142.585 169.275 143.925 169.505 ;
        RECT 119.145 168.595 121.885 169.275 ;
        RECT 121.895 168.595 124.635 169.275 ;
        RECT 124.655 168.595 133.935 169.275 ;
        RECT 134.315 168.595 143.925 169.275 ;
        RECT 144.445 168.680 144.875 169.465 ;
        RECT 144.895 168.595 150.405 169.405 ;
        RECT 150.415 168.595 155.925 169.405 ;
        RECT 156.855 168.595 158.225 169.405 ;
        RECT 57.645 168.575 57.805 168.595 ;
        RECT 57.635 168.385 57.805 168.575 ;
        RECT 58.090 168.435 58.210 168.545 ;
        RECT 58.555 168.385 58.725 168.575 ;
        RECT 59.935 168.385 60.105 168.575 ;
        RECT 61.775 168.405 61.945 168.595 ;
        RECT 63.165 168.575 63.325 168.595 ;
        RECT 63.155 168.405 63.325 168.575 ;
        RECT 67.755 168.405 67.925 168.595 ;
        RECT 69.130 168.435 69.250 168.545 ;
        RECT 71.435 168.385 71.605 168.575 ;
        RECT 75.300 168.385 75.470 168.575 ;
        RECT 78.795 168.385 78.965 168.575 ;
        RECT 79.265 168.430 79.425 168.540 ;
        RECT 80.175 168.405 80.345 168.595 ;
        RECT 82.475 168.575 82.625 168.595 ;
        RECT 82.475 168.405 82.645 168.575 ;
        RECT 82.935 168.405 83.105 168.595 ;
        RECT 84.315 168.405 84.485 168.575 ;
        RECT 84.775 168.545 84.945 168.575 ;
        RECT 84.770 168.435 84.945 168.545 ;
        RECT 84.775 168.405 84.945 168.435 ;
        RECT 85.240 168.405 85.410 168.595 ;
        RECT 87.085 168.430 87.245 168.540 ;
        RECT 88.910 168.405 89.080 168.595 ;
        RECT 90.305 168.440 90.465 168.550 ;
        RECT 84.315 168.385 84.475 168.405 ;
        RECT 46.890 168.355 47.825 168.385 ;
        RECT 44.760 168.155 47.825 168.355 ;
        RECT 42.315 167.475 43.235 167.705 ;
        RECT 44.615 167.675 47.825 168.155 ;
        RECT 44.615 167.475 45.545 167.675 ;
        RECT 46.875 167.475 47.825 167.675 ;
        RECT 48.035 167.565 49.965 168.385 ;
        RECT 48.035 167.475 48.985 167.565 ;
        RECT 50.135 167.475 53.790 168.385 ;
        RECT 54.285 167.515 54.715 168.300 ;
        RECT 54.735 167.705 57.945 168.385 ;
        RECT 54.735 167.475 55.870 167.705 ;
        RECT 58.415 167.605 59.785 168.385 ;
        RECT 59.795 167.705 68.985 168.385 ;
        RECT 64.305 167.485 65.235 167.705 ;
        RECT 68.065 167.475 68.985 167.705 ;
        RECT 69.455 167.705 71.745 168.385 ;
        RECT 71.985 167.705 75.885 168.385 ;
        RECT 69.455 167.475 70.375 167.705 ;
        RECT 74.955 167.475 75.885 167.705 ;
        RECT 75.895 167.475 79.065 168.385 ;
        RECT 80.045 167.515 80.475 168.300 ;
        RECT 80.820 167.475 84.475 168.385 ;
        RECT 84.780 168.385 84.945 168.405 ;
        RECT 90.750 168.385 90.920 168.575 ;
        RECT 91.220 168.385 91.390 168.575 ;
        RECT 92.595 168.405 92.765 168.595 ;
        RECT 93.520 168.405 93.690 168.595 ;
        RECT 94.430 168.435 94.550 168.545 ;
        RECT 98.115 168.385 98.285 168.575 ;
        RECT 100.415 168.405 100.585 168.575 ;
        RECT 100.885 168.430 101.045 168.540 ;
        RECT 100.415 168.385 100.580 168.405 ;
        RECT 101.795 168.385 101.965 168.575 ;
        RECT 102.710 168.405 102.880 168.595 ;
        RECT 105.935 168.405 106.105 168.595 ;
        RECT 106.390 168.435 106.510 168.545 ;
        RECT 106.860 168.405 107.030 168.595 ;
        RECT 107.315 168.385 107.485 168.575 ;
        RECT 107.775 168.385 107.945 168.575 ;
        RECT 116.975 168.405 117.145 168.595 ;
        RECT 121.575 168.405 121.745 168.595 ;
        RECT 122.035 168.405 122.205 168.595 ;
        RECT 124.795 168.405 124.965 168.595 ;
        RECT 127.095 168.385 127.265 168.575 ;
        RECT 127.555 168.385 127.725 168.575 ;
        RECT 131.230 168.435 131.350 168.545 ;
        RECT 132.165 168.430 132.325 168.540 ;
        RECT 134.455 168.405 134.625 168.595 ;
        RECT 136.750 168.385 136.920 168.575 ;
        RECT 137.220 168.385 137.390 168.575 ;
        RECT 142.270 168.385 142.440 168.575 ;
        RECT 142.735 168.385 142.905 168.575 ;
        RECT 144.110 168.435 144.230 168.545 ;
        RECT 144.575 168.385 144.745 168.575 ;
        RECT 145.035 168.405 145.205 168.595 ;
        RECT 149.635 168.385 149.805 168.575 ;
        RECT 150.095 168.385 150.265 168.575 ;
        RECT 150.555 168.405 150.725 168.595 ;
        RECT 151.935 168.385 152.105 168.575 ;
        RECT 155.615 168.385 155.785 168.575 ;
        RECT 156.085 168.440 156.245 168.550 ;
        RECT 157.915 168.385 158.085 168.595 ;
        RECT 84.780 167.705 86.615 168.385 ;
        RECT 85.685 167.475 86.615 167.705 ;
        RECT 88.145 167.475 91.065 168.385 ;
        RECT 91.075 167.475 93.995 168.385 ;
        RECT 94.850 167.705 98.315 168.385 ;
        RECT 98.745 167.705 100.580 168.385 ;
        RECT 94.850 167.475 95.770 167.705 ;
        RECT 98.745 167.475 99.675 167.705 ;
        RECT 101.655 167.475 105.715 168.385 ;
        RECT 105.805 167.515 106.235 168.300 ;
        RECT 106.265 167.475 107.615 168.385 ;
        RECT 107.635 167.705 116.740 168.385 ;
        RECT 117.035 167.705 127.405 168.385 ;
        RECT 117.035 167.475 119.245 167.705 ;
        RECT 121.965 167.485 122.895 167.705 ;
        RECT 127.415 167.575 131.085 168.385 ;
        RECT 131.565 167.515 131.995 168.300 ;
        RECT 133.175 167.475 137.065 168.385 ;
        RECT 137.075 167.475 139.685 168.385 ;
        RECT 139.975 167.475 142.585 168.385 ;
        RECT 142.595 167.575 144.425 168.385 ;
        RECT 144.545 167.705 148.010 168.385 ;
        RECT 147.090 167.475 148.010 167.705 ;
        RECT 148.115 167.705 149.945 168.385 ;
        RECT 149.955 167.705 151.785 168.385 ;
        RECT 148.115 167.475 149.460 167.705 ;
        RECT 150.440 167.475 151.785 167.705 ;
        RECT 151.795 167.575 155.465 168.385 ;
        RECT 155.475 167.575 156.845 168.385 ;
        RECT 156.855 167.575 158.225 168.385 ;
      LAYER nwell ;
        RECT 2.560 164.355 158.420 167.185 ;
      LAYER pwell ;
        RECT 2.755 163.155 4.125 163.965 ;
        RECT 5.495 163.835 6.415 164.055 ;
        RECT 12.495 163.955 13.415 164.065 ;
        RECT 11.080 163.835 13.415 163.955 ;
        RECT 4.135 163.155 13.415 163.835 ;
        RECT 13.795 163.155 15.165 163.935 ;
        RECT 15.645 163.240 16.075 164.025 ;
        RECT 16.095 163.835 17.025 164.065 ;
        RECT 16.095 163.155 19.995 163.835 ;
        RECT 20.235 163.155 22.065 163.965 ;
        RECT 22.075 163.155 25.730 164.065 ;
        RECT 26.675 163.155 28.045 163.935 ;
        RECT 28.055 163.835 28.985 164.065 ;
        RECT 28.055 163.155 31.955 163.835 ;
        RECT 32.280 163.155 41.385 163.835 ;
        RECT 41.405 163.240 41.835 164.025 ;
        RECT 41.855 163.155 45.510 164.065 ;
        RECT 48.755 163.835 49.685 164.065 ;
        RECT 57.405 163.835 58.335 164.055 ;
        RECT 61.165 163.835 62.085 164.065 ;
        RECT 65.295 163.835 66.225 164.065 ;
        RECT 46.005 163.155 48.745 163.835 ;
        RECT 48.755 163.155 52.655 163.835 ;
        RECT 52.895 163.155 62.085 163.835 ;
        RECT 62.325 163.155 66.225 163.835 ;
        RECT 67.165 163.240 67.595 164.025 ;
        RECT 67.615 163.155 76.720 163.835 ;
        RECT 76.815 163.155 78.645 163.965 ;
        RECT 81.855 163.835 82.785 164.065 ;
        RECT 85.555 163.835 86.900 164.065 ;
        RECT 78.885 163.155 82.785 163.835 ;
        RECT 82.795 163.155 85.535 163.835 ;
        RECT 85.555 163.155 87.385 163.835 ;
        RECT 88.325 163.155 89.675 164.065 ;
        RECT 90.165 163.155 91.515 164.065 ;
        RECT 91.555 163.155 92.905 164.065 ;
        RECT 92.925 163.240 93.355 164.025 ;
        RECT 93.575 163.835 95.785 164.065 ;
        RECT 98.505 163.835 99.435 164.055 ;
        RECT 104.510 163.835 105.430 164.065 ;
        RECT 108.295 163.835 110.505 164.065 ;
        RECT 113.225 163.835 114.155 164.055 ;
        RECT 93.575 163.155 103.945 163.835 ;
        RECT 104.510 163.155 107.975 163.835 ;
        RECT 108.295 163.155 118.665 163.835 ;
        RECT 118.685 163.240 119.115 164.025 ;
        RECT 122.395 163.835 123.735 164.065 ;
        RECT 126.565 163.835 127.495 164.055 ;
        RECT 132.055 163.835 133.395 164.065 ;
        RECT 136.225 163.835 137.155 164.055 ;
        RECT 119.135 163.155 121.875 163.835 ;
        RECT 122.395 163.155 132.005 163.835 ;
        RECT 132.055 163.155 141.665 163.835 ;
        RECT 141.675 163.155 144.425 163.965 ;
        RECT 144.445 163.240 144.875 164.025 ;
        RECT 147.655 163.835 149.000 164.065 ;
        RECT 144.905 163.155 147.645 163.835 ;
        RECT 147.655 163.155 149.485 163.835 ;
        RECT 149.495 163.155 155.005 163.965 ;
        RECT 155.015 163.155 156.845 163.965 ;
        RECT 156.855 163.155 158.225 163.965 ;
        RECT 2.895 162.945 3.065 163.155 ;
        RECT 4.275 162.965 4.445 163.155 ;
        RECT 6.115 162.945 6.285 163.135 ;
        RECT 6.850 162.945 7.020 163.135 ;
        RECT 10.715 162.945 10.885 163.135 ;
        RECT 14.855 162.965 15.025 163.155 ;
        RECT 15.310 162.995 15.430 163.105 ;
        RECT 16.510 162.965 16.680 163.155 ;
        RECT 20.375 162.965 20.545 163.155 ;
        RECT 22.220 162.965 22.390 163.155 ;
        RECT 23.135 162.945 23.305 163.135 ;
        RECT 23.595 162.945 23.765 163.135 ;
        RECT 25.905 163.000 26.065 163.110 ;
        RECT 26.815 162.945 26.985 163.155 ;
        RECT 28.470 162.965 28.640 163.155 ;
        RECT 29.125 162.990 29.285 163.100 ;
        RECT 31.875 162.965 32.045 163.135 ;
        RECT 31.875 162.945 32.025 162.965 ;
        RECT 41.075 162.945 41.245 163.155 ;
        RECT 42.000 162.965 42.170 163.155 ;
        RECT 45.670 162.995 45.790 163.105 ;
        RECT 48.435 162.965 48.605 163.155 ;
        RECT 49.170 162.965 49.340 163.155 ;
        RECT 50.275 162.945 50.445 163.135 ;
        RECT 50.730 162.995 50.850 163.105 ;
        RECT 51.200 162.945 51.370 163.135 ;
        RECT 53.035 162.965 53.205 163.155 ;
        RECT 54.880 162.945 55.050 163.135 ;
        RECT 59.015 162.945 59.185 163.135 ;
        RECT 59.470 162.995 59.590 163.105 ;
        RECT 63.610 162.945 63.780 163.135 ;
        RECT 64.075 162.945 64.245 163.135 ;
        RECT 65.640 162.965 65.810 163.155 ;
        RECT 66.385 163.000 66.545 163.110 ;
        RECT 67.755 162.965 67.925 163.155 ;
        RECT 76.680 162.945 76.850 163.135 ;
        RECT 76.955 162.965 77.125 163.155 ;
        RECT 79.715 162.945 79.885 163.135 ;
        RECT 82.200 162.965 82.370 163.155 ;
        RECT 82.935 162.965 83.105 163.155 ;
        RECT 84.040 162.945 84.210 163.135 ;
        RECT 84.785 162.990 84.945 163.100 ;
        RECT 87.075 162.965 87.245 163.155 ;
        RECT 87.545 163.000 87.705 163.110 ;
        RECT 88.455 162.945 88.625 163.135 ;
        RECT 89.375 162.965 89.545 163.155 ;
        RECT 89.830 162.995 89.950 163.105 ;
        RECT 90.295 162.965 90.465 163.155 ;
        RECT 90.750 162.945 90.920 163.135 ;
        RECT 92.140 162.945 92.310 163.135 ;
        RECT 92.590 163.100 92.760 163.155 ;
        RECT 92.590 162.990 92.765 163.100 ;
        RECT 92.590 162.965 92.760 162.990 ;
        RECT 93.515 162.945 93.685 163.135 ;
        RECT 98.575 162.945 98.745 163.135 ;
        RECT 99.035 162.945 99.205 163.135 ;
        RECT 103.635 162.965 103.805 163.155 ;
        RECT 104.090 162.995 104.210 163.105 ;
        RECT 105.200 162.945 105.370 163.135 ;
        RECT 107.775 162.965 107.945 163.155 ;
        RECT 116.515 162.945 116.685 163.135 ;
        RECT 118.355 162.965 118.525 163.155 ;
        RECT 119.275 162.965 119.445 163.155 ;
        RECT 120.380 162.945 120.550 163.135 ;
        RECT 122.035 163.105 122.205 163.135 ;
        RECT 122.030 162.995 122.205 163.105 ;
        RECT 122.035 162.945 122.205 162.995 ;
        RECT 122.500 162.945 122.670 163.135 ;
        RECT 123.870 162.995 123.990 163.105 ;
        RECT 127.740 162.945 127.910 163.135 ;
        RECT 129.395 162.945 129.565 163.135 ;
        RECT 129.855 162.945 130.025 163.135 ;
        RECT 131.230 162.995 131.350 163.105 ;
        RECT 131.695 162.965 131.865 163.155 ;
        RECT 135.560 162.945 135.730 163.135 ;
        RECT 136.295 162.945 136.465 163.135 ;
        RECT 141.355 162.965 141.525 163.155 ;
        RECT 141.815 162.965 141.985 163.155 ;
        RECT 146.875 162.945 147.045 163.135 ;
        RECT 147.335 162.945 147.505 163.155 ;
        RECT 149.175 162.965 149.345 163.155 ;
        RECT 149.635 162.965 149.805 163.155 ;
        RECT 152.855 162.945 153.025 163.135 ;
        RECT 155.155 162.965 155.325 163.155 ;
        RECT 156.530 162.995 156.650 163.105 ;
        RECT 157.915 162.945 158.085 163.155 ;
        RECT 2.755 162.135 4.125 162.945 ;
        RECT 5.055 162.165 6.425 162.945 ;
        RECT 6.435 162.265 10.335 162.945 ;
        RECT 10.575 162.265 19.765 162.945 ;
        RECT 6.435 162.035 7.365 162.265 ;
        RECT 15.085 162.045 16.015 162.265 ;
        RECT 18.845 162.035 19.765 162.265 ;
        RECT 19.870 162.265 23.335 162.945 ;
        RECT 19.870 162.035 20.790 162.265 ;
        RECT 23.455 162.035 26.665 162.945 ;
        RECT 26.675 162.135 28.505 162.945 ;
        RECT 28.525 162.075 28.955 162.860 ;
        RECT 30.095 162.125 32.025 162.945 ;
        RECT 32.280 162.265 41.385 162.945 ;
        RECT 41.395 162.265 50.585 162.945 ;
        RECT 30.095 162.035 31.045 162.125 ;
        RECT 41.395 162.035 42.315 162.265 ;
        RECT 45.145 162.045 46.075 162.265 ;
        RECT 51.055 162.035 53.975 162.945 ;
        RECT 54.285 162.075 54.715 162.860 ;
        RECT 54.735 162.035 57.655 162.945 ;
        RECT 57.955 162.165 59.325 162.945 ;
        RECT 59.795 162.265 63.925 162.945 ;
        RECT 63.935 162.265 73.125 162.945 ;
        RECT 73.365 162.265 77.265 162.945 ;
        RECT 77.285 162.265 80.025 162.945 ;
        RECT 62.585 162.035 63.925 162.265 ;
        RECT 68.445 162.045 69.375 162.265 ;
        RECT 72.205 162.035 73.125 162.265 ;
        RECT 76.335 162.035 77.265 162.265 ;
        RECT 80.045 162.075 80.475 162.860 ;
        RECT 80.725 162.265 84.625 162.945 ;
        RECT 83.695 162.035 84.625 162.265 ;
        RECT 85.555 162.265 88.765 162.945 ;
        RECT 85.555 162.035 86.690 162.265 ;
        RECT 88.875 162.035 91.065 162.945 ;
        RECT 91.075 162.035 92.425 162.945 ;
        RECT 93.375 162.265 95.205 162.945 ;
        RECT 93.860 162.035 95.205 162.265 ;
        RECT 95.310 162.265 98.775 162.945 ;
        RECT 98.895 162.265 101.635 162.945 ;
        RECT 101.885 162.265 105.785 162.945 ;
        RECT 95.310 162.035 96.230 162.265 ;
        RECT 104.855 162.035 105.785 162.265 ;
        RECT 105.805 162.075 106.235 162.860 ;
        RECT 106.455 162.265 116.825 162.945 ;
        RECT 117.065 162.265 120.965 162.945 ;
        RECT 106.455 162.035 108.665 162.265 ;
        RECT 111.385 162.045 112.315 162.265 ;
        RECT 120.035 162.035 120.965 162.265 ;
        RECT 120.975 162.165 122.345 162.945 ;
        RECT 122.355 162.035 123.705 162.945 ;
        RECT 124.425 162.265 128.325 162.945 ;
        RECT 127.395 162.035 128.325 162.265 ;
        RECT 128.335 162.165 129.705 162.945 ;
        RECT 129.715 162.165 131.085 162.945 ;
        RECT 131.565 162.075 131.995 162.860 ;
        RECT 132.245 162.265 136.145 162.945 ;
        RECT 135.215 162.035 136.145 162.265 ;
        RECT 136.155 162.165 137.525 162.945 ;
        RECT 137.575 162.265 147.185 162.945 ;
        RECT 137.575 162.035 138.915 162.265 ;
        RECT 141.745 162.045 142.675 162.265 ;
        RECT 147.195 162.135 152.705 162.945 ;
        RECT 152.715 162.135 156.385 162.945 ;
        RECT 156.855 162.135 158.225 162.945 ;
      LAYER nwell ;
        RECT 2.560 158.915 158.420 161.745 ;
      LAYER pwell ;
        RECT 2.755 157.715 4.125 158.525 ;
        RECT 8.645 158.395 9.575 158.615 ;
        RECT 12.405 158.395 13.325 158.625 ;
        RECT 4.135 157.715 13.325 158.395 ;
        RECT 13.335 157.715 14.705 158.495 ;
        RECT 15.645 157.800 16.075 158.585 ;
        RECT 16.095 158.395 17.025 158.625 ;
        RECT 16.095 157.715 19.995 158.395 ;
        RECT 20.235 157.715 22.065 158.525 ;
        RECT 22.535 157.715 26.190 158.625 ;
        RECT 26.215 157.715 28.965 158.525 ;
        RECT 32.175 158.395 33.105 158.625 ;
        RECT 29.205 157.715 33.105 158.395 ;
        RECT 34.035 157.715 37.690 158.625 ;
        RECT 37.715 157.715 41.370 158.625 ;
        RECT 41.405 157.800 41.835 158.585 ;
        RECT 41.855 158.395 42.785 158.625 ;
        RECT 46.305 158.395 47.235 158.625 ;
        RECT 51.495 158.395 52.425 158.625 ;
        RECT 41.855 157.715 45.755 158.395 ;
        RECT 46.305 157.715 48.140 158.395 ;
        RECT 48.525 157.715 52.425 158.395 ;
        RECT 52.435 158.395 53.355 158.625 ;
        RECT 56.185 158.395 57.115 158.615 ;
        RECT 52.435 157.715 61.625 158.395 ;
        RECT 61.635 157.715 63.005 158.495 ;
        RECT 63.015 158.395 63.945 158.625 ;
        RECT 63.015 157.715 66.915 158.395 ;
        RECT 67.165 157.800 67.595 158.585 ;
        RECT 72.585 158.395 73.515 158.615 ;
        RECT 76.345 158.395 77.265 158.625 ;
        RECT 68.075 157.715 77.265 158.395 ;
        RECT 77.275 158.395 78.615 158.625 ;
        RECT 83.235 158.395 84.165 158.625 ;
        RECT 85.995 158.395 86.925 158.625 ;
        RECT 77.275 157.715 81.405 158.395 ;
        RECT 81.415 157.715 84.165 158.395 ;
        RECT 84.175 157.715 86.925 158.395 ;
        RECT 86.935 157.715 88.305 158.495 ;
        RECT 88.800 158.425 90.155 158.625 ;
        RECT 88.800 158.395 91.480 158.425 ;
        RECT 88.315 157.745 91.480 158.395 ;
        RECT 88.315 157.715 90.155 157.745 ;
        RECT 91.535 157.715 92.905 158.525 ;
        RECT 92.925 157.800 93.355 158.585 ;
        RECT 93.385 157.715 96.115 158.625 ;
        RECT 101.565 158.395 102.495 158.615 ;
        RECT 105.325 158.395 106.245 158.625 ;
        RECT 108.060 158.425 109.005 158.625 ;
        RECT 97.055 157.715 106.245 158.395 ;
        RECT 106.255 157.745 109.005 158.425 ;
        RECT 2.895 157.505 3.065 157.715 ;
        RECT 4.275 157.505 4.445 157.715 ;
        RECT 6.110 157.555 6.230 157.665 ;
        RECT 9.980 157.505 10.150 157.695 ;
        RECT 10.715 157.505 10.885 157.695 ;
        RECT 14.395 157.525 14.565 157.715 ;
        RECT 14.865 157.560 15.025 157.670 ;
        RECT 16.510 157.525 16.680 157.715 ;
        RECT 20.375 157.525 20.545 157.715 ;
        RECT 22.210 157.555 22.330 157.665 ;
        RECT 22.680 157.525 22.850 157.715 ;
        RECT 23.135 157.505 23.305 157.695 ;
        RECT 26.355 157.505 26.525 157.715 ;
        RECT 27.735 157.505 27.905 157.695 ;
        RECT 28.190 157.555 28.310 157.665 ;
        RECT 29.390 157.505 29.560 157.695 ;
        RECT 32.520 157.525 32.690 157.715 ;
        RECT 33.265 157.550 33.425 157.670 ;
        RECT 34.180 157.505 34.350 157.715 ;
        RECT 37.860 157.505 38.030 157.715 ;
        RECT 41.070 157.555 41.190 157.665 ;
        RECT 41.535 157.505 41.705 157.695 ;
        RECT 42.270 157.525 42.440 157.715 ;
        RECT 47.975 157.695 48.140 157.715 ;
        RECT 2.755 156.695 4.125 157.505 ;
        RECT 4.135 156.695 5.965 157.505 ;
        RECT 6.665 156.825 10.565 157.505 ;
        RECT 10.575 156.825 19.765 157.505 ;
        RECT 9.635 156.595 10.565 156.825 ;
        RECT 15.085 156.605 16.015 156.825 ;
        RECT 18.845 156.595 19.765 156.825 ;
        RECT 19.870 156.825 23.335 157.505 ;
        RECT 19.870 156.595 20.790 156.825 ;
        RECT 23.455 156.595 26.665 157.505 ;
        RECT 26.675 156.725 28.045 157.505 ;
        RECT 28.525 156.635 28.955 157.420 ;
        RECT 28.975 156.825 32.875 157.505 ;
        RECT 28.975 156.595 29.905 156.825 ;
        RECT 34.035 156.595 37.690 157.505 ;
        RECT 37.720 157.275 39.925 157.505 ;
        RECT 37.720 156.595 40.865 157.275 ;
        RECT 41.395 156.825 44.135 157.505 ;
        RECT 44.295 157.475 44.465 157.695 ;
        RECT 47.975 157.525 48.145 157.695 ;
        RECT 46.455 157.475 47.825 157.505 ;
        RECT 44.155 156.795 47.825 157.475 ;
        RECT 46.440 156.595 47.825 156.795 ;
        RECT 47.835 157.475 48.780 157.505 ;
        RECT 50.735 157.475 50.905 157.695 ;
        RECT 51.840 157.525 52.010 157.715 ;
        RECT 47.835 157.275 50.905 157.475 ;
        RECT 51.055 157.475 52.450 157.505 ;
        RECT 53.495 157.475 53.665 157.695 ;
        RECT 53.950 157.555 54.070 157.665 ;
        RECT 54.735 157.475 56.130 157.505 ;
        RECT 57.175 157.475 57.345 157.695 ;
        RECT 57.630 157.555 57.750 157.665 ;
        RECT 58.095 157.505 58.265 157.695 ;
        RECT 60.865 157.550 61.025 157.660 ;
        RECT 61.315 157.525 61.485 157.715 ;
        RECT 61.775 157.525 61.945 157.715 ;
        RECT 62.050 157.505 62.220 157.695 ;
        RECT 63.430 157.525 63.600 157.715 ;
        RECT 65.915 157.505 66.085 157.695 ;
        RECT 67.750 157.555 67.870 157.665 ;
        RECT 68.215 157.525 68.385 157.715 ;
        RECT 75.125 157.550 75.285 157.660 ;
        RECT 76.040 157.505 76.210 157.695 ;
        RECT 77.420 157.525 77.590 157.715 ;
        RECT 80.630 157.555 80.750 157.665 ;
        RECT 81.095 157.505 81.265 157.695 ;
        RECT 81.555 157.525 81.725 157.715 ;
        RECT 84.315 157.525 84.485 157.715 ;
        RECT 87.075 157.525 87.245 157.715 ;
        RECT 88.455 157.525 88.625 157.715 ;
        RECT 91.675 157.505 91.845 157.715 ;
        RECT 92.135 157.505 92.305 157.695 ;
        RECT 93.515 157.525 93.685 157.715 ;
        RECT 94.905 157.550 95.065 157.660 ;
        RECT 96.285 157.560 96.445 157.670 ;
        RECT 97.195 157.525 97.365 157.715 ;
        RECT 99.220 157.505 99.390 157.695 ;
        RECT 100.875 157.505 101.045 157.695 ;
        RECT 101.330 157.555 101.450 157.665 ;
        RECT 101.795 157.505 101.965 157.695 ;
        RECT 105.475 157.505 105.645 157.695 ;
        RECT 106.400 157.525 106.570 157.745 ;
        RECT 108.060 157.715 109.005 157.745 ;
        RECT 109.475 157.715 118.580 158.395 ;
        RECT 118.685 157.800 119.115 158.585 ;
        RECT 119.135 158.395 120.065 158.625 ;
        RECT 119.135 157.715 123.035 158.395 ;
        RECT 123.275 157.715 125.885 158.625 ;
        RECT 127.085 158.395 128.015 158.625 ;
        RECT 126.180 157.715 128.015 158.395 ;
        RECT 128.345 157.715 129.695 158.625 ;
        RECT 129.715 157.715 131.085 158.495 ;
        RECT 132.015 158.395 132.945 158.625 ;
        RECT 137.075 158.395 138.005 158.625 ;
        RECT 132.015 157.715 135.915 158.395 ;
        RECT 137.075 157.715 140.975 158.395 ;
        RECT 141.215 157.715 143.965 158.525 ;
        RECT 144.445 157.800 144.875 158.585 ;
        RECT 144.895 157.715 150.405 158.525 ;
        RECT 150.415 157.715 155.925 158.525 ;
        RECT 156.855 157.715 158.225 158.525 ;
        RECT 106.670 157.505 106.840 157.695 ;
        RECT 109.150 157.555 109.270 157.665 ;
        RECT 109.615 157.525 109.785 157.715 ;
        RECT 110.530 157.555 110.650 157.665 ;
        RECT 111.000 157.505 111.170 157.695 ;
        RECT 114.215 157.505 114.385 157.695 ;
        RECT 119.550 157.525 119.720 157.715 ;
        RECT 123.420 157.525 123.590 157.715 ;
        RECT 126.180 157.695 126.345 157.715 ;
        RECT 123.870 157.555 123.990 157.665 ;
        RECT 125.255 157.505 125.425 157.695 ;
        RECT 125.990 157.505 126.160 157.695 ;
        RECT 126.175 157.525 126.345 157.695 ;
        RECT 128.475 157.525 128.645 157.715 ;
        RECT 129.850 157.555 129.970 157.665 ;
        RECT 130.315 157.505 130.485 157.695 ;
        RECT 130.775 157.525 130.945 157.715 ;
        RECT 131.245 157.560 131.405 157.670 ;
        RECT 132.430 157.525 132.600 157.715 ;
        RECT 136.305 157.560 136.465 157.670 ;
        RECT 137.490 157.525 137.660 157.715 ;
        RECT 141.355 157.505 141.525 157.715 ;
        RECT 141.815 157.505 141.985 157.695 ;
        RECT 144.110 157.555 144.230 157.665 ;
        RECT 145.035 157.525 145.205 157.715 ;
        RECT 150.555 157.525 150.725 157.715 ;
        RECT 151.475 157.505 151.645 157.695 ;
        RECT 156.085 157.560 156.245 157.670 ;
        RECT 157.915 157.505 158.085 157.715 ;
        RECT 47.835 156.795 51.045 157.275 ;
        RECT 47.835 156.595 48.780 156.795 ;
        RECT 50.115 156.595 51.045 156.795 ;
        RECT 51.055 156.795 53.790 157.475 ;
        RECT 51.055 156.595 52.465 156.795 ;
        RECT 54.285 156.635 54.715 157.420 ;
        RECT 54.735 156.795 57.470 157.475 ;
        RECT 57.955 156.825 60.695 157.505 ;
        RECT 61.635 156.825 65.535 157.505 ;
        RECT 65.775 156.825 74.965 157.505 ;
        RECT 54.735 156.595 56.145 156.795 ;
        RECT 61.635 156.595 62.565 156.825 ;
        RECT 70.285 156.605 71.215 156.825 ;
        RECT 74.045 156.595 74.965 156.825 ;
        RECT 75.895 156.825 80.025 157.505 ;
        RECT 75.895 156.595 77.235 156.825 ;
        RECT 80.045 156.635 80.475 157.420 ;
        RECT 80.955 156.825 82.785 157.505 ;
        RECT 81.440 156.595 82.785 156.825 ;
        RECT 82.795 156.825 91.985 157.505 ;
        RECT 91.995 156.825 94.735 157.505 ;
        RECT 95.905 156.825 99.805 157.505 ;
        RECT 82.795 156.595 83.715 156.825 ;
        RECT 86.545 156.605 87.475 156.825 ;
        RECT 98.875 156.595 99.805 156.825 ;
        RECT 99.815 156.725 101.185 157.505 ;
        RECT 101.655 156.725 103.025 157.505 ;
        RECT 103.045 156.825 105.785 157.505 ;
        RECT 105.805 156.635 106.235 157.420 ;
        RECT 106.255 156.825 110.155 157.505 ;
        RECT 110.860 157.275 113.065 157.505 ;
        RECT 106.255 156.595 107.185 156.825 ;
        RECT 110.860 156.595 114.005 157.275 ;
        RECT 114.075 156.825 123.685 157.505 ;
        RECT 118.585 156.605 119.515 156.825 ;
        RECT 122.345 156.595 123.685 156.825 ;
        RECT 124.195 156.725 125.565 157.505 ;
        RECT 125.575 156.825 129.475 157.505 ;
        RECT 125.575 156.595 126.505 156.825 ;
        RECT 130.175 156.725 131.545 157.505 ;
        RECT 131.565 156.635 131.995 157.420 ;
        RECT 132.055 156.825 141.665 157.505 ;
        RECT 141.675 156.825 151.285 157.505 ;
        RECT 132.055 156.595 133.395 156.825 ;
        RECT 136.225 156.605 137.155 156.825 ;
        RECT 146.185 156.605 147.115 156.825 ;
        RECT 149.945 156.595 151.285 156.825 ;
        RECT 151.335 156.695 156.845 157.505 ;
        RECT 156.855 156.695 158.225 157.505 ;
      LAYER nwell ;
        RECT 2.560 153.475 158.420 156.305 ;
      LAYER pwell ;
        RECT 2.755 152.275 4.125 153.085 ;
        RECT 8.645 152.955 9.575 153.175 ;
        RECT 12.405 152.955 13.325 153.185 ;
        RECT 4.135 152.275 13.325 152.955 ;
        RECT 13.335 152.275 14.705 153.055 ;
        RECT 15.645 152.360 16.075 153.145 ;
        RECT 16.095 152.955 17.025 153.185 ;
        RECT 16.095 152.275 19.995 152.955 ;
        RECT 20.235 152.275 23.445 153.185 ;
        RECT 28.425 152.955 29.355 153.175 ;
        RECT 32.185 152.955 33.105 153.185 ;
        RECT 23.915 152.275 33.105 152.955 ;
        RECT 33.210 152.955 34.130 153.185 ;
        RECT 39.080 152.985 40.465 153.185 ;
        RECT 33.210 152.275 36.675 152.955 ;
        RECT 36.795 152.305 40.465 152.985 ;
        RECT 41.405 152.360 41.835 153.145 ;
        RECT 41.855 152.985 43.240 153.185 ;
        RECT 2.895 152.065 3.065 152.275 ;
        RECT 4.275 152.085 4.445 152.275 ;
        RECT 5.195 152.065 5.365 152.255 ;
        RECT 9.345 152.065 9.515 152.255 ;
        RECT 9.795 152.065 9.965 152.255 ;
        RECT 14.395 152.085 14.565 152.275 ;
        RECT 14.865 152.120 15.025 152.230 ;
        RECT 16.510 152.085 16.680 152.275 ;
        RECT 20.375 152.085 20.545 152.275 ;
        RECT 22.215 152.065 22.385 152.255 ;
        RECT 22.685 152.110 22.845 152.220 ;
        RECT 23.590 152.115 23.710 152.225 ;
        RECT 24.055 152.085 24.225 152.275 ;
        RECT 24.515 152.065 24.685 152.255 ;
        RECT 24.960 152.065 25.130 152.255 ;
        RECT 29.100 152.065 29.270 152.255 ;
        RECT 32.785 152.065 32.955 152.255 ;
        RECT 36.025 152.110 36.185 152.220 ;
        RECT 36.475 152.085 36.645 152.275 ;
        RECT 36.935 152.085 37.105 152.305 ;
        RECT 39.095 152.275 40.465 152.305 ;
        RECT 41.855 152.305 45.525 152.985 ;
        RECT 41.855 152.275 43.225 152.305 ;
        RECT 40.155 152.065 40.325 152.255 ;
        RECT 40.625 152.225 40.785 152.230 ;
        RECT 40.610 152.120 40.785 152.225 ;
        RECT 40.610 152.115 40.730 152.120 ;
        RECT 43.835 152.065 44.005 152.255 ;
        RECT 44.280 152.065 44.450 152.255 ;
        RECT 45.215 152.085 45.385 152.305 ;
        RECT 45.535 152.275 46.905 153.055 ;
        RECT 46.915 152.985 47.860 153.185 ;
        RECT 49.195 152.985 50.125 153.185 ;
        RECT 46.915 152.505 50.125 152.985 ;
        RECT 46.915 152.305 49.985 152.505 ;
        RECT 46.915 152.275 47.860 152.305 ;
        RECT 45.675 152.085 45.845 152.275 ;
        RECT 47.970 152.115 48.090 152.225 ;
        RECT 48.435 152.065 48.605 152.255 ;
        RECT 49.815 152.085 49.985 152.305 ;
        RECT 51.150 152.275 55.185 153.185 ;
        RECT 59.705 152.955 60.635 153.175 ;
        RECT 63.465 152.955 64.385 153.185 ;
        RECT 66.200 152.985 67.145 153.185 ;
        RECT 55.195 152.275 64.385 152.955 ;
        RECT 64.395 152.305 67.145 152.985 ;
        RECT 67.165 152.360 67.595 153.145 ;
        RECT 67.615 152.955 68.545 153.185 ;
        RECT 71.850 152.955 72.770 153.185 ;
        RECT 79.530 152.985 80.485 153.185 ;
        RECT 54.870 152.255 55.040 152.275 ;
        RECT 50.285 152.120 50.445 152.230 ;
        RECT 51.655 152.065 51.825 152.255 ;
        RECT 54.870 152.085 55.045 152.255 ;
        RECT 55.335 152.085 55.505 152.275 ;
        RECT 54.875 152.065 55.045 152.085 ;
        RECT 56.530 152.065 56.700 152.255 ;
        RECT 60.670 152.065 60.840 152.255 ;
        RECT 64.540 152.085 64.710 152.305 ;
        RECT 66.200 152.275 67.145 152.305 ;
        RECT 67.615 152.275 71.515 152.955 ;
        RECT 71.850 152.275 75.315 152.955 ;
        RECT 75.445 152.275 78.185 152.955 ;
        RECT 78.205 152.305 80.485 152.985 ;
        RECT 67.755 152.065 67.925 152.255 ;
        RECT 68.030 152.085 68.200 152.275 ;
        RECT 68.210 152.065 68.380 152.255 ;
        RECT 75.115 152.085 75.285 152.275 ;
        RECT 77.875 152.085 78.045 152.275 ;
        RECT 78.330 152.255 78.500 152.305 ;
        RECT 79.530 152.275 80.485 152.305 ;
        RECT 80.495 152.985 81.450 153.185 ;
        RECT 80.495 152.305 82.775 152.985 ;
        RECT 86.455 152.955 87.385 153.185 ;
        RECT 80.495 152.275 81.450 152.305 ;
        RECT 78.330 152.085 78.505 152.255 ;
        RECT 78.335 152.065 78.505 152.085 ;
        RECT 78.795 152.065 78.965 152.255 ;
        RECT 80.635 152.065 80.805 152.255 ;
        RECT 82.480 152.085 82.650 152.305 ;
        RECT 83.485 152.275 87.385 152.955 ;
        RECT 87.395 152.275 88.765 153.085 ;
        RECT 88.775 152.955 89.705 153.185 ;
        RECT 88.775 152.275 92.675 152.955 ;
        RECT 92.925 152.360 93.355 153.145 ;
        RECT 93.375 152.275 94.745 153.055 ;
        RECT 82.930 152.115 83.050 152.225 ;
        RECT 86.800 152.085 86.970 152.275 ;
        RECT 87.535 152.085 87.705 152.275 ;
        RECT 89.190 152.085 89.360 152.275 ;
        RECT 89.840 152.065 90.010 152.255 ;
        RECT 94.435 152.085 94.605 152.275 ;
        RECT 95.695 152.235 96.585 153.185 ;
        RECT 100.715 152.955 101.645 153.185 ;
        RECT 97.745 152.275 101.645 152.955 ;
        RECT 101.655 152.275 103.485 153.085 ;
        RECT 108.005 152.955 108.935 153.175 ;
        RECT 111.765 152.955 113.105 153.185 ;
        RECT 103.495 152.275 113.105 152.955 ;
        RECT 113.155 152.275 114.525 153.055 ;
        RECT 117.735 152.955 118.665 153.185 ;
        RECT 114.765 152.275 118.665 152.955 ;
        RECT 118.685 152.360 119.115 153.145 ;
        RECT 120.940 152.985 121.885 153.185 ;
        RECT 119.135 152.305 121.885 152.985 ;
        RECT 126.405 152.955 127.335 153.175 ;
        RECT 130.165 152.955 131.085 153.185 ;
        RECT 94.905 152.120 95.065 152.230 ;
        RECT 95.365 152.110 95.525 152.220 ;
        RECT 95.815 152.085 95.985 152.235 ;
        RECT 96.275 152.105 96.445 152.235 ;
        RECT 96.745 152.120 96.905 152.230 ;
        RECT 97.205 152.110 97.365 152.220 ;
        RECT 2.755 151.255 4.125 152.065 ;
        RECT 5.055 151.285 6.425 152.065 ;
        RECT 6.435 151.155 9.645 152.065 ;
        RECT 9.655 151.385 18.845 152.065 ;
        RECT 14.165 151.165 15.095 151.385 ;
        RECT 17.925 151.155 18.845 151.385 ;
        RECT 18.950 151.385 22.415 152.065 ;
        RECT 18.950 151.155 19.870 151.385 ;
        RECT 23.465 151.155 24.815 152.065 ;
        RECT 24.845 151.155 28.505 152.065 ;
        RECT 28.525 151.195 28.955 151.980 ;
        RECT 28.985 151.155 32.645 152.065 ;
        RECT 32.655 151.155 35.865 152.065 ;
        RECT 36.890 151.385 40.355 152.065 ;
        RECT 36.890 151.155 37.810 151.385 ;
        RECT 40.935 151.155 44.145 152.065 ;
        RECT 44.165 151.155 47.825 152.065 ;
        RECT 48.295 151.155 51.505 152.065 ;
        RECT 51.525 151.155 54.255 152.065 ;
        RECT 54.285 151.195 54.715 151.980 ;
        RECT 54.735 151.285 56.105 152.065 ;
        RECT 56.115 151.385 60.015 152.065 ;
        RECT 60.255 151.385 64.155 152.065 ;
        RECT 64.490 151.385 67.955 152.065 ;
        RECT 56.115 151.155 57.045 151.385 ;
        RECT 60.255 151.155 61.185 151.385 ;
        RECT 64.490 151.155 65.410 151.385 ;
        RECT 68.095 151.155 69.445 152.065 ;
        RECT 69.540 151.385 78.645 152.065 ;
        RECT 78.655 151.255 80.025 152.065 ;
        RECT 80.045 151.195 80.475 151.980 ;
        RECT 80.495 151.385 89.685 152.065 ;
        RECT 85.005 151.165 85.935 151.385 ;
        RECT 88.765 151.155 89.685 151.385 ;
        RECT 89.695 151.155 95.205 152.065 ;
        RECT 96.155 151.155 97.045 152.105 ;
        RECT 98.120 152.065 98.290 152.255 ;
        RECT 101.060 152.085 101.230 152.275 ;
        RECT 101.795 152.085 101.965 152.275 ;
        RECT 102.255 152.085 102.425 152.255 ;
        RECT 103.635 152.085 103.805 152.275 ;
        RECT 102.260 152.065 102.425 152.085 ;
        RECT 104.555 152.065 104.725 152.255 ;
        RECT 106.405 152.110 106.565 152.220 ;
        RECT 107.775 152.105 107.945 152.255 ;
        RECT 97.975 151.385 102.105 152.065 ;
        RECT 102.260 151.385 104.095 152.065 ;
        RECT 97.975 151.155 99.315 151.385 ;
        RECT 103.165 151.155 104.095 151.385 ;
        RECT 104.415 151.255 105.785 152.065 ;
        RECT 105.805 151.195 106.235 151.980 ;
        RECT 107.175 151.155 108.065 152.105 ;
        RECT 113.295 152.085 113.465 152.275 ;
        RECT 113.755 152.065 113.925 152.255 ;
        RECT 114.215 152.085 114.385 152.255 ;
        RECT 118.080 152.085 118.250 152.275 ;
        RECT 119.280 152.085 119.450 152.305 ;
        RECT 120.940 152.275 121.885 152.305 ;
        RECT 121.895 152.275 131.085 152.955 ;
        RECT 122.035 152.085 122.205 152.275 ;
        RECT 114.220 152.065 114.385 152.085 ;
        RECT 125.715 152.065 125.885 152.255 ;
        RECT 126.170 152.065 126.340 152.255 ;
        RECT 130.960 152.065 131.130 152.255 ;
        RECT 132.035 152.235 132.925 153.185 ;
        RECT 136.645 152.955 137.985 153.185 ;
        RECT 133.855 152.275 137.985 152.955 ;
        RECT 137.995 152.275 139.365 153.055 ;
        RECT 139.375 152.275 140.745 153.055 ;
        RECT 140.755 152.275 144.425 153.085 ;
        RECT 144.445 152.360 144.875 153.145 ;
        RECT 144.895 152.275 150.405 153.085 ;
        RECT 150.415 152.275 155.925 153.085 ;
        RECT 156.855 152.275 158.225 153.085 ;
        RECT 131.245 152.120 131.405 152.230 ;
        RECT 132.155 152.225 132.325 152.235 ;
        RECT 132.150 152.115 132.325 152.225 ;
        RECT 132.155 152.085 132.325 152.115 ;
        RECT 132.615 152.065 132.785 152.235 ;
        RECT 133.085 152.120 133.245 152.230 ;
        RECT 137.670 152.085 137.840 152.275 ;
        RECT 138.135 152.085 138.305 152.275 ;
        RECT 140.435 152.085 140.605 152.275 ;
        RECT 140.895 152.085 141.065 152.275 ;
        RECT 144.115 152.065 144.285 152.255 ;
        RECT 144.575 152.065 144.745 152.255 ;
        RECT 145.035 152.085 145.205 152.275 ;
        RECT 150.095 152.065 150.265 152.255 ;
        RECT 150.555 152.085 150.725 152.275 ;
        RECT 155.615 152.065 155.785 152.255 ;
        RECT 156.085 152.120 156.245 152.230 ;
        RECT 157.915 152.065 158.085 152.275 ;
        RECT 108.310 151.155 114.040 152.065 ;
        RECT 114.220 151.385 116.055 152.065 ;
        RECT 115.125 151.155 116.055 151.385 ;
        RECT 116.415 151.385 126.025 152.065 ;
        RECT 116.415 151.155 117.755 151.385 ;
        RECT 120.585 151.165 121.515 151.385 ;
        RECT 126.055 151.155 127.405 152.065 ;
        RECT 127.645 151.385 131.545 152.065 ;
        RECT 130.615 151.155 131.545 151.385 ;
        RECT 131.565 151.195 131.995 151.980 ;
        RECT 132.475 151.385 141.665 152.065 ;
        RECT 141.685 151.385 144.425 152.065 ;
        RECT 136.985 151.165 137.915 151.385 ;
        RECT 140.745 151.155 141.665 151.385 ;
        RECT 144.435 151.255 149.945 152.065 ;
        RECT 149.955 151.255 155.465 152.065 ;
        RECT 155.475 151.255 156.845 152.065 ;
        RECT 156.855 151.255 158.225 152.065 ;
      LAYER nwell ;
        RECT 2.560 148.035 158.420 150.865 ;
      LAYER pwell ;
        RECT 2.755 146.835 4.125 147.645 ;
        RECT 8.645 147.515 9.575 147.735 ;
        RECT 12.405 147.515 13.325 147.745 ;
        RECT 4.135 146.835 13.325 147.515 ;
        RECT 13.335 146.835 14.705 147.615 ;
        RECT 15.645 146.920 16.075 147.705 ;
        RECT 16.095 147.515 17.025 147.745 ;
        RECT 20.330 147.515 21.250 147.745 ;
        RECT 16.095 146.835 19.995 147.515 ;
        RECT 20.330 146.835 23.795 147.515 ;
        RECT 23.915 146.835 25.285 147.615 ;
        RECT 25.755 146.835 28.965 147.745 ;
        RECT 28.975 146.835 32.185 147.745 ;
        RECT 32.205 146.835 35.865 147.745 ;
        RECT 35.875 146.835 37.705 147.515 ;
        RECT 37.730 146.835 41.385 147.745 ;
        RECT 41.405 146.920 41.835 147.705 ;
        RECT 41.935 146.835 44.145 147.745 ;
        RECT 44.155 146.835 47.810 147.745 ;
        RECT 47.845 146.835 51.505 147.745 ;
        RECT 51.525 146.835 55.185 147.745 ;
        RECT 56.530 147.545 57.485 147.745 ;
        RECT 55.205 146.865 57.485 147.545 ;
        RECT 2.895 146.625 3.065 146.835 ;
        RECT 4.275 146.645 4.445 146.835 ;
        RECT 5.185 146.625 5.355 146.815 ;
        RECT 8.690 146.625 8.860 146.815 ;
        RECT 12.830 146.625 13.000 146.815 ;
        RECT 14.395 146.645 14.565 146.835 ;
        RECT 14.865 146.680 15.025 146.790 ;
        RECT 16.510 146.645 16.680 146.835 ;
        RECT 16.690 146.675 16.810 146.785 ;
        RECT 17.155 146.625 17.325 146.815 ;
        RECT 23.145 146.625 23.315 146.815 ;
        RECT 23.595 146.625 23.765 146.835 ;
        RECT 24.975 146.815 25.145 146.835 ;
        RECT 24.960 146.645 25.145 146.815 ;
        RECT 25.430 146.675 25.550 146.785 ;
        RECT 25.895 146.645 26.065 146.835 ;
        RECT 29.115 146.645 29.285 146.835 ;
        RECT 24.960 146.625 25.130 146.645 ;
        RECT 30.955 146.625 31.125 146.815 ;
        RECT 32.320 146.645 32.490 146.835 ;
        RECT 34.635 146.625 34.805 146.815 ;
        RECT 35.095 146.625 35.265 146.815 ;
        RECT 36.015 146.645 36.185 146.835 ;
        RECT 38.775 146.625 38.945 146.815 ;
        RECT 41.070 146.645 41.240 146.835 ;
        RECT 43.830 146.645 44.000 146.835 ;
        RECT 44.300 146.645 44.470 146.835 ;
        RECT 47.960 146.645 48.130 146.835 ;
        RECT 48.420 146.625 48.590 146.815 ;
        RECT 51.640 146.645 51.810 146.835 ;
        RECT 52.125 146.670 52.285 146.780 ;
        RECT 53.035 146.625 53.205 146.815 ;
        RECT 55.330 146.645 55.500 146.865 ;
        RECT 56.530 146.835 57.485 146.865 ;
        RECT 57.495 147.515 58.415 147.745 ;
        RECT 61.245 147.515 62.175 147.735 ;
        RECT 57.495 146.835 66.685 147.515 ;
        RECT 67.165 146.920 67.595 147.705 ;
        RECT 67.615 146.835 68.985 147.615 ;
        RECT 73.505 147.515 74.435 147.735 ;
        RECT 77.265 147.515 78.185 147.745 ;
        RECT 68.995 146.835 78.185 147.515 ;
        RECT 78.195 147.515 79.535 147.745 ;
        RECT 85.535 147.515 86.465 147.745 ;
        RECT 78.195 146.835 82.325 147.515 ;
        RECT 82.565 146.835 86.465 147.515 ;
        RECT 87.395 147.515 88.740 147.745 ;
        RECT 87.395 146.835 89.225 147.515 ;
        RECT 89.775 146.835 92.775 147.745 ;
        RECT 92.925 146.920 93.355 147.705 ;
        RECT 97.885 147.515 98.815 147.735 ;
        RECT 101.645 147.515 102.565 147.745 ;
        RECT 93.375 146.835 102.565 147.515 ;
        RECT 102.575 146.835 104.405 147.645 ;
        RECT 104.630 146.835 110.360 147.745 ;
        RECT 110.855 146.835 112.205 147.745 ;
        RECT 115.025 147.515 116.365 147.745 ;
        RECT 112.235 146.835 116.365 147.515 ;
        RECT 117.295 146.835 118.645 147.745 ;
        RECT 118.685 146.920 119.115 147.705 ;
        RECT 119.595 146.835 122.805 147.745 ;
        RECT 123.010 146.835 126.485 147.745 ;
        RECT 129.695 147.515 130.625 147.745 ;
        RECT 126.725 146.835 130.625 147.515 ;
        RECT 131.555 146.835 133.385 147.745 ;
        RECT 138.365 147.515 139.295 147.735 ;
        RECT 142.015 147.515 144.225 147.745 ;
        RECT 133.855 146.835 144.225 147.515 ;
        RECT 144.445 146.920 144.875 147.705 ;
        RECT 144.895 146.835 150.405 147.645 ;
        RECT 150.415 146.835 155.925 147.645 ;
        RECT 156.855 146.835 158.225 147.645 ;
        RECT 55.800 146.625 55.970 146.815 ;
        RECT 56.250 146.675 56.370 146.785 ;
        RECT 60.120 146.625 60.290 146.815 ;
        RECT 60.855 146.625 61.025 146.815 ;
        RECT 62.695 146.625 62.865 146.815 ;
        RECT 66.375 146.645 66.545 146.835 ;
        RECT 66.830 146.675 66.950 146.785 ;
        RECT 68.675 146.645 68.845 146.835 ;
        RECT 69.135 146.645 69.305 146.835 ;
        RECT 75.300 146.625 75.470 146.815 ;
        RECT 78.340 146.645 78.510 146.835 ;
        RECT 79.710 146.625 79.880 146.815 ;
        RECT 84.040 146.625 84.210 146.815 ;
        RECT 84.775 146.625 84.945 146.815 ;
        RECT 85.880 146.645 86.050 146.835 ;
        RECT 86.625 146.785 86.785 146.790 ;
        RECT 86.610 146.680 86.785 146.785 ;
        RECT 86.610 146.675 86.730 146.680 ;
        RECT 87.075 146.645 87.245 146.815 ;
        RECT 88.915 146.645 89.085 146.835 ;
        RECT 89.370 146.675 89.490 146.785 ;
        RECT 87.080 146.625 87.245 146.645 ;
        RECT 89.835 146.625 90.005 146.835 ;
        RECT 92.590 146.675 92.710 146.785 ;
        RECT 93.055 146.625 93.225 146.815 ;
        RECT 93.515 146.645 93.685 146.835 ;
        RECT 95.825 146.670 95.985 146.780 ;
        RECT 97.195 146.665 97.365 146.815 ;
        RECT 97.665 146.670 97.825 146.780 ;
        RECT 2.755 145.815 4.125 146.625 ;
        RECT 5.055 145.715 8.265 146.625 ;
        RECT 8.275 145.945 12.175 146.625 ;
        RECT 12.415 145.945 16.315 146.625 ;
        RECT 8.275 145.715 9.205 145.945 ;
        RECT 12.415 145.715 13.345 145.945 ;
        RECT 17.015 145.715 20.225 146.625 ;
        RECT 20.235 145.715 23.445 146.625 ;
        RECT 23.455 145.845 24.825 146.625 ;
        RECT 24.845 145.715 28.505 146.625 ;
        RECT 28.525 145.755 28.955 146.540 ;
        RECT 29.905 145.715 31.255 146.625 ;
        RECT 31.370 145.945 34.835 146.625 ;
        RECT 35.065 145.945 38.530 146.625 ;
        RECT 38.635 145.945 47.825 146.625 ;
        RECT 31.370 145.715 32.290 145.945 ;
        RECT 37.610 145.715 38.530 145.945 ;
        RECT 43.145 145.725 44.075 145.945 ;
        RECT 46.905 145.715 47.825 145.945 ;
        RECT 48.305 145.715 51.965 146.625 ;
        RECT 52.895 145.845 54.265 146.625 ;
        RECT 54.285 145.755 54.715 146.540 ;
        RECT 54.735 145.715 56.085 146.625 ;
        RECT 56.805 145.945 60.705 146.625 ;
        RECT 60.715 145.945 62.545 146.625 ;
        RECT 62.555 145.945 71.745 146.625 ;
        RECT 71.985 145.945 75.885 146.625 ;
        RECT 75.895 145.945 80.025 146.625 ;
        RECT 59.775 145.715 60.705 145.945 ;
        RECT 61.200 145.715 62.545 145.945 ;
        RECT 67.065 145.725 67.995 145.945 ;
        RECT 70.825 145.715 71.745 145.945 ;
        RECT 74.955 145.715 75.885 145.945 ;
        RECT 78.685 145.715 80.025 145.945 ;
        RECT 80.045 145.755 80.475 146.540 ;
        RECT 80.725 145.945 84.625 146.625 ;
        RECT 83.695 145.715 84.625 145.945 ;
        RECT 84.635 145.815 86.465 146.625 ;
        RECT 87.080 145.945 88.915 146.625 ;
        RECT 87.985 145.715 88.915 145.945 ;
        RECT 89.695 145.715 92.100 146.625 ;
        RECT 92.915 145.715 95.665 146.625 ;
        RECT 96.595 145.715 97.485 146.665 ;
        RECT 100.415 146.645 100.585 146.815 ;
        RECT 100.875 146.645 101.045 146.815 ;
        RECT 102.715 146.645 102.885 146.835 ;
        RECT 103.185 146.670 103.345 146.780 ;
        RECT 104.555 146.665 104.725 146.815 ;
        RECT 105.025 146.670 105.185 146.780 ;
        RECT 100.415 146.625 100.580 146.645 ;
        RECT 98.745 145.945 100.580 146.625 ;
        RECT 100.880 146.625 101.045 146.645 ;
        RECT 100.880 145.945 102.715 146.625 ;
        RECT 98.745 145.715 99.675 145.945 ;
        RECT 101.785 145.715 102.715 145.945 ;
        RECT 103.955 145.715 104.845 146.665 ;
        RECT 110.075 146.645 110.245 146.835 ;
        RECT 110.530 146.675 110.650 146.785 ;
        RECT 111.000 146.645 111.170 146.835 ;
        RECT 111.915 146.625 112.085 146.815 ;
        RECT 116.050 146.625 116.220 146.835 ;
        RECT 116.525 146.670 116.685 146.790 ;
        RECT 117.440 146.625 117.610 146.815 ;
        RECT 118.360 146.645 118.530 146.835 ;
        RECT 119.270 146.675 119.390 146.785 ;
        RECT 122.505 146.645 122.675 146.835 ;
        RECT 126.170 146.645 126.340 146.835 ;
        RECT 127.090 146.675 127.210 146.785 ;
        RECT 130.040 146.645 130.210 146.835 ;
        RECT 130.785 146.680 130.945 146.790 ;
        RECT 130.960 146.625 131.130 146.815 ;
        RECT 132.155 146.625 132.325 146.815 ;
        RECT 133.070 146.645 133.240 146.835 ;
        RECT 133.995 146.785 134.165 146.835 ;
        RECT 133.530 146.675 133.650 146.785 ;
        RECT 133.990 146.675 134.165 146.785 ;
        RECT 133.995 146.645 134.165 146.675 ;
        RECT 134.455 146.625 134.625 146.815 ;
        RECT 144.575 146.625 144.745 146.815 ;
        RECT 145.035 146.645 145.205 146.835 ;
        RECT 145.955 146.625 146.125 146.815 ;
        RECT 146.415 146.625 146.585 146.815 ;
        RECT 150.555 146.645 150.725 146.835 ;
        RECT 151.935 146.625 152.105 146.815 ;
        RECT 155.615 146.625 155.785 146.815 ;
        RECT 156.085 146.680 156.245 146.790 ;
        RECT 157.915 146.625 158.085 146.835 ;
        RECT 105.805 145.755 106.235 146.540 ;
        RECT 106.470 145.715 112.200 146.625 ;
        RECT 112.235 145.945 116.365 146.625 ;
        RECT 115.025 145.715 116.365 145.945 ;
        RECT 117.295 145.715 126.820 146.625 ;
        RECT 127.645 145.945 131.545 146.625 ;
        RECT 130.615 145.715 131.545 145.945 ;
        RECT 131.565 145.755 131.995 146.540 ;
        RECT 132.030 145.715 133.845 146.625 ;
        RECT 134.315 145.945 143.505 146.625 ;
        RECT 138.825 145.725 139.755 145.945 ;
        RECT 142.585 145.715 143.505 145.945 ;
        RECT 143.515 145.845 144.885 146.625 ;
        RECT 144.895 145.845 146.265 146.625 ;
        RECT 146.275 145.815 151.785 146.625 ;
        RECT 151.795 145.815 155.465 146.625 ;
        RECT 155.475 145.815 156.845 146.625 ;
        RECT 156.855 145.815 158.225 146.625 ;
      LAYER nwell ;
        RECT 2.560 142.595 158.420 145.425 ;
      LAYER pwell ;
        RECT 2.755 141.395 4.125 142.205 ;
        RECT 5.495 142.075 6.415 142.295 ;
        RECT 12.495 142.195 13.415 142.305 ;
        RECT 11.080 142.075 13.415 142.195 ;
        RECT 4.135 141.395 13.415 142.075 ;
        RECT 13.795 141.395 15.165 142.175 ;
        RECT 15.645 141.480 16.075 142.265 ;
        RECT 16.095 142.075 17.025 142.305 ;
        RECT 16.095 141.395 19.995 142.075 ;
        RECT 20.695 141.395 23.905 142.305 ;
        RECT 23.915 141.395 25.285 142.175 ;
        RECT 25.850 142.075 26.770 142.305 ;
        RECT 33.945 142.075 34.875 142.295 ;
        RECT 37.705 142.075 38.625 142.305 ;
        RECT 25.850 141.395 29.315 142.075 ;
        RECT 29.435 141.395 38.625 142.075 ;
        RECT 38.645 141.395 41.375 142.305 ;
        RECT 41.405 141.480 41.835 142.265 ;
        RECT 41.855 142.075 42.785 142.305 ;
        RECT 46.090 142.075 47.010 142.305 ;
        RECT 41.855 141.395 45.755 142.075 ;
        RECT 46.090 141.395 49.555 142.075 ;
        RECT 49.675 141.395 53.330 142.305 ;
        RECT 56.555 142.075 57.485 142.305 ;
        RECT 53.585 141.395 57.485 142.075 ;
        RECT 57.865 142.195 58.785 142.305 ;
        RECT 57.865 142.075 60.200 142.195 ;
        RECT 64.865 142.075 65.785 142.295 ;
        RECT 57.865 141.395 67.145 142.075 ;
        RECT 67.165 141.480 67.595 142.265 ;
        RECT 67.760 141.395 70.825 142.305 ;
        RECT 71.755 142.105 72.685 142.305 ;
        RECT 74.020 142.105 74.965 142.305 ;
        RECT 71.755 141.625 74.965 142.105 ;
        RECT 78.685 142.075 80.025 142.305 ;
        RECT 71.895 141.425 74.965 141.625 ;
        RECT 2.895 141.185 3.065 141.395 ;
        RECT 4.275 141.345 4.445 141.395 ;
        RECT 4.270 141.235 4.445 141.345 ;
        RECT 4.275 141.205 4.445 141.235 ;
        RECT 4.735 141.185 4.905 141.375 ;
        RECT 10.715 141.185 10.885 141.375 ;
        RECT 11.175 141.185 11.345 141.375 ;
        RECT 14.855 141.205 15.025 141.395 ;
        RECT 15.310 141.235 15.430 141.345 ;
        RECT 16.510 141.205 16.680 141.395 ;
        RECT 20.370 141.235 20.490 141.345 ;
        RECT 23.605 141.205 23.775 141.395 ;
        RECT 24.055 141.185 24.225 141.395 ;
        RECT 24.790 141.185 24.960 141.375 ;
        RECT 25.430 141.235 25.550 141.345 ;
        RECT 29.115 141.205 29.285 141.395 ;
        RECT 29.390 141.185 29.560 141.375 ;
        RECT 29.575 141.205 29.745 141.395 ;
        RECT 33.530 141.185 33.700 141.375 ;
        RECT 40.800 141.185 40.970 141.375 ;
        RECT 41.075 141.205 41.245 141.395 ;
        RECT 42.270 141.205 42.440 141.395 ;
        RECT 43.835 141.185 44.005 141.375 ;
        RECT 44.570 141.185 44.740 141.375 ;
        RECT 48.430 141.235 48.550 141.345 ;
        RECT 48.895 141.185 49.065 141.375 ;
        RECT 49.355 141.205 49.525 141.395 ;
        RECT 49.820 141.205 49.990 141.395 ;
        RECT 53.680 141.185 53.850 141.375 ;
        RECT 54.875 141.185 55.045 141.375 ;
        RECT 56.900 141.205 57.070 141.395 ;
        RECT 66.835 141.205 67.005 141.395 ;
        RECT 67.295 141.185 67.465 141.375 ;
        RECT 67.750 141.235 67.870 141.345 ;
        RECT 70.510 141.205 70.680 141.395 ;
        RECT 70.975 141.185 71.145 141.375 ;
        RECT 71.895 141.205 72.065 141.425 ;
        RECT 74.020 141.395 74.965 141.425 ;
        RECT 75.895 141.395 80.025 142.075 ;
        RECT 80.035 141.395 81.405 142.205 ;
        RECT 83.220 142.105 84.165 142.305 ;
        RECT 81.415 141.425 84.165 142.105 ;
        RECT 74.650 141.185 74.820 141.375 ;
        RECT 75.125 141.240 75.285 141.350 ;
        RECT 78.790 141.185 78.960 141.375 ;
        RECT 79.265 141.230 79.425 141.340 ;
        RECT 79.710 141.205 79.880 141.395 ;
        RECT 80.175 141.205 80.345 141.395 ;
        RECT 81.560 141.205 81.730 141.425 ;
        RECT 83.220 141.395 84.165 141.425 ;
        RECT 84.175 141.395 86.925 142.205 ;
        RECT 87.035 141.395 89.225 142.305 ;
        RECT 89.235 141.395 92.445 142.305 ;
        RECT 92.925 141.480 93.355 142.265 ;
        RECT 93.375 141.395 97.045 142.205 ;
        RECT 97.975 141.395 100.725 142.305 ;
        RECT 100.755 141.395 102.105 142.305 ;
        RECT 102.670 141.395 106.705 142.305 ;
        RECT 106.715 141.395 113.225 142.305 ;
        RECT 116.405 142.075 117.745 142.305 ;
        RECT 113.615 141.395 117.745 142.075 ;
        RECT 118.685 141.480 119.115 142.265 ;
        RECT 119.150 141.395 122.805 142.305 ;
        RECT 122.815 141.395 126.290 142.305 ;
        RECT 126.495 141.395 129.415 142.305 ;
        RECT 129.725 141.395 132.455 142.305 ;
        RECT 133.395 141.395 139.905 142.305 ;
        RECT 140.295 141.395 142.905 142.305 ;
        RECT 143.055 141.395 144.405 142.305 ;
        RECT 144.445 141.480 144.875 142.265 ;
        RECT 144.905 141.395 147.645 142.075 ;
        RECT 147.655 141.395 153.165 142.205 ;
        RECT 153.175 141.395 156.845 142.205 ;
        RECT 156.855 141.395 158.225 142.205 ;
        RECT 84.315 141.205 84.485 141.395 ;
        RECT 86.155 141.185 86.325 141.375 ;
        RECT 86.615 141.185 86.785 141.375 ;
        RECT 87.995 141.185 88.165 141.375 ;
        RECT 88.910 141.205 89.080 141.395 ;
        RECT 92.135 141.185 92.305 141.395 ;
        RECT 92.595 141.345 92.765 141.375 ;
        RECT 92.590 141.235 92.765 141.345 ;
        RECT 92.595 141.185 92.765 141.235 ;
        RECT 93.515 141.205 93.685 141.395 ;
        RECT 96.285 141.230 96.445 141.340 ;
        RECT 97.200 141.185 97.370 141.375 ;
        RECT 98.115 141.205 98.285 141.395 ;
        RECT 100.870 141.205 101.040 141.395 ;
        RECT 106.390 141.375 106.560 141.395 ;
        RECT 102.250 141.235 102.370 141.345 ;
        RECT 104.090 141.185 104.260 141.375 ;
        RECT 104.555 141.185 104.725 141.375 ;
        RECT 106.390 141.205 106.570 141.375 ;
        RECT 106.860 141.205 107.030 141.395 ;
        RECT 106.400 141.185 106.570 141.205 ;
        RECT 110.540 141.185 110.710 141.375 ;
        RECT 2.755 140.375 4.125 141.185 ;
        RECT 4.595 140.275 7.805 141.185 ;
        RECT 7.815 140.275 11.025 141.185 ;
        RECT 11.035 140.505 20.315 141.185 ;
        RECT 12.395 140.285 13.315 140.505 ;
        RECT 17.980 140.385 20.315 140.505 ;
        RECT 19.395 140.275 20.315 140.385 ;
        RECT 20.790 140.505 24.255 141.185 ;
        RECT 24.375 140.505 28.275 141.185 ;
        RECT 20.790 140.275 21.710 140.505 ;
        RECT 24.375 140.275 25.305 140.505 ;
        RECT 28.525 140.315 28.955 141.100 ;
        RECT 28.975 140.505 32.875 141.185 ;
        RECT 33.115 140.505 37.015 141.185 ;
        RECT 37.485 140.505 41.385 141.185 ;
        RECT 41.405 140.505 44.145 141.185 ;
        RECT 44.155 140.505 48.055 141.185 ;
        RECT 28.975 140.275 29.905 140.505 ;
        RECT 33.115 140.275 34.045 140.505 ;
        RECT 40.455 140.275 41.385 140.505 ;
        RECT 44.155 140.275 45.085 140.505 ;
        RECT 48.755 140.405 50.125 141.185 ;
        RECT 50.365 140.505 54.265 141.185 ;
        RECT 53.335 140.275 54.265 140.505 ;
        RECT 54.285 140.315 54.715 141.100 ;
        RECT 54.735 140.505 63.925 141.185 ;
        RECT 59.245 140.285 60.175 140.505 ;
        RECT 63.005 140.275 63.925 140.505 ;
        RECT 64.030 140.505 67.495 141.185 ;
        RECT 69.445 141.155 71.285 141.185 ;
        RECT 68.120 140.505 71.285 141.155 ;
        RECT 64.030 140.275 64.950 140.505 ;
        RECT 68.120 140.475 70.800 140.505 ;
        RECT 69.445 140.275 70.800 140.475 ;
        RECT 71.310 140.275 74.965 141.185 ;
        RECT 75.235 140.275 79.105 141.185 ;
        RECT 80.045 140.315 80.475 141.100 ;
        RECT 80.625 140.275 86.465 141.185 ;
        RECT 86.475 140.375 87.845 141.185 ;
        RECT 87.855 140.275 91.065 141.185 ;
        RECT 91.085 140.275 92.435 141.185 ;
        RECT 92.455 140.375 96.125 141.185 ;
        RECT 97.055 140.505 100.725 141.185 ;
        RECT 97.055 140.275 97.980 140.505 ;
        RECT 100.750 140.275 104.405 141.185 ;
        RECT 104.415 140.375 105.785 141.185 ;
        RECT 105.805 140.315 106.235 141.100 ;
        RECT 106.255 140.505 110.350 141.185 ;
        RECT 106.740 140.275 110.350 140.505 ;
        RECT 110.395 140.275 112.585 141.185 ;
        RECT 112.840 141.155 113.010 141.375 ;
        RECT 116.055 141.185 116.225 141.375 ;
        RECT 117.430 141.205 117.600 141.395 ;
        RECT 117.905 141.240 118.065 141.350 ;
        RECT 119.275 141.185 119.445 141.375 ;
        RECT 122.490 141.205 122.660 141.395 ;
        RECT 122.960 141.205 123.130 141.395 ;
        RECT 124.330 141.185 124.500 141.375 ;
        RECT 124.790 141.235 124.910 141.345 ;
        RECT 125.260 141.185 125.430 141.375 ;
        RECT 126.640 141.205 126.810 141.395 ;
        RECT 129.855 141.205 130.025 141.395 ;
        RECT 131.235 141.185 131.405 141.375 ;
        RECT 132.155 141.185 132.325 141.375 ;
        RECT 132.625 141.240 132.785 141.350 ;
        RECT 133.540 141.205 133.710 141.395 ;
        RECT 140.440 141.375 140.610 141.395 ;
        RECT 134.925 141.230 135.085 141.340 ;
        RECT 140.430 141.205 140.610 141.375 ;
        RECT 140.430 141.185 140.600 141.205 ;
        RECT 114.970 141.155 115.905 141.185 ;
        RECT 112.840 140.955 115.905 141.155 ;
        RECT 112.695 140.475 115.905 140.955 ;
        RECT 112.695 140.275 113.625 140.475 ;
        RECT 114.955 140.275 115.905 140.475 ;
        RECT 115.955 140.275 119.125 141.185 ;
        RECT 119.135 140.275 121.885 141.185 ;
        RECT 122.035 140.275 124.645 141.185 ;
        RECT 125.115 140.275 128.770 141.185 ;
        RECT 128.805 140.275 131.535 141.185 ;
        RECT 131.565 140.315 131.995 141.100 ;
        RECT 132.015 140.275 134.765 141.185 ;
        RECT 135.875 140.275 140.745 141.185 ;
        RECT 140.900 141.155 141.070 141.375 ;
        RECT 143.200 141.205 143.370 141.395 ;
        RECT 143.030 141.155 143.965 141.185 ;
        RECT 140.900 140.955 143.965 141.155 ;
        RECT 140.755 140.475 143.965 140.955 ;
        RECT 140.755 140.275 141.685 140.475 ;
        RECT 143.015 140.275 143.965 140.475 ;
        RECT 143.975 141.155 144.910 141.185 ;
        RECT 146.870 141.155 147.040 141.375 ;
        RECT 147.335 141.205 147.505 141.395 ;
        RECT 147.795 141.205 147.965 141.395 ;
        RECT 148.260 141.185 148.430 141.375 ;
        RECT 148.715 141.185 148.885 141.375 ;
        RECT 153.315 141.205 153.485 141.395 ;
        RECT 154.235 141.185 154.405 141.375 ;
        RECT 157.915 141.185 158.085 141.395 ;
        RECT 143.975 140.955 147.040 141.155 ;
        RECT 143.975 140.475 147.185 140.955 ;
        RECT 143.975 140.275 144.925 140.475 ;
        RECT 146.255 140.275 147.185 140.475 ;
        RECT 147.195 140.275 148.545 141.185 ;
        RECT 148.575 140.375 154.085 141.185 ;
        RECT 154.095 140.375 156.845 141.185 ;
        RECT 156.855 140.375 158.225 141.185 ;
      LAYER nwell ;
        RECT 2.560 137.155 158.420 139.985 ;
      LAYER pwell ;
        RECT 2.755 135.955 4.125 136.765 ;
        RECT 8.645 136.635 9.575 136.855 ;
        RECT 12.405 136.635 13.325 136.865 ;
        RECT 4.135 135.955 13.325 136.635 ;
        RECT 14.255 135.955 15.625 136.735 ;
        RECT 15.645 136.040 16.075 136.825 ;
        RECT 16.095 136.635 17.025 136.865 ;
        RECT 16.095 135.955 19.995 136.635 ;
        RECT 20.235 135.955 22.065 136.765 ;
        RECT 26.585 136.635 27.515 136.855 ;
        RECT 30.345 136.635 31.265 136.865 ;
        RECT 22.075 135.955 31.265 136.635 ;
        RECT 32.195 136.635 33.115 136.865 ;
        RECT 35.945 136.635 36.875 136.855 ;
        RECT 32.195 135.955 41.385 136.635 ;
        RECT 41.405 136.040 41.835 136.825 ;
        RECT 47.285 136.635 48.215 136.855 ;
        RECT 51.045 136.635 51.965 136.865 ;
        RECT 42.775 135.955 51.965 136.635 ;
        RECT 52.435 135.955 53.805 136.735 ;
        RECT 53.815 136.635 54.745 136.865 ;
        RECT 62.465 136.635 63.395 136.855 ;
        RECT 66.225 136.635 67.145 136.865 ;
        RECT 53.815 135.955 57.715 136.635 ;
        RECT 57.955 135.955 67.145 136.635 ;
        RECT 67.165 136.040 67.595 136.825 ;
        RECT 67.625 135.955 68.975 136.865 ;
        RECT 68.995 135.955 71.605 136.865 ;
        RECT 71.855 135.955 74.965 136.865 ;
        RECT 74.975 135.955 76.805 136.765 ;
        RECT 79.095 136.635 80.025 136.865 ;
        RECT 77.275 135.955 80.025 136.635 ;
        RECT 80.035 135.955 81.850 136.865 ;
        RECT 81.875 135.955 83.245 136.765 ;
        RECT 83.355 135.955 86.465 136.865 ;
        RECT 86.475 136.665 87.420 136.865 ;
        RECT 86.475 135.985 89.225 136.665 ;
        RECT 86.475 135.955 87.420 135.985 ;
        RECT 2.895 135.745 3.065 135.955 ;
        RECT 4.275 135.905 4.445 135.955 ;
        RECT 4.270 135.795 4.445 135.905 ;
        RECT 4.275 135.765 4.445 135.795 ;
        RECT 4.735 135.745 4.905 135.935 ;
        RECT 7.035 135.745 7.205 135.935 ;
        RECT 7.505 135.790 7.665 135.900 ;
        RECT 8.690 135.745 8.860 135.935 ;
        RECT 12.555 135.745 12.725 135.935 ;
        RECT 13.485 135.800 13.645 135.910 ;
        RECT 15.315 135.765 15.485 135.955 ;
        RECT 16.510 135.765 16.680 135.955 ;
        RECT 20.375 135.765 20.545 135.955 ;
        RECT 21.755 135.745 21.925 135.935 ;
        RECT 22.215 135.765 22.385 135.955 ;
        RECT 23.135 135.745 23.305 135.935 ;
        RECT 24.790 135.745 24.960 135.935 ;
        RECT 31.415 135.745 31.585 135.935 ;
        RECT 31.875 135.745 32.045 135.935 ;
        RECT 41.075 135.765 41.245 135.955 ;
        RECT 42.005 135.800 42.165 135.910 ;
        RECT 42.915 135.765 43.085 135.955 ;
        RECT 50.735 135.745 50.905 135.935 ;
        RECT 52.115 135.905 52.285 135.935 ;
        RECT 52.110 135.795 52.285 135.905 ;
        RECT 52.115 135.745 52.285 135.795 ;
        RECT 52.575 135.745 52.745 135.955 ;
        RECT 53.950 135.795 54.070 135.905 ;
        RECT 54.230 135.765 54.400 135.955 ;
        RECT 54.875 135.745 55.045 135.935 ;
        RECT 56.255 135.745 56.425 135.935 ;
        RECT 58.095 135.765 58.265 135.955 ;
        RECT 66.375 135.745 66.545 135.935 ;
        RECT 66.840 135.745 67.010 135.935 ;
        RECT 68.675 135.765 68.845 135.955 ;
        RECT 69.140 135.765 69.310 135.955 ;
        RECT 70.975 135.745 71.145 135.935 ;
        RECT 71.895 135.765 72.065 135.955 ;
        RECT 73.270 135.745 73.440 135.935 ;
        RECT 74.650 135.745 74.820 135.935 ;
        RECT 75.115 135.745 75.285 135.955 ;
        RECT 76.950 135.795 77.070 135.905 ;
        RECT 77.415 135.765 77.585 135.955 ;
        RECT 77.875 135.745 78.045 135.935 ;
        RECT 79.710 135.795 79.830 135.905 ;
        RECT 80.640 135.745 80.810 135.935 ;
        RECT 81.555 135.765 81.725 135.955 ;
        RECT 82.015 135.745 82.185 135.955 ;
        RECT 83.395 135.765 83.565 135.955 ;
        RECT 85.235 135.765 85.405 135.935 ;
        RECT 85.235 135.745 85.400 135.765 ;
        RECT 2.755 134.935 4.125 135.745 ;
        RECT 4.595 134.965 5.965 135.745 ;
        RECT 5.975 134.965 7.345 135.745 ;
        RECT 8.275 135.065 12.175 135.745 ;
        RECT 12.415 135.065 21.605 135.745 ;
        RECT 8.275 134.835 9.205 135.065 ;
        RECT 16.925 134.845 17.855 135.065 ;
        RECT 20.685 134.835 21.605 135.065 ;
        RECT 21.615 134.935 22.985 135.745 ;
        RECT 22.995 134.965 24.365 135.745 ;
        RECT 24.375 135.065 28.275 135.745 ;
        RECT 24.375 134.835 25.305 135.065 ;
        RECT 28.525 134.875 28.955 135.660 ;
        RECT 28.985 135.065 31.725 135.745 ;
        RECT 31.735 135.065 40.925 135.745 ;
        RECT 36.245 134.845 37.175 135.065 ;
        RECT 40.005 134.835 40.925 135.065 ;
        RECT 41.855 135.065 51.045 135.745 ;
        RECT 41.855 134.835 42.775 135.065 ;
        RECT 45.605 134.845 46.535 135.065 ;
        RECT 51.055 134.965 52.425 135.745 ;
        RECT 52.435 134.965 53.805 135.745 ;
        RECT 54.285 134.875 54.715 135.660 ;
        RECT 54.735 134.965 56.105 135.745 ;
        RECT 56.115 135.065 65.305 135.745 ;
        RECT 60.625 134.845 61.555 135.065 ;
        RECT 64.385 134.835 65.305 135.065 ;
        RECT 65.315 134.965 66.685 135.745 ;
        RECT 66.695 135.065 70.825 135.745 ;
        RECT 66.695 134.835 68.035 135.065 ;
        RECT 70.835 134.935 72.205 135.745 ;
        RECT 72.235 134.835 73.585 135.745 ;
        RECT 73.615 134.835 74.965 135.745 ;
        RECT 74.985 134.835 77.715 135.745 ;
        RECT 77.735 135.065 79.565 135.745 ;
        RECT 78.220 134.835 79.565 135.065 ;
        RECT 80.045 134.875 80.475 135.660 ;
        RECT 80.495 134.835 81.845 135.745 ;
        RECT 81.875 134.935 83.245 135.745 ;
        RECT 83.565 135.065 85.400 135.745 ;
        RECT 85.700 135.715 85.870 135.935 ;
        RECT 88.450 135.795 88.570 135.905 ;
        RECT 87.360 135.715 88.305 135.745 ;
        RECT 88.910 135.715 89.080 135.985 ;
        RECT 89.235 135.955 92.155 136.865 ;
        RECT 92.925 136.040 93.355 136.825 ;
        RECT 93.375 135.955 96.125 136.765 ;
        RECT 96.135 136.665 97.080 136.865 ;
        RECT 98.415 136.665 99.345 136.865 ;
        RECT 96.135 136.185 99.345 136.665 ;
        RECT 96.135 135.985 99.205 136.185 ;
        RECT 96.135 135.955 97.080 135.985 ;
        RECT 89.380 135.765 89.550 135.955 ;
        RECT 92.590 135.745 92.760 135.935 ;
        RECT 93.055 135.745 93.225 135.935 ;
        RECT 93.515 135.765 93.685 135.955 ;
        RECT 95.810 135.795 95.930 135.905 ;
        RECT 97.200 135.745 97.370 135.935 ;
        RECT 99.035 135.765 99.205 135.985 ;
        RECT 99.355 135.955 102.105 136.765 ;
        RECT 102.575 136.665 103.520 136.865 ;
        RECT 104.855 136.665 105.785 136.865 ;
        RECT 102.575 136.185 105.785 136.665 ;
        RECT 102.575 135.985 105.645 136.185 ;
        RECT 102.575 135.955 103.520 135.985 ;
        RECT 99.495 135.765 99.665 135.955 ;
        RECT 100.870 135.745 101.040 135.935 ;
        RECT 102.250 135.795 102.370 135.905 ;
        RECT 104.550 135.745 104.720 135.935 ;
        RECT 105.025 135.790 105.185 135.900 ;
        RECT 105.475 135.765 105.645 135.985 ;
        RECT 105.860 135.955 112.030 136.865 ;
        RECT 112.235 136.635 113.185 136.865 ;
        RECT 114.955 136.635 116.330 136.865 ;
        RECT 117.280 136.635 118.650 136.865 ;
        RECT 112.235 136.185 116.330 136.635 ;
        RECT 112.235 135.955 114.945 136.185 ;
        RECT 105.935 135.765 106.105 135.955 ;
        RECT 106.395 135.745 106.565 135.935 ;
        RECT 108.235 135.745 108.405 135.935 ;
        RECT 113.765 135.790 113.925 135.900 ;
        RECT 116.055 135.765 116.225 136.185 ;
        RECT 116.375 135.955 118.650 136.635 ;
        RECT 118.685 136.040 119.115 136.825 ;
        RECT 119.150 135.955 120.965 136.865 ;
        RECT 123.715 136.635 124.645 136.865 ;
        RECT 121.895 135.955 124.645 136.635 ;
        RECT 124.655 136.665 125.600 136.865 ;
        RECT 124.655 135.985 127.405 136.665 ;
        RECT 124.655 135.955 125.600 135.985 ;
        RECT 116.520 135.765 116.690 135.955 ;
        RECT 117.890 135.745 118.060 135.935 ;
        RECT 119.275 135.765 119.445 135.955 ;
        RECT 121.115 135.745 121.285 135.935 ;
        RECT 121.575 135.745 121.745 135.935 ;
        RECT 122.035 135.765 122.205 135.955 ;
        RECT 127.090 135.935 127.260 135.985 ;
        RECT 127.760 135.955 130.165 136.865 ;
        RECT 130.175 135.955 132.005 136.765 ;
        RECT 132.025 135.955 134.755 136.865 ;
        RECT 134.775 136.665 136.185 136.865 ;
        RECT 137.545 136.775 139.135 136.865 ;
        RECT 134.775 135.985 137.510 136.665 ;
        RECT 134.775 135.955 136.170 135.985 ;
        RECT 125.715 135.745 125.885 135.935 ;
        RECT 126.185 135.790 126.345 135.900 ;
        RECT 127.085 135.765 127.260 135.935 ;
        RECT 129.855 135.765 130.025 135.955 ;
        RECT 127.085 135.745 127.255 135.765 ;
        RECT 130.315 135.745 130.485 135.955 ;
        RECT 132.155 135.745 132.325 135.955 ;
        RECT 134.455 135.745 134.625 135.935 ;
        RECT 137.215 135.765 137.385 135.985 ;
        RECT 137.545 135.955 140.115 136.775 ;
        RECT 140.375 135.955 142.585 136.865 ;
        RECT 142.595 135.955 144.425 136.765 ;
        RECT 144.445 136.040 144.875 136.825 ;
        RECT 145.205 136.635 146.135 136.865 ;
        RECT 147.680 136.635 149.025 136.865 ;
        RECT 145.205 135.955 147.040 136.635 ;
        RECT 147.195 135.955 149.025 136.635 ;
        RECT 149.035 135.955 154.545 136.765 ;
        RECT 154.555 135.955 156.385 136.765 ;
        RECT 156.855 135.955 158.225 136.765 ;
        RECT 139.975 135.935 140.115 135.955 ;
        RECT 137.675 135.765 137.845 135.935 ;
        RECT 137.680 135.745 137.845 135.765 ;
        RECT 139.975 135.745 140.145 135.935 ;
        RECT 142.270 135.765 142.440 135.955 ;
        RECT 142.735 135.765 142.905 135.955 ;
        RECT 146.875 135.935 147.040 135.955 ;
        RECT 145.495 135.745 145.665 135.935 ;
        RECT 146.875 135.765 147.045 135.935 ;
        RECT 147.335 135.765 147.505 135.955 ;
        RECT 149.175 135.765 149.345 135.955 ;
        RECT 151.015 135.745 151.185 135.935 ;
        RECT 154.695 135.765 154.865 135.955 ;
        RECT 156.530 135.795 156.650 135.905 ;
        RECT 157.915 135.745 158.085 135.955 ;
        RECT 90.110 135.715 91.065 135.745 ;
        RECT 83.565 134.835 84.495 135.065 ;
        RECT 85.555 135.035 88.305 135.715 ;
        RECT 88.785 135.035 91.065 135.715 ;
        RECT 87.360 134.835 88.305 135.035 ;
        RECT 90.110 134.835 91.065 135.035 ;
        RECT 91.075 134.835 92.905 135.745 ;
        RECT 92.915 134.935 95.665 135.745 ;
        RECT 96.135 134.835 97.485 135.745 ;
        RECT 97.600 135.065 101.185 135.745 ;
        RECT 100.265 134.835 101.185 135.065 ;
        RECT 101.210 134.835 104.865 135.745 ;
        RECT 105.805 134.875 106.235 135.660 ;
        RECT 106.255 134.935 108.085 135.745 ;
        RECT 108.100 134.835 113.410 135.745 ;
        RECT 114.730 134.835 118.205 135.745 ;
        RECT 118.215 134.835 121.425 135.745 ;
        RECT 121.435 134.935 122.805 135.745 ;
        RECT 122.815 134.835 125.925 135.745 ;
        RECT 126.955 134.835 130.165 135.745 ;
        RECT 130.175 134.935 131.545 135.745 ;
        RECT 131.565 134.875 131.995 135.660 ;
        RECT 132.015 135.065 134.305 135.745 ;
        RECT 133.385 134.835 134.305 135.065 ;
        RECT 134.415 134.835 137.525 135.745 ;
        RECT 137.680 135.065 139.515 135.745 ;
        RECT 138.585 134.835 139.515 135.065 ;
        RECT 139.835 134.935 145.345 135.745 ;
        RECT 145.355 134.935 150.865 135.745 ;
        RECT 150.875 134.935 156.385 135.745 ;
        RECT 156.855 134.935 158.225 135.745 ;
      LAYER nwell ;
        RECT 2.560 131.715 158.420 134.545 ;
      LAYER pwell ;
        RECT 2.755 130.515 4.125 131.325 ;
        RECT 4.135 130.515 5.505 131.295 ;
        RECT 10.025 131.195 10.955 131.415 ;
        RECT 13.785 131.195 14.705 131.425 ;
        RECT 5.515 130.515 14.705 131.195 ;
        RECT 15.645 130.600 16.075 131.385 ;
        RECT 16.095 131.195 17.025 131.425 ;
        RECT 16.095 130.515 19.995 131.195 ;
        RECT 21.155 130.515 22.525 131.295 ;
        RECT 27.045 131.195 27.975 131.415 ;
        RECT 30.805 131.195 31.725 131.425 ;
        RECT 34.390 131.195 35.310 131.425 ;
        RECT 22.535 130.515 31.725 131.195 ;
        RECT 31.845 130.515 35.310 131.195 ;
        RECT 35.415 131.195 36.345 131.425 ;
        RECT 35.415 130.515 39.315 131.195 ;
        RECT 40.015 130.515 41.385 131.295 ;
        RECT 41.405 130.600 41.835 131.385 ;
        RECT 41.855 130.515 43.225 131.295 ;
        RECT 46.435 131.195 47.365 131.425 ;
        RECT 43.465 130.515 47.365 131.195 ;
        RECT 47.375 131.225 48.785 131.425 ;
        RECT 47.375 130.545 50.110 131.225 ;
        RECT 50.135 131.195 51.065 131.425 ;
        RECT 54.275 131.195 55.205 131.425 ;
        RECT 47.375 130.515 48.770 130.545 ;
        RECT 2.895 130.305 3.065 130.515 ;
        RECT 4.275 130.305 4.445 130.515 ;
        RECT 5.655 130.325 5.825 130.515 ;
        RECT 7.030 130.355 7.150 130.465 ;
        RECT 8.415 130.305 8.585 130.495 ;
        RECT 8.875 130.305 9.045 130.495 ;
        RECT 10.255 130.305 10.425 130.495 ;
        RECT 14.865 130.360 15.025 130.470 ;
        RECT 16.510 130.325 16.680 130.515 ;
        RECT 19.455 130.305 19.625 130.495 ;
        RECT 20.385 130.360 20.545 130.470 ;
        RECT 22.215 130.325 22.385 130.515 ;
        RECT 22.675 130.325 22.845 130.515 ;
        RECT 29.125 130.350 29.285 130.460 ;
        RECT 30.035 130.305 30.205 130.495 ;
        RECT 31.415 130.305 31.585 130.495 ;
        RECT 31.875 130.325 32.045 130.515 ;
        RECT 35.830 130.325 36.000 130.515 ;
        RECT 39.690 130.355 39.810 130.465 ;
        RECT 40.155 130.325 40.325 130.515 ;
        RECT 40.615 130.305 40.785 130.495 ;
        RECT 41.995 130.325 42.165 130.515 ;
        RECT 46.780 130.325 46.950 130.515 ;
        RECT 49.815 130.325 49.985 130.545 ;
        RECT 50.135 130.515 54.035 131.195 ;
        RECT 54.275 130.515 58.175 131.195 ;
        RECT 58.415 130.515 63.925 131.325 ;
        RECT 63.935 130.515 66.685 131.325 ;
        RECT 67.165 130.600 67.595 131.385 ;
        RECT 68.075 130.515 73.585 131.425 ;
        RECT 73.595 131.225 74.550 131.425 ;
        RECT 73.595 130.545 75.875 131.225 ;
        RECT 73.595 130.515 74.550 130.545 ;
        RECT 50.550 130.325 50.720 130.515 ;
        RECT 53.035 130.305 53.205 130.495 ;
        RECT 53.505 130.350 53.665 130.460 ;
        RECT 54.690 130.325 54.860 130.515 ;
        RECT 54.870 130.355 54.990 130.465 ;
        RECT 55.335 130.305 55.505 130.495 ;
        RECT 56.715 130.305 56.885 130.495 ;
        RECT 58.555 130.325 58.725 130.515 ;
        RECT 64.075 130.325 64.245 130.515 ;
        RECT 65.915 130.305 66.085 130.495 ;
        RECT 66.830 130.355 66.950 130.465 ;
        RECT 67.750 130.355 67.870 130.465 ;
        RECT 68.670 130.355 68.790 130.465 ;
        RECT 73.270 130.325 73.440 130.515 ;
        RECT 74.190 130.305 74.360 130.495 ;
        RECT 75.580 130.325 75.750 130.545 ;
        RECT 75.895 130.515 78.300 131.425 ;
        RECT 78.655 130.515 80.485 131.325 ;
        RECT 80.955 131.195 83.780 131.425 ;
        RECT 80.955 130.515 84.485 131.195 ;
        RECT 84.635 130.515 85.985 131.425 ;
        RECT 86.015 130.515 88.765 131.325 ;
        RECT 88.775 130.515 90.545 131.425 ;
        RECT 90.615 130.515 92.445 131.325 ;
        RECT 92.925 130.600 93.355 131.385 ;
        RECT 93.375 130.515 94.745 131.325 ;
        RECT 94.755 130.515 97.965 131.425 ;
        RECT 97.975 130.515 99.345 131.325 ;
        RECT 99.355 130.515 102.565 131.425 ;
        RECT 102.575 130.515 103.945 131.325 ;
        RECT 103.955 130.515 107.610 131.425 ;
        RECT 107.635 130.515 110.385 131.425 ;
        RECT 112.915 131.335 113.865 131.425 ;
        RECT 110.395 130.515 111.765 131.325 ;
        RECT 111.935 130.515 113.865 131.335 ;
        RECT 114.275 130.515 118.665 131.425 ;
        RECT 118.685 130.600 119.115 131.385 ;
        RECT 119.135 131.225 120.080 131.425 ;
        RECT 121.415 131.225 122.345 131.425 ;
        RECT 119.135 130.745 122.345 131.225 ;
        RECT 119.135 130.545 122.205 130.745 ;
        RECT 119.135 130.515 120.080 130.545 ;
        RECT 76.035 130.325 76.205 130.515 ;
        RECT 77.415 130.305 77.585 130.495 ;
        RECT 77.875 130.305 78.045 130.495 ;
        RECT 78.795 130.325 78.965 130.515 ;
        RECT 84.285 130.495 84.485 130.515 ;
        RECT 85.700 130.495 85.870 130.515 ;
        RECT 79.710 130.355 79.830 130.465 ;
        RECT 80.630 130.355 80.750 130.465 ;
        RECT 83.855 130.305 84.025 130.495 ;
        RECT 84.315 130.305 84.485 130.495 ;
        RECT 85.695 130.325 85.870 130.495 ;
        RECT 86.155 130.325 86.325 130.515 ;
        RECT 87.995 130.325 88.165 130.495 ;
        RECT 88.920 130.325 89.090 130.515 ;
        RECT 90.755 130.325 90.925 130.515 ;
        RECT 85.715 130.305 85.865 130.325 ;
        RECT 88.000 130.305 88.165 130.325 ;
        RECT 91.210 130.305 91.380 130.495 ;
        RECT 92.590 130.355 92.710 130.465 ;
        RECT 93.515 130.325 93.685 130.515 ;
        RECT 93.515 130.305 93.665 130.325 ;
        RECT 93.975 130.305 94.145 130.495 ;
        RECT 94.885 130.325 95.055 130.515 ;
        RECT 98.115 130.325 98.285 130.515 ;
        RECT 99.485 130.325 99.655 130.515 ;
        RECT 102.715 130.325 102.885 130.515 ;
        RECT 104.100 130.305 104.270 130.515 ;
        RECT 105.470 130.355 105.590 130.465 ;
        RECT 106.400 130.305 106.570 130.495 ;
        RECT 107.775 130.325 107.945 130.515 ;
        RECT 110.535 130.325 110.705 130.515 ;
        RECT 111.935 130.495 112.085 130.515 ;
        RECT 111.915 130.325 112.085 130.495 ;
        RECT 111.915 130.305 112.065 130.325 ;
        RECT 112.375 130.305 112.545 130.495 ;
        RECT 115.130 130.355 115.250 130.465 ;
        RECT 115.600 130.305 115.770 130.495 ;
        RECT 118.350 130.325 118.520 130.515 ;
        RECT 118.825 130.350 118.985 130.460 ;
        RECT 121.115 130.305 121.285 130.495 ;
        RECT 122.035 130.325 122.205 130.545 ;
        RECT 122.355 130.515 123.725 131.325 ;
        RECT 123.735 131.195 126.560 131.425 ;
        RECT 123.735 130.515 127.265 131.195 ;
        RECT 127.435 130.515 128.785 131.425 ;
        RECT 128.795 130.515 131.545 131.425 ;
        RECT 131.570 130.515 135.225 131.425 ;
        RECT 135.235 130.515 138.445 131.425 ;
        RECT 138.455 130.515 140.860 131.425 ;
        RECT 141.215 130.515 143.965 131.325 ;
        RECT 144.445 130.600 144.875 131.385 ;
        RECT 144.895 130.515 150.405 131.325 ;
        RECT 150.415 130.515 155.925 131.325 ;
        RECT 156.855 130.515 158.225 131.325 ;
        RECT 122.495 130.325 122.665 130.515 ;
        RECT 127.065 130.495 127.265 130.515 ;
        RECT 124.790 130.305 124.960 130.495 ;
        RECT 125.255 130.305 125.425 130.495 ;
        RECT 127.095 130.325 127.265 130.495 ;
        RECT 128.470 130.325 128.640 130.515 ;
        RECT 128.935 130.305 129.105 130.495 ;
        RECT 130.310 130.305 130.480 130.495 ;
        RECT 131.235 130.325 131.405 130.515 ;
        RECT 132.165 130.350 132.325 130.460 ;
        RECT 134.910 130.325 135.080 130.515 ;
        RECT 138.145 130.325 138.315 130.515 ;
        RECT 138.595 130.305 138.765 130.515 ;
        RECT 139.055 130.305 139.225 130.495 ;
        RECT 140.435 130.305 140.605 130.495 ;
        RECT 141.355 130.325 141.525 130.515 ;
        RECT 144.110 130.355 144.230 130.465 ;
        RECT 145.035 130.325 145.205 130.515 ;
        RECT 145.955 130.305 146.125 130.495 ;
        RECT 150.555 130.325 150.725 130.515 ;
        RECT 151.475 130.305 151.645 130.495 ;
        RECT 156.085 130.360 156.245 130.470 ;
        RECT 157.915 130.305 158.085 130.515 ;
        RECT 2.755 129.495 4.125 130.305 ;
        RECT 4.135 129.495 6.885 130.305 ;
        RECT 7.355 129.525 8.725 130.305 ;
        RECT 8.735 129.495 10.105 130.305 ;
        RECT 10.115 129.625 19.305 130.305 ;
        RECT 19.315 129.625 28.505 130.305 ;
        RECT 14.625 129.405 15.555 129.625 ;
        RECT 18.385 129.395 19.305 129.625 ;
        RECT 23.825 129.405 24.755 129.625 ;
        RECT 27.585 129.395 28.505 129.625 ;
        RECT 28.525 129.435 28.955 130.220 ;
        RECT 29.895 129.525 31.265 130.305 ;
        RECT 31.275 129.625 40.465 130.305 ;
        RECT 40.475 129.625 49.665 130.305 ;
        RECT 35.785 129.405 36.715 129.625 ;
        RECT 39.545 129.395 40.465 129.625 ;
        RECT 44.985 129.405 45.915 129.625 ;
        RECT 48.745 129.395 49.665 129.625 ;
        RECT 49.770 129.625 53.235 130.305 ;
        RECT 49.770 129.395 50.690 129.625 ;
        RECT 54.285 129.435 54.715 130.220 ;
        RECT 55.195 129.525 56.565 130.305 ;
        RECT 56.575 129.625 65.765 130.305 ;
        RECT 61.085 129.405 62.015 129.625 ;
        RECT 64.845 129.395 65.765 129.625 ;
        RECT 65.775 129.495 68.525 130.305 ;
        RECT 68.995 129.395 74.505 130.305 ;
        RECT 74.515 129.395 77.625 130.305 ;
        RECT 77.735 129.495 79.565 130.305 ;
        RECT 80.045 129.435 80.475 130.220 ;
        RECT 80.955 129.395 84.065 130.305 ;
        RECT 84.175 129.495 85.545 130.305 ;
        RECT 85.715 129.485 87.645 130.305 ;
        RECT 88.000 129.625 89.835 130.305 ;
        RECT 86.695 129.395 87.645 129.485 ;
        RECT 88.905 129.395 89.835 129.625 ;
        RECT 90.175 129.395 91.525 130.305 ;
        RECT 91.735 129.485 93.665 130.305 ;
        RECT 91.735 129.395 92.685 129.485 ;
        RECT 93.890 129.395 103.910 130.305 ;
        RECT 103.955 129.395 105.305 130.305 ;
        RECT 105.805 129.435 106.235 130.220 ;
        RECT 106.255 129.395 109.910 130.305 ;
        RECT 110.135 129.485 112.065 130.305 ;
        RECT 112.235 129.495 114.985 130.305 ;
        RECT 110.135 129.395 111.085 129.485 ;
        RECT 115.455 129.395 118.375 130.305 ;
        RECT 119.595 129.395 121.410 130.305 ;
        RECT 121.520 129.625 125.105 130.305 ;
        RECT 124.185 129.395 125.105 129.625 ;
        RECT 125.115 129.495 128.785 130.305 ;
        RECT 128.795 129.495 130.165 130.305 ;
        RECT 130.195 129.395 131.545 130.305 ;
        RECT 131.565 129.435 131.995 130.220 ;
        RECT 133.065 129.395 138.905 130.305 ;
        RECT 138.925 129.395 140.275 130.305 ;
        RECT 140.295 129.495 145.805 130.305 ;
        RECT 145.815 129.495 151.325 130.305 ;
        RECT 151.335 129.495 156.845 130.305 ;
        RECT 156.855 129.495 158.225 130.305 ;
      LAYER nwell ;
        RECT 2.560 126.275 158.420 129.105 ;
      LAYER pwell ;
        RECT 2.755 125.075 4.125 125.885 ;
        RECT 4.135 125.075 7.805 125.885 ;
        RECT 7.815 125.075 9.185 125.885 ;
        RECT 9.195 125.755 10.125 125.985 ;
        RECT 9.195 125.075 13.095 125.755 ;
        RECT 13.795 125.075 15.165 125.855 ;
        RECT 15.645 125.160 16.075 125.945 ;
        RECT 16.095 125.075 18.845 125.885 ;
        RECT 18.950 125.755 19.870 125.985 ;
        RECT 18.950 125.075 22.415 125.755 ;
        RECT 22.535 125.075 28.045 125.885 ;
        RECT 29.070 125.755 29.990 125.985 ;
        RECT 29.070 125.075 32.535 125.755 ;
        RECT 33.575 125.075 34.945 125.855 ;
        RECT 34.955 125.755 35.885 125.985 ;
        RECT 34.955 125.075 38.855 125.755 ;
        RECT 40.015 125.075 41.385 125.855 ;
        RECT 41.405 125.160 41.835 125.945 ;
        RECT 42.315 125.075 43.685 125.855 ;
        RECT 43.695 125.755 44.625 125.985 ;
        RECT 43.695 125.075 47.595 125.755 ;
        RECT 47.835 125.075 49.205 125.885 ;
        RECT 53.725 125.755 54.655 125.975 ;
        RECT 57.485 125.755 58.405 125.985 ;
        RECT 49.215 125.075 58.405 125.755 ;
        RECT 58.415 125.755 59.345 125.985 ;
        RECT 58.415 125.075 62.315 125.755 ;
        RECT 62.555 125.075 66.225 125.885 ;
        RECT 67.165 125.160 67.595 125.945 ;
        RECT 67.615 125.075 73.125 125.985 ;
        RECT 73.135 125.075 74.505 125.885 ;
        RECT 74.515 125.785 75.460 125.985 ;
        RECT 74.515 125.105 77.265 125.785 ;
        RECT 74.515 125.075 75.460 125.105 ;
        RECT 2.895 124.865 3.065 125.075 ;
        RECT 4.275 124.865 4.445 125.075 ;
        RECT 7.955 124.885 8.125 125.075 ;
        RECT 9.610 124.885 9.780 125.075 ;
        RECT 9.795 124.865 9.965 125.055 ;
        RECT 13.470 124.915 13.590 125.025 ;
        RECT 14.855 124.885 15.025 125.075 ;
        RECT 15.315 125.025 15.485 125.055 ;
        RECT 15.310 124.915 15.485 125.025 ;
        RECT 15.315 124.865 15.485 124.915 ;
        RECT 16.235 124.885 16.405 125.075 ;
        RECT 20.835 124.865 21.005 125.055 ;
        RECT 22.215 124.885 22.385 125.075 ;
        RECT 22.675 124.885 22.845 125.075 ;
        RECT 26.355 124.865 26.525 125.055 ;
        RECT 28.205 125.025 28.365 125.030 ;
        RECT 28.190 124.920 28.365 125.025 ;
        RECT 28.190 124.915 28.310 124.920 ;
        RECT 29.115 124.865 29.285 125.055 ;
        RECT 32.335 124.885 32.505 125.075 ;
        RECT 32.805 124.920 32.965 125.030 ;
        RECT 34.635 124.865 34.805 125.075 ;
        RECT 35.370 124.885 35.540 125.075 ;
        RECT 38.310 124.915 38.430 125.025 ;
        RECT 39.245 124.920 39.405 125.030 ;
        RECT 41.075 124.885 41.245 125.075 ;
        RECT 41.995 125.025 42.165 125.055 ;
        RECT 41.990 124.915 42.165 125.025 ;
        RECT 41.995 124.865 42.165 124.915 ;
        RECT 42.455 124.865 42.625 125.055 ;
        RECT 43.375 124.885 43.545 125.075 ;
        RECT 44.110 124.885 44.280 125.075 ;
        RECT 47.975 124.885 48.145 125.075 ;
        RECT 49.355 124.885 49.525 125.075 ;
        RECT 51.195 124.865 51.365 125.055 ;
        RECT 51.655 124.865 51.825 125.055 ;
        RECT 54.875 124.865 55.045 125.055 ;
        RECT 58.830 124.885 59.000 125.075 ;
        RECT 60.395 124.865 60.565 125.055 ;
        RECT 62.695 124.885 62.865 125.075 ;
        RECT 65.915 124.865 66.085 125.055 ;
        RECT 66.385 124.920 66.545 125.030 ;
        RECT 72.810 124.865 72.980 125.075 ;
        RECT 73.275 124.865 73.445 125.075 ;
        RECT 76.950 124.885 77.120 125.105 ;
        RECT 77.275 125.075 80.025 125.985 ;
        RECT 80.035 125.075 82.785 125.885 ;
        RECT 83.265 125.075 85.995 125.985 ;
        RECT 87.820 125.785 88.765 125.985 ;
        RECT 86.015 125.105 88.765 125.785 ;
        RECT 77.415 124.885 77.585 125.075 ;
        RECT 77.870 124.865 78.040 125.055 ;
        RECT 79.260 124.865 79.430 125.055 ;
        RECT 79.710 124.915 79.830 125.025 ;
        RECT 80.175 124.885 80.345 125.075 ;
        RECT 82.930 124.915 83.050 125.025 ;
        RECT 83.395 124.885 83.565 125.075 ;
        RECT 86.160 125.055 86.330 125.105 ;
        RECT 87.820 125.075 88.765 125.105 ;
        RECT 88.975 125.895 89.925 125.985 ;
        RECT 88.975 125.075 90.905 125.895 ;
        RECT 91.075 125.075 92.905 125.885 ;
        RECT 92.925 125.160 93.355 125.945 ;
        RECT 94.745 125.755 95.665 125.985 ;
        RECT 93.375 125.075 95.665 125.755 ;
        RECT 96.135 125.755 97.060 125.985 ;
        RECT 96.135 125.075 99.805 125.755 ;
        RECT 99.815 125.075 101.165 125.985 ;
        RECT 102.115 125.755 103.045 125.985 ;
        RECT 107.485 125.755 108.415 125.985 ;
        RECT 110.245 125.755 111.175 125.985 ;
        RECT 102.115 125.075 106.015 125.755 ;
        RECT 107.485 125.075 109.320 125.755 ;
        RECT 110.245 125.075 112.080 125.755 ;
        RECT 113.155 125.075 116.365 125.985 ;
        RECT 116.685 125.755 117.615 125.985 ;
        RECT 116.685 125.075 118.520 125.755 ;
        RECT 118.685 125.160 119.115 125.945 ;
        RECT 119.155 125.075 120.505 125.985 ;
        RECT 120.515 125.075 121.865 125.985 ;
        RECT 121.895 125.075 125.550 125.985 ;
        RECT 125.575 125.075 128.785 125.985 ;
        RECT 128.795 125.075 131.545 125.885 ;
        RECT 132.015 125.075 134.765 125.985 ;
        RECT 136.110 125.785 137.065 125.985 ;
        RECT 134.785 125.105 137.065 125.785 ;
        RECT 90.755 125.055 90.905 125.075 ;
        RECT 86.155 124.885 86.330 125.055 ;
        RECT 90.750 124.885 90.925 125.055 ;
        RECT 91.215 124.885 91.385 125.075 ;
        RECT 93.515 124.885 93.685 125.075 ;
        RECT 86.155 124.865 86.325 124.885 ;
        RECT 90.750 124.865 90.920 124.885 ;
        RECT 93.975 124.865 94.145 125.055 ;
        RECT 94.425 124.865 94.595 125.055 ;
        RECT 95.810 124.915 95.930 125.025 ;
        RECT 96.280 124.885 96.450 125.075 ;
        RECT 97.650 124.915 97.770 125.025 ;
        RECT 99.035 124.865 99.205 125.055 ;
        RECT 99.495 124.865 99.665 125.055 ;
        RECT 99.960 124.885 100.130 125.075 ;
        RECT 101.345 124.920 101.505 125.030 ;
        RECT 102.530 124.885 102.700 125.075 ;
        RECT 109.155 125.055 109.320 125.075 ;
        RECT 111.915 125.055 112.080 125.075 ;
        RECT 103.175 124.865 103.345 125.055 ;
        RECT 106.405 124.920 106.565 125.030 ;
        RECT 107.775 124.865 107.945 125.055 ;
        RECT 108.230 124.915 108.350 125.025 ;
        RECT 108.700 124.865 108.870 125.055 ;
        RECT 109.155 124.885 109.325 125.055 ;
        RECT 109.610 124.915 109.730 125.025 ;
        RECT 111.915 124.885 112.085 125.055 ;
        RECT 112.385 124.920 112.545 125.030 ;
        RECT 113.295 124.885 113.465 125.075 ;
        RECT 118.355 125.055 118.520 125.075 ;
        RECT 116.515 124.885 116.685 125.055 ;
        RECT 116.485 124.865 116.685 124.885 ;
        RECT 116.980 124.865 117.150 125.055 ;
        RECT 118.355 125.025 118.525 125.055 ;
        RECT 118.350 124.915 118.525 125.025 ;
        RECT 118.355 124.885 118.525 124.915 ;
        RECT 118.815 124.865 118.985 125.055 ;
        RECT 120.190 124.885 120.360 125.075 ;
        RECT 121.580 125.055 121.750 125.075 ;
        RECT 121.575 124.885 121.750 125.055 ;
        RECT 122.040 124.885 122.210 125.075 ;
        RECT 121.575 124.865 121.745 124.885 ;
        RECT 127.560 124.865 127.730 125.055 ;
        RECT 128.485 124.885 128.655 125.075 ;
        RECT 128.935 124.885 129.105 125.075 ;
        RECT 129.855 124.865 130.025 125.055 ;
        RECT 131.690 124.915 131.810 125.025 ;
        RECT 132.155 124.885 132.325 125.075 ;
        RECT 134.910 125.055 135.080 125.105 ;
        RECT 136.110 125.075 137.065 125.105 ;
        RECT 137.075 125.075 142.585 125.885 ;
        RECT 142.595 125.075 144.425 125.885 ;
        RECT 144.445 125.160 144.875 125.945 ;
        RECT 144.895 125.075 150.405 125.885 ;
        RECT 150.415 125.075 155.925 125.885 ;
        RECT 156.855 125.075 158.225 125.885 ;
        RECT 134.910 124.885 135.085 125.055 ;
        RECT 137.215 124.885 137.385 125.075 ;
        RECT 134.915 124.865 135.085 124.885 ;
        RECT 137.675 124.865 137.845 125.055 ;
        RECT 138.135 124.865 138.305 125.055 ;
        RECT 142.735 124.885 142.905 125.075 ;
        RECT 143.655 124.865 143.825 125.055 ;
        RECT 145.035 124.885 145.205 125.075 ;
        RECT 149.175 124.865 149.345 125.055 ;
        RECT 150.555 124.885 150.725 125.075 ;
        RECT 154.695 124.865 154.865 125.055 ;
        RECT 156.085 124.920 156.245 125.030 ;
        RECT 156.530 124.915 156.650 125.025 ;
        RECT 157.915 124.865 158.085 125.075 ;
        RECT 2.755 124.055 4.125 124.865 ;
        RECT 4.135 124.055 9.645 124.865 ;
        RECT 9.655 124.055 15.165 124.865 ;
        RECT 15.175 124.055 20.685 124.865 ;
        RECT 20.695 124.055 26.205 124.865 ;
        RECT 26.215 124.055 28.045 124.865 ;
        RECT 28.525 123.995 28.955 124.780 ;
        RECT 28.975 124.055 34.485 124.865 ;
        RECT 34.495 124.055 38.165 124.865 ;
        RECT 38.730 124.185 42.195 124.865 ;
        RECT 38.730 123.955 39.650 124.185 ;
        RECT 42.315 124.055 47.825 124.865 ;
        RECT 47.930 124.185 51.395 124.865 ;
        RECT 47.930 123.955 48.850 124.185 ;
        RECT 51.515 124.055 54.265 124.865 ;
        RECT 54.285 123.995 54.715 124.780 ;
        RECT 54.735 124.055 60.245 124.865 ;
        RECT 60.255 124.055 65.765 124.865 ;
        RECT 65.775 124.055 67.605 124.865 ;
        RECT 67.615 123.955 73.125 124.865 ;
        RECT 73.135 124.055 74.965 124.865 ;
        RECT 75.265 123.955 78.185 124.865 ;
        RECT 78.195 123.955 79.545 124.865 ;
        RECT 80.045 123.995 80.475 124.780 ;
        RECT 80.625 123.955 86.465 124.865 ;
        RECT 86.475 123.955 91.065 124.865 ;
        RECT 91.075 124.185 94.285 124.865 ;
        RECT 91.075 123.955 92.210 124.185 ;
        RECT 94.295 123.955 97.505 124.865 ;
        RECT 97.985 123.955 99.335 124.865 ;
        RECT 99.355 124.055 103.025 124.865 ;
        RECT 103.045 123.955 105.775 124.865 ;
        RECT 105.805 123.995 106.235 124.780 ;
        RECT 106.255 123.955 108.070 124.865 ;
        RECT 108.555 123.955 112.945 124.865 ;
        RECT 113.155 124.185 116.685 124.865 ;
        RECT 113.155 123.955 115.980 124.185 ;
        RECT 116.835 123.955 118.185 124.865 ;
        RECT 118.685 123.955 121.415 124.865 ;
        RECT 121.435 123.955 127.275 124.865 ;
        RECT 127.415 123.955 128.765 124.865 ;
        RECT 129.730 123.955 131.545 124.865 ;
        RECT 131.565 123.995 131.995 124.780 ;
        RECT 132.015 123.955 135.225 124.865 ;
        RECT 135.235 124.185 137.985 124.865 ;
        RECT 135.235 123.955 136.165 124.185 ;
        RECT 137.995 124.055 143.505 124.865 ;
        RECT 143.515 124.055 149.025 124.865 ;
        RECT 149.035 124.055 154.545 124.865 ;
        RECT 154.555 124.055 156.385 124.865 ;
        RECT 156.855 124.055 158.225 124.865 ;
      LAYER nwell ;
        RECT 2.560 120.835 158.420 123.665 ;
      LAYER pwell ;
        RECT 2.755 119.635 4.125 120.445 ;
        RECT 4.135 119.635 9.645 120.445 ;
        RECT 9.655 119.635 15.165 120.445 ;
        RECT 15.645 119.720 16.075 120.505 ;
        RECT 16.095 119.635 21.605 120.445 ;
        RECT 21.615 119.635 27.125 120.445 ;
        RECT 27.135 119.635 32.645 120.445 ;
        RECT 32.655 119.635 38.165 120.445 ;
        RECT 38.175 119.635 40.925 120.445 ;
        RECT 41.405 119.720 41.835 120.505 ;
        RECT 41.855 119.635 47.365 120.445 ;
        RECT 47.375 119.635 52.885 120.445 ;
        RECT 52.895 119.635 58.405 120.445 ;
        RECT 58.415 119.635 63.925 120.445 ;
        RECT 63.935 119.635 66.685 120.445 ;
        RECT 67.165 119.720 67.595 120.505 ;
        RECT 67.615 119.635 71.285 120.445 ;
        RECT 71.295 119.635 72.665 120.445 ;
        RECT 72.985 120.315 73.915 120.545 ;
        RECT 72.985 119.635 74.820 120.315 ;
        RECT 75.435 119.635 78.605 120.545 ;
        RECT 78.655 119.635 84.165 120.445 ;
        RECT 84.215 119.635 87.385 120.545 ;
        RECT 87.395 119.635 90.145 120.445 ;
        RECT 90.925 120.315 91.855 120.545 ;
        RECT 90.925 119.635 92.760 120.315 ;
        RECT 92.925 119.720 93.355 120.505 ;
        RECT 94.295 120.345 95.240 120.545 ;
        RECT 96.575 120.345 97.505 120.545 ;
        RECT 94.295 119.865 97.505 120.345 ;
        RECT 94.295 119.665 97.365 119.865 ;
        RECT 94.295 119.635 95.240 119.665 ;
        RECT 2.895 119.425 3.065 119.635 ;
        RECT 4.275 119.425 4.445 119.635 ;
        RECT 9.795 119.425 9.965 119.635 ;
        RECT 15.315 119.585 15.485 119.615 ;
        RECT 15.310 119.475 15.485 119.585 ;
        RECT 15.315 119.425 15.485 119.475 ;
        RECT 16.235 119.445 16.405 119.635 ;
        RECT 20.835 119.425 21.005 119.615 ;
        RECT 21.755 119.445 21.925 119.635 ;
        RECT 26.355 119.425 26.525 119.615 ;
        RECT 27.275 119.445 27.445 119.635 ;
        RECT 28.190 119.475 28.310 119.585 ;
        RECT 29.115 119.425 29.285 119.615 ;
        RECT 32.795 119.445 32.965 119.635 ;
        RECT 34.635 119.425 34.805 119.615 ;
        RECT 38.315 119.445 38.485 119.635 ;
        RECT 40.155 119.425 40.325 119.615 ;
        RECT 41.070 119.475 41.190 119.585 ;
        RECT 41.995 119.445 42.165 119.635 ;
        RECT 45.675 119.425 45.845 119.615 ;
        RECT 47.515 119.445 47.685 119.635 ;
        RECT 51.195 119.425 51.365 119.615 ;
        RECT 53.035 119.445 53.205 119.635 ;
        RECT 53.950 119.475 54.070 119.585 ;
        RECT 54.875 119.425 55.045 119.615 ;
        RECT 58.555 119.445 58.725 119.635 ;
        RECT 60.395 119.425 60.565 119.615 ;
        RECT 64.075 119.445 64.245 119.635 ;
        RECT 65.915 119.425 66.085 119.615 ;
        RECT 66.830 119.475 66.950 119.585 ;
        RECT 67.755 119.445 67.925 119.635 ;
        RECT 71.435 119.425 71.605 119.635 ;
        RECT 74.655 119.615 74.820 119.635 ;
        RECT 74.655 119.445 74.825 119.615 ;
        RECT 75.110 119.475 75.230 119.585 ;
        RECT 76.955 119.425 77.125 119.615 ;
        RECT 78.335 119.445 78.505 119.635 ;
        RECT 78.795 119.445 78.965 119.635 ;
        RECT 79.710 119.475 79.830 119.585 ;
        RECT 80.635 119.425 80.805 119.615 ;
        RECT 84.315 119.445 84.485 119.635 ;
        RECT 86.155 119.425 86.325 119.615 ;
        RECT 87.535 119.445 87.705 119.635 ;
        RECT 92.595 119.615 92.760 119.635 ;
        RECT 90.290 119.475 90.410 119.585 ;
        RECT 91.675 119.425 91.845 119.615 ;
        RECT 92.595 119.445 92.765 119.615 ;
        RECT 93.525 119.480 93.685 119.590 ;
        RECT 96.735 119.425 96.905 119.615 ;
        RECT 97.195 119.585 97.365 119.665 ;
        RECT 97.535 119.635 98.885 120.545 ;
        RECT 99.815 119.635 102.985 120.545 ;
        RECT 103.135 119.635 106.245 120.545 ;
        RECT 106.275 119.635 107.625 120.545 ;
        RECT 107.635 119.635 109.005 120.445 ;
        RECT 109.115 119.635 112.225 120.545 ;
        RECT 112.235 119.635 117.745 120.445 ;
        RECT 118.685 119.720 119.115 120.505 ;
        RECT 119.135 119.635 121.885 120.445 ;
        RECT 121.895 119.635 125.065 120.545 ;
        RECT 125.115 119.635 126.465 120.545 ;
        RECT 126.505 119.635 127.855 120.545 ;
        RECT 127.875 119.635 131.545 120.445 ;
        RECT 132.015 119.635 133.845 120.545 ;
        RECT 133.855 119.635 139.365 120.445 ;
        RECT 139.375 119.635 143.045 120.445 ;
        RECT 143.055 119.635 144.425 120.445 ;
        RECT 144.445 119.720 144.875 120.505 ;
        RECT 144.895 119.635 150.405 120.445 ;
        RECT 150.415 119.635 155.925 120.445 ;
        RECT 156.855 119.635 158.225 120.445 ;
        RECT 97.190 119.475 97.365 119.585 ;
        RECT 97.195 119.445 97.365 119.475 ;
        RECT 97.650 119.615 97.820 119.635 ;
        RECT 97.650 119.445 97.830 119.615 ;
        RECT 97.660 119.425 97.830 119.445 ;
        RECT 99.035 119.425 99.205 119.615 ;
        RECT 102.715 119.445 102.885 119.635 ;
        RECT 103.175 119.445 103.345 119.635 ;
        RECT 106.390 119.615 106.560 119.635 ;
        RECT 104.555 119.425 104.725 119.615 ;
        RECT 106.390 119.445 106.565 119.615 ;
        RECT 107.775 119.445 107.945 119.635 ;
        RECT 109.155 119.445 109.325 119.635 ;
        RECT 106.395 119.425 106.565 119.445 ;
        RECT 111.915 119.425 112.085 119.615 ;
        RECT 112.375 119.445 112.545 119.635 ;
        RECT 117.435 119.425 117.605 119.615 ;
        RECT 117.905 119.480 118.065 119.590 ;
        RECT 119.275 119.445 119.445 119.635 ;
        RECT 122.955 119.425 123.125 119.615 ;
        RECT 124.795 119.445 124.965 119.635 ;
        RECT 126.180 119.445 126.350 119.635 ;
        RECT 126.635 119.445 126.805 119.635 ;
        RECT 128.015 119.445 128.185 119.635 ;
        RECT 128.475 119.425 128.645 119.615 ;
        RECT 131.230 119.475 131.350 119.585 ;
        RECT 131.690 119.475 131.810 119.585 ;
        RECT 132.155 119.425 132.325 119.615 ;
        RECT 133.530 119.445 133.700 119.635 ;
        RECT 133.995 119.445 134.165 119.635 ;
        RECT 137.675 119.425 137.845 119.615 ;
        RECT 139.515 119.445 139.685 119.635 ;
        RECT 143.195 119.425 143.365 119.635 ;
        RECT 145.035 119.445 145.205 119.635 ;
        RECT 148.715 119.425 148.885 119.615 ;
        RECT 150.555 119.445 150.725 119.635 ;
        RECT 154.235 119.425 154.405 119.615 ;
        RECT 156.085 119.480 156.245 119.590 ;
        RECT 157.915 119.425 158.085 119.635 ;
        RECT 2.755 118.615 4.125 119.425 ;
        RECT 4.135 118.615 9.645 119.425 ;
        RECT 9.655 118.615 15.165 119.425 ;
        RECT 15.175 118.615 20.685 119.425 ;
        RECT 20.695 118.615 26.205 119.425 ;
        RECT 26.215 118.615 28.045 119.425 ;
        RECT 28.525 118.555 28.955 119.340 ;
        RECT 28.975 118.615 34.485 119.425 ;
        RECT 34.495 118.615 40.005 119.425 ;
        RECT 40.015 118.615 45.525 119.425 ;
        RECT 45.535 118.615 51.045 119.425 ;
        RECT 51.055 118.615 53.805 119.425 ;
        RECT 54.285 118.555 54.715 119.340 ;
        RECT 54.735 118.615 60.245 119.425 ;
        RECT 60.255 118.615 65.765 119.425 ;
        RECT 65.775 118.615 71.285 119.425 ;
        RECT 71.295 118.615 76.805 119.425 ;
        RECT 76.815 118.615 79.565 119.425 ;
        RECT 80.045 118.555 80.475 119.340 ;
        RECT 80.495 118.615 86.005 119.425 ;
        RECT 86.015 118.615 91.525 119.425 ;
        RECT 91.535 118.615 94.285 119.425 ;
        RECT 94.325 118.515 97.045 119.425 ;
        RECT 97.515 118.515 98.865 119.425 ;
        RECT 98.895 118.615 104.405 119.425 ;
        RECT 104.415 118.615 105.785 119.425 ;
        RECT 105.805 118.555 106.235 119.340 ;
        RECT 106.255 118.615 111.765 119.425 ;
        RECT 111.775 118.615 117.285 119.425 ;
        RECT 117.295 118.615 122.805 119.425 ;
        RECT 122.815 118.615 128.325 119.425 ;
        RECT 128.335 118.615 131.085 119.425 ;
        RECT 131.565 118.555 131.995 119.340 ;
        RECT 132.015 118.615 137.525 119.425 ;
        RECT 137.535 118.615 143.045 119.425 ;
        RECT 143.055 118.615 148.565 119.425 ;
        RECT 148.575 118.615 154.085 119.425 ;
        RECT 154.095 118.615 156.845 119.425 ;
        RECT 156.855 118.615 158.225 119.425 ;
      LAYER nwell ;
        RECT 2.560 115.395 158.420 118.225 ;
      LAYER pwell ;
        RECT 2.755 114.195 4.125 115.005 ;
        RECT 4.135 114.195 9.645 115.005 ;
        RECT 9.655 114.195 15.165 115.005 ;
        RECT 15.645 114.280 16.075 115.065 ;
        RECT 16.095 114.195 21.605 115.005 ;
        RECT 21.615 114.195 27.125 115.005 ;
        RECT 27.135 114.195 28.505 115.005 ;
        RECT 28.525 114.280 28.955 115.065 ;
        RECT 28.975 114.195 34.485 115.005 ;
        RECT 34.495 114.195 40.005 115.005 ;
        RECT 40.015 114.195 41.385 115.005 ;
        RECT 41.405 114.280 41.835 115.065 ;
        RECT 41.855 114.195 47.365 115.005 ;
        RECT 47.375 114.195 52.885 115.005 ;
        RECT 52.895 114.195 54.265 115.005 ;
        RECT 54.285 114.280 54.715 115.065 ;
        RECT 54.735 114.195 60.245 115.005 ;
        RECT 60.255 114.195 65.765 115.005 ;
        RECT 65.775 114.195 67.145 115.005 ;
        RECT 67.165 114.280 67.595 115.065 ;
        RECT 67.615 114.195 73.125 115.005 ;
        RECT 73.135 114.195 78.645 115.005 ;
        RECT 78.655 114.195 80.025 115.005 ;
        RECT 80.045 114.280 80.475 115.065 ;
        RECT 80.495 114.195 86.005 115.005 ;
        RECT 86.015 114.195 91.525 115.005 ;
        RECT 91.535 114.195 92.905 115.005 ;
        RECT 92.925 114.280 93.355 115.065 ;
        RECT 93.375 114.195 98.885 115.005 ;
        RECT 98.895 114.195 104.405 115.005 ;
        RECT 104.415 114.195 105.785 115.005 ;
        RECT 105.805 114.280 106.235 115.065 ;
        RECT 106.255 114.195 111.765 115.005 ;
        RECT 111.775 114.195 117.285 115.005 ;
        RECT 117.295 114.195 118.665 115.005 ;
        RECT 118.685 114.280 119.115 115.065 ;
        RECT 119.135 114.195 124.645 115.005 ;
        RECT 124.655 114.195 130.165 115.005 ;
        RECT 130.175 114.195 131.545 115.005 ;
        RECT 131.565 114.280 131.995 115.065 ;
        RECT 132.015 114.195 137.525 115.005 ;
        RECT 137.535 114.195 143.045 115.005 ;
        RECT 143.055 114.195 144.425 115.005 ;
        RECT 144.445 114.280 144.875 115.065 ;
        RECT 144.895 114.195 150.405 115.005 ;
        RECT 150.415 114.195 155.925 115.005 ;
        RECT 156.855 114.195 158.225 115.005 ;
        RECT 2.895 114.005 3.065 114.195 ;
        RECT 4.275 114.005 4.445 114.195 ;
        RECT 9.795 114.005 9.965 114.195 ;
        RECT 15.310 114.035 15.430 114.145 ;
        RECT 16.235 114.005 16.405 114.195 ;
        RECT 21.755 114.005 21.925 114.195 ;
        RECT 27.275 114.005 27.445 114.195 ;
        RECT 29.115 114.005 29.285 114.195 ;
        RECT 34.635 114.005 34.805 114.195 ;
        RECT 40.155 114.005 40.325 114.195 ;
        RECT 41.995 114.005 42.165 114.195 ;
        RECT 47.515 114.005 47.685 114.195 ;
        RECT 53.035 114.005 53.205 114.195 ;
        RECT 54.875 114.005 55.045 114.195 ;
        RECT 60.395 114.005 60.565 114.195 ;
        RECT 65.915 114.005 66.085 114.195 ;
        RECT 67.755 114.005 67.925 114.195 ;
        RECT 73.275 114.005 73.445 114.195 ;
        RECT 78.795 114.005 78.965 114.195 ;
        RECT 80.635 114.005 80.805 114.195 ;
        RECT 86.155 114.005 86.325 114.195 ;
        RECT 91.675 114.005 91.845 114.195 ;
        RECT 93.515 114.005 93.685 114.195 ;
        RECT 99.035 114.005 99.205 114.195 ;
        RECT 104.555 114.005 104.725 114.195 ;
        RECT 106.395 114.005 106.565 114.195 ;
        RECT 111.915 114.005 112.085 114.195 ;
        RECT 117.435 114.005 117.605 114.195 ;
        RECT 119.275 114.005 119.445 114.195 ;
        RECT 124.795 114.005 124.965 114.195 ;
        RECT 130.315 114.005 130.485 114.195 ;
        RECT 132.155 114.005 132.325 114.195 ;
        RECT 137.675 114.005 137.845 114.195 ;
        RECT 143.195 114.005 143.365 114.195 ;
        RECT 145.035 114.005 145.205 114.195 ;
        RECT 150.555 114.005 150.725 114.195 ;
        RECT 156.085 114.040 156.245 114.150 ;
        RECT 157.915 114.005 158.085 114.195 ;
        RECT 105.870 11.460 107.880 55.740 ;
        RECT 109.870 36.760 111.880 82.740 ;
        RECT 112.870 36.760 114.880 82.740 ;
        RECT 115.870 36.760 117.880 82.740 ;
        RECT 118.870 36.760 120.880 82.740 ;
        RECT 121.870 36.760 123.880 82.740 ;
        RECT 124.870 36.760 126.880 82.740 ;
        RECT 127.870 36.760 129.880 82.740 ;
        RECT 130.870 36.760 132.880 82.740 ;
        RECT 103.470 11.060 107.880 11.460 ;
        RECT 105.870 9.760 107.880 11.060 ;
        RECT 109.870 9.760 111.880 35.740 ;
        RECT 112.870 9.760 114.880 35.740 ;
        RECT 115.870 9.760 117.880 35.740 ;
        RECT 118.870 9.760 120.880 35.740 ;
        RECT 121.870 9.760 123.880 35.740 ;
        RECT 124.870 9.760 126.880 35.740 ;
        RECT 127.870 9.760 129.880 35.740 ;
      LAYER li1 ;
        RECT 2.750 220.085 158.230 220.255 ;
        RECT 2.835 218.995 4.045 220.085 ;
        RECT 2.835 218.285 3.355 218.825 ;
        RECT 3.525 218.455 4.045 218.995 ;
        RECT 4.675 219.090 5.025 219.915 ;
        RECT 5.195 219.260 5.525 220.085 ;
        RECT 5.695 219.090 5.865 219.915 ;
        RECT 6.035 219.260 6.290 220.085 ;
        RECT 6.460 219.090 6.705 219.915 ;
        RECT 6.885 219.285 7.170 220.085 ;
        RECT 7.350 219.365 7.680 219.875 ;
        RECT 4.675 219.065 6.705 219.090 ;
        RECT 4.675 218.920 6.745 219.065 ;
        RECT 4.675 218.335 4.905 218.920 ;
        RECT 6.575 218.895 6.745 218.920 ;
        RECT 7.350 218.725 7.600 219.365 ;
        RECT 7.950 219.215 8.120 219.825 ;
        RECT 8.290 219.395 8.620 220.085 ;
        RECT 8.850 219.535 9.090 219.825 ;
        RECT 9.290 219.705 9.710 220.085 ;
        RECT 9.890 219.615 10.520 219.865 ;
        RECT 10.970 219.705 11.300 220.085 ;
        RECT 9.890 219.535 10.060 219.615 ;
        RECT 11.470 219.535 11.640 219.825 ;
        RECT 11.820 219.705 12.200 220.085 ;
        RECT 12.440 219.700 13.270 219.870 ;
        RECT 8.850 219.365 10.060 219.535 ;
        RECT 5.075 218.505 7.600 218.725 ;
        RECT 2.835 217.535 4.045 218.285 ;
        RECT 4.675 218.165 6.705 218.335 ;
        RECT 4.675 217.715 5.025 218.165 ;
        RECT 5.195 217.535 5.525 217.995 ;
        RECT 5.695 217.715 5.865 218.165 ;
        RECT 6.035 217.535 6.290 217.995 ;
        RECT 6.460 217.715 6.705 218.165 ;
        RECT 6.885 217.535 7.170 217.995 ;
        RECT 7.350 217.795 7.600 218.505 ;
        RECT 7.780 219.195 8.120 219.215 ;
        RECT 7.780 219.025 9.720 219.195 ;
        RECT 7.780 218.130 7.990 219.025 ;
        RECT 9.890 218.855 10.060 219.365 ;
        RECT 10.230 219.105 10.750 219.415 ;
        RECT 8.160 218.685 10.060 218.855 ;
        RECT 8.160 218.625 8.490 218.685 ;
        RECT 8.640 218.455 8.970 218.515 ;
        RECT 8.310 218.185 8.970 218.455 ;
        RECT 7.780 217.800 8.120 218.130 ;
        RECT 8.300 217.535 8.960 218.015 ;
        RECT 9.140 217.925 9.310 218.685 ;
        RECT 10.230 218.515 10.410 218.925 ;
        RECT 9.480 218.345 9.810 218.465 ;
        RECT 10.580 218.345 10.750 219.105 ;
        RECT 9.480 218.175 10.750 218.345 ;
        RECT 10.920 219.285 12.270 219.535 ;
        RECT 10.920 218.515 11.090 219.285 ;
        RECT 12.020 219.025 12.270 219.285 ;
        RECT 11.260 218.855 11.510 219.015 ;
        RECT 12.440 218.855 12.610 219.700 ;
        RECT 13.505 219.415 13.675 219.915 ;
        RECT 13.845 219.585 14.175 220.085 ;
        RECT 12.780 219.025 13.280 219.405 ;
        RECT 13.505 219.245 14.200 219.415 ;
        RECT 11.260 218.685 12.610 218.855 ;
        RECT 12.190 218.645 12.610 218.685 ;
        RECT 10.920 218.175 11.320 218.515 ;
        RECT 11.610 218.185 12.020 218.515 ;
        RECT 9.140 217.755 9.990 217.925 ;
        RECT 10.550 217.535 10.890 217.995 ;
        RECT 11.070 217.745 11.320 218.175 ;
        RECT 11.610 217.535 12.020 217.975 ;
        RECT 12.190 217.915 12.360 218.645 ;
        RECT 12.530 218.095 12.880 218.465 ;
        RECT 13.060 218.155 13.280 219.025 ;
        RECT 13.450 218.455 13.860 219.075 ;
        RECT 14.030 218.275 14.200 219.245 ;
        RECT 13.505 218.085 14.200 218.275 ;
        RECT 12.190 217.715 13.205 217.915 ;
        RECT 13.505 217.755 13.675 218.085 ;
        RECT 13.845 217.535 14.175 217.915 ;
        RECT 14.390 217.795 14.615 219.915 ;
        RECT 14.785 219.585 15.115 220.085 ;
        RECT 15.285 219.415 15.455 219.915 ;
        RECT 14.790 219.245 15.455 219.415 ;
        RECT 14.790 218.255 15.020 219.245 ;
        RECT 15.190 218.425 15.540 219.075 ;
        RECT 15.715 218.920 16.005 220.085 ;
        RECT 16.180 218.935 16.440 220.085 ;
        RECT 16.615 219.010 16.870 219.915 ;
        RECT 17.040 219.325 17.370 220.085 ;
        RECT 17.585 219.155 17.755 219.915 ;
        RECT 18.020 219.415 18.275 219.915 ;
        RECT 18.445 219.585 18.775 220.085 ;
        RECT 18.020 219.245 18.770 219.415 ;
        RECT 14.790 218.085 15.455 218.255 ;
        RECT 14.785 217.535 15.115 217.915 ;
        RECT 15.285 217.795 15.455 218.085 ;
        RECT 15.715 217.535 16.005 218.260 ;
        RECT 16.180 217.535 16.440 218.375 ;
        RECT 16.615 218.280 16.785 219.010 ;
        RECT 17.040 218.985 17.755 219.155 ;
        RECT 17.040 218.775 17.210 218.985 ;
        RECT 16.955 218.445 17.210 218.775 ;
        RECT 16.615 217.705 16.870 218.280 ;
        RECT 17.040 218.255 17.210 218.445 ;
        RECT 17.490 218.435 17.845 218.805 ;
        RECT 18.020 218.425 18.370 219.075 ;
        RECT 18.540 218.255 18.770 219.245 ;
        RECT 17.040 218.085 17.755 218.255 ;
        RECT 17.040 217.535 17.370 217.915 ;
        RECT 17.585 217.705 17.755 218.085 ;
        RECT 18.020 218.085 18.770 218.255 ;
        RECT 18.020 217.795 18.275 218.085 ;
        RECT 18.445 217.535 18.775 217.915 ;
        RECT 18.945 217.795 19.115 219.915 ;
        RECT 19.285 219.115 19.610 219.900 ;
        RECT 19.780 219.625 20.030 220.085 ;
        RECT 20.200 219.585 20.450 219.915 ;
        RECT 20.665 219.585 21.345 219.915 ;
        RECT 20.200 219.455 20.370 219.585 ;
        RECT 19.975 219.285 20.370 219.455 ;
        RECT 19.345 218.065 19.805 219.115 ;
        RECT 19.975 217.925 20.145 219.285 ;
        RECT 20.540 219.025 21.005 219.415 ;
        RECT 20.315 218.215 20.665 218.835 ;
        RECT 20.835 218.435 21.005 219.025 ;
        RECT 21.175 218.805 21.345 219.585 ;
        RECT 21.515 219.485 21.685 219.825 ;
        RECT 21.920 219.655 22.250 220.085 ;
        RECT 22.420 219.485 22.590 219.825 ;
        RECT 22.885 219.625 23.255 220.085 ;
        RECT 21.515 219.315 22.590 219.485 ;
        RECT 23.425 219.455 23.595 219.915 ;
        RECT 23.830 219.575 24.700 219.915 ;
        RECT 24.870 219.625 25.120 220.085 ;
        RECT 23.035 219.285 23.595 219.455 ;
        RECT 23.035 219.145 23.205 219.285 ;
        RECT 21.705 218.975 23.205 219.145 ;
        RECT 23.900 219.115 24.360 219.405 ;
        RECT 21.175 218.635 22.865 218.805 ;
        RECT 20.835 218.215 21.190 218.435 ;
        RECT 21.360 217.925 21.530 218.635 ;
        RECT 21.735 218.215 22.525 218.465 ;
        RECT 22.695 218.455 22.865 218.635 ;
        RECT 23.035 218.285 23.205 218.975 ;
        RECT 19.475 217.535 19.805 217.895 ;
        RECT 19.975 217.755 20.470 217.925 ;
        RECT 20.675 217.755 21.530 217.925 ;
        RECT 22.405 217.535 22.735 217.995 ;
        RECT 22.945 217.895 23.205 218.285 ;
        RECT 23.395 219.105 24.360 219.115 ;
        RECT 24.530 219.195 24.700 219.575 ;
        RECT 25.290 219.535 25.460 219.825 ;
        RECT 25.640 219.705 25.970 220.085 ;
        RECT 25.290 219.365 26.090 219.535 ;
        RECT 23.395 218.945 24.070 219.105 ;
        RECT 24.530 219.025 25.750 219.195 ;
        RECT 23.395 218.155 23.605 218.945 ;
        RECT 24.530 218.935 24.700 219.025 ;
        RECT 23.775 218.155 24.125 218.775 ;
        RECT 24.295 218.765 24.700 218.935 ;
        RECT 24.295 217.985 24.465 218.765 ;
        RECT 24.635 218.315 24.855 218.595 ;
        RECT 25.035 218.485 25.575 218.855 ;
        RECT 25.920 218.745 26.090 219.365 ;
        RECT 26.265 219.025 26.435 220.085 ;
        RECT 26.645 219.075 26.935 219.915 ;
        RECT 27.105 219.245 27.275 220.085 ;
        RECT 27.485 219.075 27.735 219.915 ;
        RECT 27.945 219.245 28.115 220.085 ;
        RECT 26.645 218.905 28.370 219.075 ;
        RECT 28.595 218.920 28.885 220.085 ;
        RECT 29.060 218.945 29.395 219.915 ;
        RECT 29.565 218.945 29.735 220.085 ;
        RECT 29.905 219.745 31.935 219.915 ;
        RECT 24.635 218.145 25.165 218.315 ;
        RECT 22.945 217.725 23.295 217.895 ;
        RECT 23.515 217.705 24.465 217.985 ;
        RECT 24.635 217.535 24.825 217.975 ;
        RECT 24.995 217.915 25.165 218.145 ;
        RECT 25.335 218.085 25.575 218.485 ;
        RECT 25.745 218.735 26.090 218.745 ;
        RECT 25.745 218.525 27.775 218.735 ;
        RECT 25.745 218.270 26.070 218.525 ;
        RECT 27.960 218.355 28.370 218.905 ;
        RECT 25.745 217.915 26.065 218.270 ;
        RECT 24.995 217.745 26.065 217.915 ;
        RECT 26.265 217.535 26.435 218.345 ;
        RECT 26.605 218.185 28.370 218.355 ;
        RECT 29.060 218.275 29.230 218.945 ;
        RECT 29.905 218.775 30.075 219.745 ;
        RECT 29.400 218.445 29.655 218.775 ;
        RECT 29.880 218.445 30.075 218.775 ;
        RECT 30.245 219.405 31.370 219.575 ;
        RECT 29.485 218.275 29.655 218.445 ;
        RECT 30.245 218.275 30.415 219.405 ;
        RECT 26.605 217.705 26.935 218.185 ;
        RECT 27.105 217.535 27.275 218.005 ;
        RECT 27.445 217.705 27.775 218.185 ;
        RECT 27.945 217.535 28.115 218.005 ;
        RECT 28.595 217.535 28.885 218.260 ;
        RECT 29.060 217.705 29.315 218.275 ;
        RECT 29.485 218.105 30.415 218.275 ;
        RECT 30.585 219.065 31.595 219.235 ;
        RECT 30.585 218.265 30.755 219.065 ;
        RECT 30.240 218.070 30.415 218.105 ;
        RECT 29.485 217.535 29.815 217.935 ;
        RECT 30.240 217.705 30.770 218.070 ;
        RECT 30.960 218.045 31.235 218.865 ;
        RECT 30.955 217.875 31.235 218.045 ;
        RECT 30.960 217.705 31.235 217.875 ;
        RECT 31.405 217.705 31.595 219.065 ;
        RECT 31.765 219.080 31.935 219.745 ;
        RECT 32.105 219.325 32.275 220.085 ;
        RECT 32.510 219.325 33.025 219.735 ;
        RECT 31.765 218.890 32.515 219.080 ;
        RECT 32.685 218.515 33.025 219.325 ;
        RECT 33.285 219.155 33.455 219.915 ;
        RECT 33.635 219.325 33.965 220.085 ;
        RECT 33.285 218.985 33.950 219.155 ;
        RECT 34.135 219.010 34.405 219.915 ;
        RECT 34.630 219.215 34.915 220.085 ;
        RECT 35.085 219.455 35.345 219.915 ;
        RECT 35.520 219.625 35.775 220.085 ;
        RECT 35.945 219.455 36.205 219.915 ;
        RECT 35.085 219.285 36.205 219.455 ;
        RECT 36.375 219.285 36.685 220.085 ;
        RECT 35.085 219.035 35.345 219.285 ;
        RECT 36.855 219.115 37.165 219.915 ;
        RECT 33.780 218.840 33.950 218.985 ;
        RECT 31.795 218.345 33.025 218.515 ;
        RECT 33.215 218.435 33.545 218.805 ;
        RECT 33.780 218.510 34.065 218.840 ;
        RECT 31.775 217.535 32.285 218.070 ;
        RECT 32.505 217.740 32.750 218.345 ;
        RECT 33.780 218.255 33.950 218.510 ;
        RECT 33.285 218.085 33.950 218.255 ;
        RECT 34.235 218.210 34.405 219.010 ;
        RECT 33.285 217.705 33.455 218.085 ;
        RECT 33.635 217.535 33.965 217.915 ;
        RECT 34.145 217.705 34.405 218.210 ;
        RECT 34.590 218.865 35.345 219.035 ;
        RECT 36.135 218.945 37.165 219.115 ;
        RECT 34.590 218.355 34.995 218.865 ;
        RECT 36.135 218.695 36.305 218.945 ;
        RECT 35.165 218.525 36.305 218.695 ;
        RECT 34.590 218.185 36.240 218.355 ;
        RECT 36.475 218.205 36.825 218.775 ;
        RECT 34.635 217.535 34.915 218.015 ;
        RECT 35.085 217.795 35.345 218.185 ;
        RECT 35.520 217.535 35.775 218.015 ;
        RECT 35.945 217.795 36.240 218.185 ;
        RECT 36.995 218.035 37.165 218.945 ;
        RECT 37.335 219.325 37.850 219.735 ;
        RECT 38.085 219.325 38.255 220.085 ;
        RECT 38.425 219.745 40.455 219.915 ;
        RECT 37.335 218.515 37.675 219.325 ;
        RECT 38.425 219.080 38.595 219.745 ;
        RECT 38.990 219.405 40.115 219.575 ;
        RECT 37.845 218.890 38.595 219.080 ;
        RECT 38.765 219.065 39.775 219.235 ;
        RECT 37.335 218.345 38.565 218.515 ;
        RECT 36.420 217.535 36.695 218.015 ;
        RECT 36.865 217.705 37.165 218.035 ;
        RECT 37.610 217.740 37.855 218.345 ;
        RECT 38.075 217.535 38.585 218.070 ;
        RECT 38.765 217.705 38.955 219.065 ;
        RECT 39.125 218.725 39.400 218.865 ;
        RECT 39.125 218.555 39.405 218.725 ;
        RECT 39.125 217.705 39.400 218.555 ;
        RECT 39.605 218.265 39.775 219.065 ;
        RECT 39.945 218.275 40.115 219.405 ;
        RECT 40.285 218.775 40.455 219.745 ;
        RECT 40.625 218.945 40.795 220.085 ;
        RECT 40.965 218.945 41.300 219.915 ;
        RECT 40.285 218.445 40.480 218.775 ;
        RECT 40.705 218.445 40.960 218.775 ;
        RECT 40.705 218.275 40.875 218.445 ;
        RECT 41.130 218.275 41.300 218.945 ;
        RECT 41.475 218.920 41.765 220.085 ;
        RECT 41.935 219.115 42.245 219.915 ;
        RECT 42.415 219.285 42.725 220.085 ;
        RECT 42.895 219.455 43.155 219.915 ;
        RECT 43.325 219.625 43.580 220.085 ;
        RECT 43.755 219.455 44.015 219.915 ;
        RECT 42.895 219.285 44.015 219.455 ;
        RECT 41.935 218.945 42.965 219.115 ;
        RECT 39.945 218.105 40.875 218.275 ;
        RECT 39.945 218.070 40.120 218.105 ;
        RECT 39.590 217.705 40.120 218.070 ;
        RECT 40.545 217.535 40.875 217.935 ;
        RECT 41.045 217.705 41.300 218.275 ;
        RECT 41.475 217.535 41.765 218.260 ;
        RECT 41.935 218.035 42.105 218.945 ;
        RECT 42.275 218.205 42.625 218.775 ;
        RECT 42.795 218.695 42.965 218.945 ;
        RECT 43.755 219.035 44.015 219.285 ;
        RECT 44.185 219.215 44.470 220.085 ;
        RECT 43.755 218.865 44.510 219.035 ;
        RECT 42.795 218.525 43.935 218.695 ;
        RECT 44.105 218.355 44.510 218.865 ;
        RECT 42.860 218.185 44.510 218.355 ;
        RECT 44.695 219.010 44.965 219.915 ;
        RECT 45.135 219.325 45.465 220.085 ;
        RECT 45.645 219.155 45.815 219.915 ;
        RECT 44.695 218.210 44.865 219.010 ;
        RECT 45.150 218.985 45.815 219.155 ;
        RECT 46.075 219.325 46.590 219.735 ;
        RECT 46.825 219.325 46.995 220.085 ;
        RECT 47.165 219.745 49.195 219.915 ;
        RECT 45.150 218.840 45.320 218.985 ;
        RECT 45.035 218.510 45.320 218.840 ;
        RECT 45.150 218.255 45.320 218.510 ;
        RECT 45.555 218.435 45.885 218.805 ;
        RECT 46.075 218.515 46.415 219.325 ;
        RECT 47.165 219.080 47.335 219.745 ;
        RECT 47.730 219.405 48.855 219.575 ;
        RECT 46.585 218.890 47.335 219.080 ;
        RECT 47.505 219.065 48.515 219.235 ;
        RECT 46.075 218.345 47.305 218.515 ;
        RECT 41.935 217.705 42.235 218.035 ;
        RECT 42.405 217.535 42.680 218.015 ;
        RECT 42.860 217.795 43.155 218.185 ;
        RECT 43.325 217.535 43.580 218.015 ;
        RECT 43.755 217.795 44.015 218.185 ;
        RECT 44.185 217.535 44.465 218.015 ;
        RECT 44.695 217.705 44.955 218.210 ;
        RECT 45.150 218.085 45.815 218.255 ;
        RECT 45.135 217.535 45.465 217.915 ;
        RECT 45.645 217.705 45.815 218.085 ;
        RECT 46.350 217.740 46.595 218.345 ;
        RECT 46.815 217.535 47.325 218.070 ;
        RECT 47.505 217.705 47.695 219.065 ;
        RECT 47.865 218.045 48.140 218.865 ;
        RECT 48.345 218.265 48.515 219.065 ;
        RECT 48.685 218.275 48.855 219.405 ;
        RECT 49.025 218.775 49.195 219.745 ;
        RECT 49.365 218.945 49.535 220.085 ;
        RECT 49.705 218.945 50.040 219.915 ;
        RECT 49.025 218.445 49.220 218.775 ;
        RECT 49.445 218.445 49.700 218.775 ;
        RECT 49.445 218.275 49.615 218.445 ;
        RECT 49.870 218.275 50.040 218.945 ;
        RECT 48.685 218.105 49.615 218.275 ;
        RECT 48.685 218.070 48.860 218.105 ;
        RECT 47.865 217.875 48.145 218.045 ;
        RECT 47.865 217.705 48.140 217.875 ;
        RECT 48.330 217.705 48.860 218.070 ;
        RECT 49.285 217.535 49.615 217.935 ;
        RECT 49.785 217.705 50.040 218.275 ;
        RECT 50.215 219.115 50.525 219.915 ;
        RECT 50.695 219.285 51.005 220.085 ;
        RECT 51.175 219.455 51.435 219.915 ;
        RECT 51.605 219.625 51.860 220.085 ;
        RECT 52.035 219.455 52.295 219.915 ;
        RECT 51.175 219.285 52.295 219.455 ;
        RECT 50.215 218.945 51.245 219.115 ;
        RECT 50.215 218.035 50.385 218.945 ;
        RECT 50.555 218.205 50.905 218.775 ;
        RECT 51.075 218.695 51.245 218.945 ;
        RECT 52.035 219.035 52.295 219.285 ;
        RECT 52.465 219.215 52.750 220.085 ;
        RECT 52.035 218.865 52.790 219.035 ;
        RECT 52.975 218.995 54.185 220.085 ;
        RECT 51.075 218.525 52.215 218.695 ;
        RECT 52.385 218.355 52.790 218.865 ;
        RECT 51.140 218.185 52.790 218.355 ;
        RECT 52.975 218.285 53.495 218.825 ;
        RECT 53.665 218.455 54.185 218.995 ;
        RECT 54.355 218.920 54.645 220.085 ;
        RECT 55.330 219.215 55.615 220.085 ;
        RECT 55.785 219.455 56.045 219.915 ;
        RECT 56.220 219.625 56.475 220.085 ;
        RECT 56.645 219.455 56.905 219.915 ;
        RECT 55.785 219.285 56.905 219.455 ;
        RECT 57.075 219.285 57.385 220.085 ;
        RECT 55.785 219.035 56.045 219.285 ;
        RECT 57.555 219.115 57.865 219.915 ;
        RECT 55.290 218.865 56.045 219.035 ;
        RECT 56.835 218.945 57.865 219.115 ;
        RECT 55.290 218.355 55.695 218.865 ;
        RECT 56.835 218.695 57.005 218.945 ;
        RECT 55.865 218.525 57.005 218.695 ;
        RECT 50.215 217.705 50.515 218.035 ;
        RECT 50.685 217.535 50.960 218.015 ;
        RECT 51.140 217.795 51.435 218.185 ;
        RECT 51.605 217.535 51.860 218.015 ;
        RECT 52.035 217.795 52.295 218.185 ;
        RECT 52.465 217.535 52.745 218.015 ;
        RECT 52.975 217.535 54.185 218.285 ;
        RECT 54.355 217.535 54.645 218.260 ;
        RECT 55.290 218.185 56.940 218.355 ;
        RECT 57.175 218.205 57.525 218.775 ;
        RECT 55.335 217.535 55.615 218.015 ;
        RECT 55.785 217.795 56.045 218.185 ;
        RECT 56.220 217.535 56.475 218.015 ;
        RECT 56.645 217.795 56.940 218.185 ;
        RECT 57.695 218.035 57.865 218.945 ;
        RECT 57.120 217.535 57.395 218.015 ;
        RECT 57.565 217.705 57.865 218.035 ;
        RECT 58.955 219.115 59.265 219.915 ;
        RECT 59.435 219.285 59.745 220.085 ;
        RECT 59.915 219.455 60.175 219.915 ;
        RECT 60.345 219.625 60.600 220.085 ;
        RECT 60.775 219.455 61.035 219.915 ;
        RECT 59.915 219.285 61.035 219.455 ;
        RECT 58.955 218.945 59.985 219.115 ;
        RECT 58.955 218.035 59.125 218.945 ;
        RECT 59.295 218.205 59.645 218.775 ;
        RECT 59.815 218.695 59.985 218.945 ;
        RECT 60.775 219.035 61.035 219.285 ;
        RECT 61.205 219.215 61.490 220.085 ;
        RECT 61.715 219.115 62.025 219.915 ;
        RECT 62.195 219.285 62.505 220.085 ;
        RECT 62.675 219.455 62.935 219.915 ;
        RECT 63.105 219.625 63.360 220.085 ;
        RECT 63.535 219.455 63.795 219.915 ;
        RECT 62.675 219.285 63.795 219.455 ;
        RECT 60.775 218.865 61.530 219.035 ;
        RECT 59.815 218.525 60.955 218.695 ;
        RECT 61.125 218.355 61.530 218.865 ;
        RECT 59.880 218.185 61.530 218.355 ;
        RECT 61.715 218.945 62.745 219.115 ;
        RECT 58.955 217.705 59.255 218.035 ;
        RECT 59.425 217.535 59.700 218.015 ;
        RECT 59.880 217.795 60.175 218.185 ;
        RECT 60.345 217.535 60.600 218.015 ;
        RECT 60.775 217.795 61.035 218.185 ;
        RECT 61.715 218.035 61.885 218.945 ;
        RECT 62.055 218.205 62.405 218.775 ;
        RECT 62.575 218.695 62.745 218.945 ;
        RECT 63.535 219.035 63.795 219.285 ;
        RECT 63.965 219.215 64.250 220.085 ;
        RECT 64.510 219.295 65.045 219.915 ;
        RECT 63.535 218.865 64.290 219.035 ;
        RECT 62.575 218.525 63.715 218.695 ;
        RECT 63.885 218.355 64.290 218.865 ;
        RECT 62.640 218.185 64.290 218.355 ;
        RECT 64.510 218.275 64.825 219.295 ;
        RECT 65.215 219.285 65.545 220.085 ;
        RECT 66.030 219.115 66.420 219.290 ;
        RECT 64.995 218.945 66.420 219.115 ;
        RECT 64.995 218.445 65.165 218.945 ;
        RECT 61.205 217.535 61.485 218.015 ;
        RECT 61.715 217.705 62.015 218.035 ;
        RECT 62.185 217.535 62.460 218.015 ;
        RECT 62.640 217.795 62.935 218.185 ;
        RECT 63.105 217.535 63.360 218.015 ;
        RECT 63.535 217.795 63.795 218.185 ;
        RECT 63.965 217.535 64.245 218.015 ;
        RECT 64.510 217.705 65.125 218.275 ;
        RECT 65.415 218.215 65.680 218.775 ;
        RECT 65.850 218.045 66.020 218.945 ;
        RECT 67.235 218.920 67.525 220.085 ;
        RECT 67.700 219.705 68.035 220.085 ;
        RECT 66.190 218.215 66.545 218.775 ;
        RECT 65.295 217.535 65.510 218.045 ;
        RECT 65.740 217.715 66.020 218.045 ;
        RECT 66.200 217.535 66.440 218.045 ;
        RECT 67.235 217.535 67.525 218.260 ;
        RECT 67.695 218.215 67.935 219.525 ;
        RECT 68.205 219.115 68.455 219.915 ;
        RECT 68.675 219.365 69.005 220.085 ;
        RECT 69.190 219.115 69.440 219.915 ;
        RECT 69.905 219.285 70.235 220.085 ;
        RECT 70.405 219.655 70.745 219.915 ;
        RECT 68.105 218.945 70.295 219.115 ;
        RECT 68.105 218.035 68.275 218.945 ;
        RECT 69.980 218.775 70.295 218.945 ;
        RECT 67.780 217.705 68.275 218.035 ;
        RECT 68.495 217.810 68.845 218.775 ;
        RECT 69.025 217.805 69.325 218.775 ;
        RECT 69.505 217.805 69.785 218.775 ;
        RECT 69.980 218.525 70.310 218.775 ;
        RECT 69.965 217.535 70.235 218.335 ;
        RECT 70.485 218.255 70.745 219.655 ;
        RECT 70.405 217.745 70.745 218.255 ;
        RECT 70.915 219.215 71.190 219.915 ;
        RECT 71.360 219.540 71.615 220.085 ;
        RECT 71.785 219.575 72.265 219.915 ;
        RECT 72.440 219.530 73.045 220.085 ;
        RECT 72.430 219.430 73.045 219.530 ;
        RECT 72.430 219.405 72.615 219.430 ;
        RECT 70.915 218.185 71.085 219.215 ;
        RECT 71.360 219.085 72.115 219.335 ;
        RECT 72.285 219.160 72.615 219.405 ;
        RECT 71.360 219.050 72.130 219.085 ;
        RECT 71.360 219.040 72.145 219.050 ;
        RECT 71.255 219.025 72.150 219.040 ;
        RECT 71.255 219.010 72.170 219.025 ;
        RECT 71.255 219.000 72.190 219.010 ;
        RECT 71.255 218.990 72.215 219.000 ;
        RECT 71.255 218.960 72.285 218.990 ;
        RECT 71.255 218.930 72.305 218.960 ;
        RECT 71.255 218.900 72.325 218.930 ;
        RECT 71.255 218.875 72.355 218.900 ;
        RECT 71.255 218.840 72.390 218.875 ;
        RECT 71.255 218.835 72.420 218.840 ;
        RECT 71.255 218.440 71.485 218.835 ;
        RECT 72.030 218.830 72.420 218.835 ;
        RECT 72.055 218.820 72.420 218.830 ;
        RECT 72.070 218.815 72.420 218.820 ;
        RECT 72.085 218.810 72.420 218.815 ;
        RECT 72.785 218.810 73.045 219.260 ;
        RECT 73.305 219.155 73.475 219.915 ;
        RECT 73.690 219.325 74.020 220.085 ;
        RECT 73.305 218.985 74.020 219.155 ;
        RECT 74.190 219.010 74.445 219.915 ;
        RECT 72.085 218.805 73.045 218.810 ;
        RECT 72.095 218.795 73.045 218.805 ;
        RECT 72.105 218.790 73.045 218.795 ;
        RECT 72.115 218.780 73.045 218.790 ;
        RECT 72.120 218.770 73.045 218.780 ;
        RECT 72.125 218.765 73.045 218.770 ;
        RECT 72.135 218.750 73.045 218.765 ;
        RECT 72.140 218.735 73.045 218.750 ;
        RECT 72.150 218.710 73.045 218.735 ;
        RECT 71.655 218.240 71.985 218.665 ;
        RECT 70.915 217.705 71.175 218.185 ;
        RECT 71.345 217.535 71.595 218.075 ;
        RECT 71.765 217.755 71.985 218.240 ;
        RECT 72.155 218.640 73.045 218.710 ;
        RECT 72.155 217.915 72.325 218.640 ;
        RECT 72.495 218.085 73.045 218.470 ;
        RECT 73.215 218.435 73.570 218.805 ;
        RECT 73.850 218.775 74.020 218.985 ;
        RECT 73.850 218.445 74.105 218.775 ;
        RECT 73.850 218.255 74.020 218.445 ;
        RECT 74.275 218.280 74.445 219.010 ;
        RECT 74.620 218.935 74.880 220.085 ;
        RECT 75.055 218.995 78.565 220.085 ;
        RECT 78.735 218.995 79.945 220.085 ;
        RECT 73.305 218.085 74.020 218.255 ;
        RECT 72.155 217.745 73.045 217.915 ;
        RECT 73.305 217.705 73.475 218.085 ;
        RECT 73.690 217.535 74.020 217.915 ;
        RECT 74.190 217.705 74.445 218.280 ;
        RECT 74.620 217.535 74.880 218.375 ;
        RECT 75.055 218.305 76.705 218.825 ;
        RECT 76.875 218.475 78.565 218.995 ;
        RECT 75.055 217.535 78.565 218.305 ;
        RECT 78.735 218.285 79.255 218.825 ;
        RECT 79.425 218.455 79.945 218.995 ;
        RECT 80.115 218.920 80.405 220.085 ;
        RECT 80.575 218.995 82.245 220.085 ;
        RECT 80.575 218.305 81.325 218.825 ;
        RECT 81.495 218.475 82.245 218.995 ;
        RECT 82.415 218.945 82.675 220.085 ;
        RECT 82.915 219.575 84.530 219.905 ;
        RECT 82.925 218.775 83.095 219.335 ;
        RECT 83.355 219.235 84.530 219.405 ;
        RECT 84.700 219.285 84.980 220.085 ;
        RECT 83.355 218.945 83.685 219.235 ;
        RECT 84.360 219.115 84.530 219.235 ;
        RECT 83.855 218.775 84.100 219.065 ;
        RECT 84.360 218.945 85.020 219.115 ;
        RECT 85.190 218.945 85.465 219.915 ;
        RECT 85.635 219.650 90.980 220.085 ;
        RECT 84.850 218.775 85.020 218.945 ;
        RECT 82.420 218.525 82.755 218.775 ;
        RECT 82.925 218.445 83.640 218.775 ;
        RECT 83.855 218.445 84.680 218.775 ;
        RECT 84.850 218.445 85.125 218.775 ;
        RECT 82.925 218.355 83.175 218.445 ;
        RECT 78.735 217.535 79.945 218.285 ;
        RECT 80.115 217.535 80.405 218.260 ;
        RECT 80.575 217.535 82.245 218.305 ;
        RECT 82.415 217.535 82.675 218.355 ;
        RECT 82.845 217.935 83.175 218.355 ;
        RECT 84.850 218.275 85.020 218.445 ;
        RECT 83.355 218.105 85.020 218.275 ;
        RECT 85.295 218.210 85.465 218.945 ;
        RECT 83.355 217.705 83.615 218.105 ;
        RECT 83.785 217.535 84.115 217.935 ;
        RECT 84.285 217.755 84.455 218.105 ;
        RECT 84.625 217.535 85.000 217.935 ;
        RECT 85.190 217.865 85.465 218.210 ;
        RECT 87.220 218.080 87.560 218.910 ;
        RECT 89.040 218.400 89.390 219.650 ;
        RECT 91.155 218.995 92.825 220.085 ;
        RECT 91.155 218.305 91.905 218.825 ;
        RECT 92.075 218.475 92.825 218.995 ;
        RECT 92.995 218.920 93.285 220.085 ;
        RECT 93.455 218.520 93.805 219.915 ;
        RECT 93.975 219.285 94.380 220.085 ;
        RECT 94.550 219.745 96.085 219.915 ;
        RECT 94.550 219.115 94.720 219.745 ;
        RECT 93.975 218.945 94.720 219.115 ;
        RECT 85.635 217.535 90.980 218.080 ;
        RECT 91.155 217.535 92.825 218.305 ;
        RECT 92.995 217.535 93.285 218.260 ;
        RECT 93.455 217.705 93.725 218.520 ;
        RECT 93.975 218.445 94.145 218.945 ;
        RECT 94.890 218.775 95.160 219.520 ;
        RECT 94.315 218.445 94.650 218.775 ;
        RECT 94.820 218.445 95.160 218.775 ;
        RECT 95.350 218.775 95.585 219.520 ;
        RECT 95.755 219.115 96.085 219.745 ;
        RECT 96.270 219.285 96.505 220.085 ;
        RECT 96.675 219.115 96.965 219.915 ;
        RECT 95.755 218.945 96.965 219.115 ;
        RECT 97.135 218.995 100.645 220.085 ;
        RECT 101.840 219.285 102.095 220.085 ;
        RECT 102.265 219.115 102.595 219.915 ;
        RECT 102.765 219.285 102.935 220.085 ;
        RECT 103.105 219.115 103.435 219.915 ;
        RECT 95.350 218.445 95.640 218.775 ;
        RECT 95.810 218.445 96.210 218.775 ;
        RECT 96.380 218.275 96.550 218.945 ;
        RECT 96.720 218.445 96.965 218.775 ;
        RECT 97.135 218.305 98.785 218.825 ;
        RECT 98.955 218.475 100.645 218.995 ;
        RECT 101.735 218.945 103.435 219.115 ;
        RECT 103.605 218.945 103.865 220.085 ;
        RECT 104.035 218.995 105.705 220.085 ;
        RECT 101.735 218.355 102.015 218.945 ;
        RECT 102.185 218.525 102.935 218.775 ;
        RECT 103.105 218.525 103.865 218.775 ;
        RECT 93.895 217.535 94.565 218.275 ;
        RECT 94.735 218.105 96.130 218.275 ;
        RECT 94.735 217.760 95.030 218.105 ;
        RECT 95.210 217.535 95.585 217.935 ;
        RECT 95.800 217.760 96.130 218.105 ;
        RECT 96.380 217.705 96.965 218.275 ;
        RECT 97.135 217.535 100.645 218.305 ;
        RECT 101.735 218.105 102.595 218.355 ;
        RECT 102.765 218.165 103.865 218.335 ;
        RECT 101.845 217.915 102.175 217.935 ;
        RECT 102.765 217.915 103.015 218.165 ;
        RECT 101.845 217.705 103.015 217.915 ;
        RECT 103.185 217.535 103.355 217.995 ;
        RECT 103.525 217.705 103.865 218.165 ;
        RECT 104.035 218.305 104.785 218.825 ;
        RECT 104.955 218.475 105.705 218.995 ;
        RECT 105.875 218.920 106.165 220.085 ;
        RECT 106.815 219.030 107.120 219.815 ;
        RECT 107.300 219.615 107.985 220.085 ;
        RECT 107.295 219.095 107.990 219.405 ;
        RECT 104.035 217.535 105.705 218.305 ;
        RECT 105.875 217.535 106.165 218.260 ;
        RECT 106.815 218.225 106.990 219.030 ;
        RECT 108.165 218.925 108.450 219.870 ;
        RECT 108.625 219.635 108.955 220.085 ;
        RECT 109.125 219.465 109.295 219.895 ;
        RECT 109.555 219.650 114.900 220.085 ;
        RECT 107.590 218.775 108.450 218.925 ;
        RECT 107.165 218.755 108.450 218.775 ;
        RECT 108.620 219.235 109.295 219.465 ;
        RECT 107.165 218.395 108.150 218.755 ;
        RECT 108.620 218.585 108.855 219.235 ;
        RECT 106.815 217.705 107.055 218.225 ;
        RECT 107.980 218.060 108.150 218.395 ;
        RECT 108.320 218.255 108.855 218.585 ;
        RECT 108.635 218.105 108.855 218.255 ;
        RECT 109.025 218.215 109.325 219.065 ;
        RECT 107.225 217.535 107.620 218.030 ;
        RECT 107.980 217.865 108.355 218.060 ;
        RECT 108.185 217.720 108.355 217.865 ;
        RECT 108.635 217.730 108.875 218.105 ;
        RECT 111.140 218.080 111.480 218.910 ;
        RECT 112.960 218.400 113.310 219.650 ;
        RECT 115.075 218.995 118.585 220.085 ;
        RECT 115.075 218.305 116.725 218.825 ;
        RECT 116.895 218.475 118.585 218.995 ;
        RECT 118.755 218.920 119.045 220.085 ;
        RECT 119.265 219.625 119.515 220.085 ;
        RECT 119.725 219.455 119.895 219.915 ;
        RECT 119.220 219.285 119.895 219.455 ;
        RECT 120.065 219.285 120.315 220.085 ;
        RECT 120.485 219.455 120.735 219.875 ;
        RECT 120.945 219.625 121.275 220.085 ;
        RECT 121.465 219.455 121.715 219.875 ;
        RECT 120.485 219.285 121.775 219.455 ;
        RECT 119.220 218.335 119.475 219.285 ;
        RECT 122.005 219.115 122.175 219.915 ;
        RECT 119.685 218.945 122.175 219.115 ;
        RECT 122.435 219.010 122.705 219.915 ;
        RECT 122.875 219.325 123.205 220.085 ;
        RECT 123.385 219.155 123.555 219.915 ;
        RECT 119.685 218.695 119.855 218.945 ;
        RECT 119.685 218.525 120.015 218.695 ;
        RECT 120.195 218.445 120.525 218.775 ;
        RECT 120.755 218.695 120.925 218.710 ;
        RECT 120.755 218.525 121.085 218.695 ;
        RECT 109.045 217.535 109.380 218.040 ;
        RECT 109.555 217.535 114.900 218.080 ;
        RECT 115.075 217.535 118.585 218.305 ;
        RECT 118.755 217.535 119.045 218.260 ;
        RECT 119.220 218.165 119.895 218.335 ;
        RECT 120.195 218.210 120.400 218.445 ;
        RECT 120.755 218.315 120.925 218.525 ;
        RECT 121.315 218.320 121.485 218.775 ;
        RECT 119.725 218.045 119.895 218.165 ;
        RECT 120.660 218.145 120.925 218.315 ;
        RECT 121.095 218.150 121.485 218.320 ;
        RECT 120.660 218.045 120.830 218.145 ;
        RECT 119.220 217.535 119.475 217.995 ;
        RECT 119.725 217.875 119.905 218.045 ;
        RECT 120.145 217.915 120.315 217.995 ;
        RECT 119.725 217.705 119.895 217.875 ;
        RECT 120.085 217.535 120.415 217.915 ;
        RECT 120.655 217.875 120.830 218.045 ;
        RECT 120.660 217.850 120.830 217.875 ;
        RECT 121.095 217.865 121.305 218.150 ;
        RECT 121.665 217.955 121.835 218.945 ;
        RECT 122.025 218.205 122.220 218.775 ;
        RECT 122.435 218.210 122.605 219.010 ;
        RECT 122.890 218.985 123.555 219.155 ;
        RECT 123.815 218.995 126.405 220.085 ;
        RECT 122.890 218.840 123.060 218.985 ;
        RECT 122.775 218.510 123.060 218.840 ;
        RECT 122.890 218.255 123.060 218.510 ;
        RECT 123.295 218.435 123.625 218.805 ;
        RECT 123.815 218.305 125.025 218.825 ;
        RECT 125.195 218.475 126.405 218.995 ;
        RECT 126.595 219.030 126.900 219.815 ;
        RECT 127.080 219.615 127.765 220.085 ;
        RECT 127.075 219.095 127.770 219.405 ;
        RECT 121.505 217.785 121.835 217.955 ;
        RECT 121.590 217.705 121.835 217.785 ;
        RECT 122.005 217.535 122.265 218.015 ;
        RECT 122.435 217.705 122.695 218.210 ;
        RECT 122.890 218.085 123.555 218.255 ;
        RECT 122.875 217.535 123.205 217.915 ;
        RECT 123.385 217.705 123.555 218.085 ;
        RECT 123.815 217.535 126.405 218.305 ;
        RECT 126.595 218.225 126.770 219.030 ;
        RECT 127.945 218.925 128.230 219.870 ;
        RECT 128.405 219.635 128.735 220.085 ;
        RECT 128.905 219.465 129.075 219.895 ;
        RECT 127.370 218.775 128.230 218.925 ;
        RECT 126.945 218.755 128.230 218.775 ;
        RECT 128.400 219.235 129.075 219.465 ;
        RECT 126.945 218.395 127.930 218.755 ;
        RECT 128.400 218.585 128.635 219.235 ;
        RECT 126.595 217.705 126.835 218.225 ;
        RECT 127.760 218.060 127.930 218.395 ;
        RECT 128.100 218.255 128.635 218.585 ;
        RECT 128.415 218.105 128.635 218.255 ;
        RECT 128.805 218.215 129.105 219.065 ;
        RECT 129.335 219.010 129.605 219.915 ;
        RECT 129.775 219.325 130.105 220.085 ;
        RECT 130.285 219.155 130.455 219.915 ;
        RECT 129.335 218.210 129.505 219.010 ;
        RECT 129.790 218.985 130.455 219.155 ;
        RECT 129.790 218.840 129.960 218.985 ;
        RECT 131.635 218.920 131.925 220.085 ;
        RECT 132.095 219.010 132.365 219.915 ;
        RECT 132.535 219.325 132.865 220.085 ;
        RECT 133.045 219.155 133.215 219.915 ;
        RECT 129.675 218.510 129.960 218.840 ;
        RECT 129.790 218.255 129.960 218.510 ;
        RECT 130.195 218.435 130.525 218.805 ;
        RECT 127.005 217.535 127.400 218.030 ;
        RECT 127.760 217.865 128.135 218.060 ;
        RECT 127.965 217.720 128.135 217.865 ;
        RECT 128.415 217.730 128.655 218.105 ;
        RECT 128.825 217.535 129.160 218.040 ;
        RECT 129.335 217.705 129.595 218.210 ;
        RECT 129.790 218.085 130.455 218.255 ;
        RECT 129.775 217.535 130.105 217.915 ;
        RECT 130.285 217.705 130.455 218.085 ;
        RECT 131.635 217.535 131.925 218.260 ;
        RECT 132.095 218.210 132.265 219.010 ;
        RECT 132.550 218.985 133.215 219.155 ;
        RECT 133.495 219.030 133.800 219.815 ;
        RECT 133.980 219.615 134.665 220.085 ;
        RECT 133.975 219.095 134.670 219.405 ;
        RECT 132.550 218.840 132.720 218.985 ;
        RECT 132.435 218.510 132.720 218.840 ;
        RECT 132.550 218.255 132.720 218.510 ;
        RECT 132.955 218.435 133.285 218.805 ;
        RECT 132.095 217.705 132.355 218.210 ;
        RECT 132.550 218.085 133.215 218.255 ;
        RECT 132.535 217.535 132.865 217.915 ;
        RECT 133.045 217.705 133.215 218.085 ;
        RECT 133.495 218.225 133.670 219.030 ;
        RECT 134.845 218.925 135.130 219.870 ;
        RECT 135.305 219.635 135.635 220.085 ;
        RECT 135.805 219.465 135.975 219.895 ;
        RECT 134.270 218.775 135.130 218.925 ;
        RECT 133.845 218.755 135.130 218.775 ;
        RECT 135.300 219.235 135.975 219.465 ;
        RECT 133.845 218.395 134.830 218.755 ;
        RECT 135.300 218.585 135.535 219.235 ;
        RECT 133.495 217.705 133.735 218.225 ;
        RECT 134.660 218.060 134.830 218.395 ;
        RECT 135.000 218.255 135.535 218.585 ;
        RECT 135.315 218.105 135.535 218.255 ;
        RECT 135.705 218.215 136.005 219.065 ;
        RECT 136.235 219.010 136.505 219.915 ;
        RECT 136.675 219.325 137.005 220.085 ;
        RECT 137.185 219.155 137.355 219.915 ;
        RECT 136.235 218.210 136.405 219.010 ;
        RECT 136.690 218.985 137.355 219.155 ;
        RECT 137.615 219.010 137.885 219.915 ;
        RECT 138.055 219.325 138.385 220.085 ;
        RECT 138.565 219.155 138.735 219.915 ;
        RECT 136.690 218.840 136.860 218.985 ;
        RECT 136.575 218.510 136.860 218.840 ;
        RECT 136.690 218.255 136.860 218.510 ;
        RECT 137.095 218.435 137.425 218.805 ;
        RECT 133.905 217.535 134.300 218.030 ;
        RECT 134.660 217.865 135.035 218.060 ;
        RECT 134.865 217.720 135.035 217.865 ;
        RECT 135.315 217.730 135.555 218.105 ;
        RECT 135.725 217.535 136.060 218.040 ;
        RECT 136.235 217.705 136.495 218.210 ;
        RECT 136.690 218.085 137.355 218.255 ;
        RECT 136.675 217.535 137.005 217.915 ;
        RECT 137.185 217.705 137.355 218.085 ;
        RECT 137.615 218.210 137.785 219.010 ;
        RECT 138.070 218.985 138.735 219.155 ;
        RECT 138.995 218.995 140.205 220.085 ;
        RECT 138.070 218.840 138.240 218.985 ;
        RECT 137.955 218.510 138.240 218.840 ;
        RECT 138.070 218.255 138.240 218.510 ;
        RECT 138.475 218.435 138.805 218.805 ;
        RECT 138.995 218.285 139.515 218.825 ;
        RECT 139.685 218.455 140.205 218.995 ;
        RECT 140.465 219.155 140.635 219.915 ;
        RECT 140.815 219.325 141.145 220.085 ;
        RECT 140.465 218.985 141.130 219.155 ;
        RECT 141.315 219.010 141.585 219.915 ;
        RECT 140.960 218.840 141.130 218.985 ;
        RECT 140.395 218.435 140.725 218.805 ;
        RECT 140.960 218.510 141.245 218.840 ;
        RECT 137.615 217.705 137.875 218.210 ;
        RECT 138.070 218.085 138.735 218.255 ;
        RECT 138.055 217.535 138.385 217.915 ;
        RECT 138.565 217.705 138.735 218.085 ;
        RECT 138.995 217.535 140.205 218.285 ;
        RECT 140.960 218.255 141.130 218.510 ;
        RECT 140.465 218.085 141.130 218.255 ;
        RECT 141.415 218.210 141.585 219.010 ;
        RECT 141.755 218.995 144.345 220.085 ;
        RECT 140.465 217.705 140.635 218.085 ;
        RECT 140.815 217.535 141.145 217.915 ;
        RECT 141.325 217.705 141.585 218.210 ;
        RECT 141.755 218.305 142.965 218.825 ;
        RECT 143.135 218.475 144.345 218.995 ;
        RECT 144.515 218.920 144.805 220.085 ;
        RECT 144.980 218.945 145.330 220.085 ;
        RECT 144.980 218.525 145.330 218.775 ;
        RECT 145.500 218.525 145.945 219.915 ;
        RECT 146.350 218.775 146.590 219.855 ;
        RECT 146.115 218.525 146.590 218.775 ;
        RECT 141.755 217.535 144.345 218.305 ;
        RECT 144.515 217.535 144.805 218.260 ;
        RECT 145.065 217.535 145.235 218.355 ;
        RECT 145.405 218.185 146.590 218.355 ;
        RECT 145.405 217.705 145.735 218.185 ;
        RECT 145.905 217.535 146.075 218.015 ;
        RECT 146.260 217.705 146.590 218.185 ;
        RECT 146.835 218.275 147.050 219.915 ;
        RECT 147.220 218.945 147.565 220.085 ;
        RECT 147.735 219.010 148.005 219.915 ;
        RECT 148.175 219.325 148.505 220.085 ;
        RECT 148.685 219.155 148.855 219.915 ;
        RECT 147.220 218.445 147.565 218.775 ;
        RECT 146.835 217.710 147.565 218.275 ;
        RECT 147.735 218.210 147.905 219.010 ;
        RECT 148.190 218.985 148.855 219.155 ;
        RECT 149.115 219.010 149.385 219.915 ;
        RECT 149.555 219.325 149.885 220.085 ;
        RECT 150.065 219.155 150.235 219.915 ;
        RECT 148.190 218.840 148.360 218.985 ;
        RECT 148.075 218.510 148.360 218.840 ;
        RECT 148.190 218.255 148.360 218.510 ;
        RECT 148.595 218.435 148.925 218.805 ;
        RECT 147.735 217.705 147.995 218.210 ;
        RECT 148.190 218.085 148.855 218.255 ;
        RECT 148.175 217.535 148.505 217.915 ;
        RECT 148.685 217.705 148.855 218.085 ;
        RECT 149.115 218.210 149.285 219.010 ;
        RECT 149.570 218.985 150.235 219.155 ;
        RECT 151.415 219.010 151.685 219.915 ;
        RECT 151.855 219.325 152.185 220.085 ;
        RECT 152.365 219.155 152.535 219.915 ;
        RECT 149.570 218.840 149.740 218.985 ;
        RECT 149.455 218.510 149.740 218.840 ;
        RECT 149.570 218.255 149.740 218.510 ;
        RECT 149.975 218.435 150.305 218.805 ;
        RECT 149.115 217.705 149.375 218.210 ;
        RECT 149.570 218.085 150.235 218.255 ;
        RECT 149.555 217.535 149.885 217.915 ;
        RECT 150.065 217.705 150.235 218.085 ;
        RECT 151.415 218.210 151.585 219.010 ;
        RECT 151.870 218.985 152.535 219.155 ;
        RECT 152.795 218.995 156.305 220.085 ;
        RECT 151.870 218.840 152.040 218.985 ;
        RECT 151.755 218.510 152.040 218.840 ;
        RECT 151.870 218.255 152.040 218.510 ;
        RECT 152.275 218.435 152.605 218.805 ;
        RECT 152.795 218.305 154.445 218.825 ;
        RECT 154.615 218.475 156.305 218.995 ;
        RECT 156.935 218.995 158.145 220.085 ;
        RECT 156.935 218.455 157.455 218.995 ;
        RECT 151.415 217.705 151.675 218.210 ;
        RECT 151.870 218.085 152.535 218.255 ;
        RECT 151.855 217.535 152.185 217.915 ;
        RECT 152.365 217.705 152.535 218.085 ;
        RECT 152.795 217.535 156.305 218.305 ;
        RECT 157.625 218.285 158.145 218.825 ;
        RECT 156.935 217.535 158.145 218.285 ;
        RECT 2.750 217.365 158.230 217.535 ;
        RECT 2.835 216.615 4.045 217.365 ;
        RECT 4.220 216.815 4.475 217.105 ;
        RECT 4.645 216.985 4.975 217.365 ;
        RECT 4.220 216.645 4.970 216.815 ;
        RECT 2.835 216.075 3.355 216.615 ;
        RECT 3.525 215.905 4.045 216.445 ;
        RECT 2.835 214.815 4.045 215.905 ;
        RECT 4.220 215.825 4.570 216.475 ;
        RECT 4.740 215.655 4.970 216.645 ;
        RECT 4.220 215.485 4.970 215.655 ;
        RECT 4.220 214.985 4.475 215.485 ;
        RECT 4.645 214.815 4.975 215.315 ;
        RECT 5.145 214.985 5.315 217.105 ;
        RECT 5.675 217.005 6.005 217.365 ;
        RECT 6.175 216.975 6.670 217.145 ;
        RECT 6.875 216.975 7.730 217.145 ;
        RECT 5.545 215.785 6.005 216.835 ;
        RECT 5.485 215.000 5.810 215.785 ;
        RECT 6.175 215.615 6.345 216.975 ;
        RECT 6.515 216.065 6.865 216.685 ;
        RECT 7.035 216.465 7.390 216.685 ;
        RECT 7.035 215.875 7.205 216.465 ;
        RECT 7.560 216.265 7.730 216.975 ;
        RECT 8.605 216.905 8.935 217.365 ;
        RECT 9.145 217.005 9.495 217.175 ;
        RECT 7.935 216.435 8.725 216.685 ;
        RECT 9.145 216.615 9.405 217.005 ;
        RECT 9.715 216.915 10.665 217.195 ;
        RECT 10.835 216.925 11.025 217.365 ;
        RECT 11.195 216.985 12.265 217.155 ;
        RECT 8.895 216.265 9.065 216.445 ;
        RECT 6.175 215.445 6.570 215.615 ;
        RECT 6.740 215.485 7.205 215.875 ;
        RECT 7.375 216.095 9.065 216.265 ;
        RECT 6.400 215.315 6.570 215.445 ;
        RECT 7.375 215.315 7.545 216.095 ;
        RECT 9.235 215.925 9.405 216.615 ;
        RECT 7.905 215.755 9.405 215.925 ;
        RECT 9.595 215.955 9.805 216.745 ;
        RECT 9.975 216.125 10.325 216.745 ;
        RECT 10.495 216.135 10.665 216.915 ;
        RECT 11.195 216.755 11.365 216.985 ;
        RECT 10.835 216.585 11.365 216.755 ;
        RECT 10.835 216.305 11.055 216.585 ;
        RECT 11.535 216.415 11.775 216.815 ;
        RECT 10.495 215.965 10.900 216.135 ;
        RECT 11.235 216.045 11.775 216.415 ;
        RECT 11.945 216.630 12.265 216.985 ;
        RECT 11.945 216.375 12.270 216.630 ;
        RECT 12.465 216.555 12.635 217.365 ;
        RECT 12.805 216.715 13.135 217.195 ;
        RECT 13.305 216.895 13.475 217.365 ;
        RECT 13.645 216.715 13.975 217.195 ;
        RECT 14.145 216.895 14.315 217.365 ;
        RECT 15.345 216.815 15.515 217.195 ;
        RECT 15.695 216.985 16.025 217.365 ;
        RECT 12.805 216.545 14.570 216.715 ;
        RECT 15.345 216.645 16.010 216.815 ;
        RECT 16.205 216.690 16.465 217.195 ;
        RECT 11.945 216.165 13.975 216.375 ;
        RECT 11.945 216.155 12.290 216.165 ;
        RECT 9.595 215.795 10.270 215.955 ;
        RECT 10.730 215.875 10.900 215.965 ;
        RECT 9.595 215.785 10.560 215.795 ;
        RECT 9.235 215.615 9.405 215.755 ;
        RECT 5.980 214.815 6.230 215.275 ;
        RECT 6.400 214.985 6.650 215.315 ;
        RECT 6.865 214.985 7.545 215.315 ;
        RECT 7.715 215.415 8.790 215.585 ;
        RECT 9.235 215.445 9.795 215.615 ;
        RECT 10.100 215.495 10.560 215.785 ;
        RECT 10.730 215.705 11.950 215.875 ;
        RECT 7.715 215.075 7.885 215.415 ;
        RECT 8.120 214.815 8.450 215.245 ;
        RECT 8.620 215.075 8.790 215.415 ;
        RECT 9.085 214.815 9.455 215.275 ;
        RECT 9.625 214.985 9.795 215.445 ;
        RECT 10.730 215.325 10.900 215.705 ;
        RECT 12.120 215.535 12.290 216.155 ;
        RECT 14.160 215.995 14.570 216.545 ;
        RECT 15.275 216.095 15.605 216.465 ;
        RECT 15.840 216.390 16.010 216.645 ;
        RECT 10.030 214.985 10.900 215.325 ;
        RECT 11.490 215.365 12.290 215.535 ;
        RECT 11.070 214.815 11.320 215.275 ;
        RECT 11.490 215.075 11.660 215.365 ;
        RECT 11.840 214.815 12.170 215.195 ;
        RECT 12.465 214.815 12.635 215.875 ;
        RECT 12.845 215.825 14.570 215.995 ;
        RECT 15.840 216.060 16.125 216.390 ;
        RECT 15.840 215.915 16.010 216.060 ;
        RECT 12.845 214.985 13.135 215.825 ;
        RECT 13.305 214.815 13.475 215.655 ;
        RECT 13.685 214.985 13.935 215.825 ;
        RECT 15.345 215.745 16.010 215.915 ;
        RECT 16.295 215.890 16.465 216.690 ;
        RECT 16.725 216.815 16.895 217.195 ;
        RECT 17.075 216.985 17.405 217.365 ;
        RECT 16.725 216.645 17.390 216.815 ;
        RECT 17.585 216.690 17.845 217.195 ;
        RECT 16.655 216.095 16.985 216.465 ;
        RECT 17.220 216.390 17.390 216.645 ;
        RECT 17.220 216.060 17.505 216.390 ;
        RECT 17.220 215.915 17.390 216.060 ;
        RECT 14.145 214.815 14.315 215.655 ;
        RECT 15.345 214.985 15.515 215.745 ;
        RECT 15.695 214.815 16.025 215.575 ;
        RECT 16.195 214.985 16.465 215.890 ;
        RECT 16.725 215.745 17.390 215.915 ;
        RECT 17.675 215.890 17.845 216.690 ;
        RECT 16.725 214.985 16.895 215.745 ;
        RECT 17.075 214.815 17.405 215.575 ;
        RECT 17.575 214.985 17.845 215.890 ;
        RECT 18.020 216.625 18.275 217.195 ;
        RECT 18.445 216.965 18.775 217.365 ;
        RECT 19.200 216.830 19.730 217.195 ;
        RECT 19.920 217.025 20.195 217.195 ;
        RECT 19.915 216.855 20.195 217.025 ;
        RECT 19.200 216.795 19.375 216.830 ;
        RECT 18.445 216.625 19.375 216.795 ;
        RECT 18.020 215.955 18.190 216.625 ;
        RECT 18.445 216.455 18.615 216.625 ;
        RECT 18.360 216.125 18.615 216.455 ;
        RECT 18.840 216.125 19.035 216.455 ;
        RECT 18.020 214.985 18.355 215.955 ;
        RECT 18.525 214.815 18.695 215.955 ;
        RECT 18.865 215.155 19.035 216.125 ;
        RECT 19.205 215.495 19.375 216.625 ;
        RECT 19.545 215.835 19.715 216.635 ;
        RECT 19.920 216.035 20.195 216.855 ;
        RECT 20.365 215.835 20.555 217.195 ;
        RECT 20.735 216.830 21.245 217.365 ;
        RECT 21.465 216.555 21.710 217.160 ;
        RECT 23.080 216.625 23.335 217.195 ;
        RECT 23.505 216.965 23.835 217.365 ;
        RECT 24.260 216.830 24.790 217.195 ;
        RECT 24.980 217.025 25.255 217.195 ;
        RECT 24.975 216.855 25.255 217.025 ;
        RECT 24.260 216.795 24.435 216.830 ;
        RECT 23.505 216.625 24.435 216.795 ;
        RECT 20.755 216.385 21.985 216.555 ;
        RECT 19.545 215.665 20.555 215.835 ;
        RECT 20.725 215.820 21.475 216.010 ;
        RECT 19.205 215.325 20.330 215.495 ;
        RECT 20.725 215.155 20.895 215.820 ;
        RECT 21.645 215.575 21.985 216.385 ;
        RECT 18.865 214.985 20.895 215.155 ;
        RECT 21.065 214.815 21.235 215.575 ;
        RECT 21.470 215.165 21.985 215.575 ;
        RECT 23.080 215.955 23.250 216.625 ;
        RECT 23.505 216.455 23.675 216.625 ;
        RECT 23.420 216.125 23.675 216.455 ;
        RECT 23.900 216.125 24.095 216.455 ;
        RECT 23.080 214.985 23.415 215.955 ;
        RECT 23.585 214.815 23.755 215.955 ;
        RECT 23.925 215.155 24.095 216.125 ;
        RECT 24.265 215.495 24.435 216.625 ;
        RECT 24.605 215.835 24.775 216.635 ;
        RECT 24.980 216.035 25.255 216.855 ;
        RECT 25.425 215.835 25.615 217.195 ;
        RECT 25.795 216.830 26.305 217.365 ;
        RECT 26.525 216.555 26.770 217.160 ;
        RECT 27.305 216.815 27.475 217.195 ;
        RECT 27.655 216.985 27.985 217.365 ;
        RECT 27.305 216.645 27.970 216.815 ;
        RECT 28.165 216.690 28.425 217.195 ;
        RECT 25.815 216.385 27.045 216.555 ;
        RECT 24.605 215.665 25.615 215.835 ;
        RECT 25.785 215.820 26.535 216.010 ;
        RECT 24.265 215.325 25.390 215.495 ;
        RECT 25.785 215.155 25.955 215.820 ;
        RECT 26.705 215.575 27.045 216.385 ;
        RECT 27.235 216.095 27.565 216.465 ;
        RECT 27.800 216.390 27.970 216.645 ;
        RECT 27.800 216.060 28.085 216.390 ;
        RECT 27.800 215.915 27.970 216.060 ;
        RECT 23.925 214.985 25.955 215.155 ;
        RECT 26.125 214.815 26.295 215.575 ;
        RECT 26.530 215.165 27.045 215.575 ;
        RECT 27.305 215.745 27.970 215.915 ;
        RECT 28.255 215.890 28.425 216.690 ;
        RECT 28.595 216.640 28.885 217.365 ;
        RECT 29.145 216.815 29.315 217.195 ;
        RECT 29.495 216.985 29.825 217.365 ;
        RECT 29.145 216.645 29.810 216.815 ;
        RECT 30.005 216.690 30.265 217.195 ;
        RECT 29.075 216.095 29.405 216.465 ;
        RECT 29.640 216.390 29.810 216.645 ;
        RECT 29.640 216.060 29.925 216.390 ;
        RECT 27.305 214.985 27.475 215.745 ;
        RECT 27.655 214.815 27.985 215.575 ;
        RECT 28.155 214.985 28.425 215.890 ;
        RECT 28.595 214.815 28.885 215.980 ;
        RECT 29.640 215.915 29.810 216.060 ;
        RECT 29.145 215.745 29.810 215.915 ;
        RECT 30.095 215.890 30.265 216.690 ;
        RECT 30.710 216.555 30.955 217.160 ;
        RECT 31.175 216.830 31.685 217.365 ;
        RECT 29.145 214.985 29.315 215.745 ;
        RECT 29.495 214.815 29.825 215.575 ;
        RECT 29.995 214.985 30.265 215.890 ;
        RECT 30.435 216.385 31.665 216.555 ;
        RECT 30.435 215.575 30.775 216.385 ;
        RECT 30.945 215.820 31.695 216.010 ;
        RECT 30.435 215.165 30.950 215.575 ;
        RECT 31.185 214.815 31.355 215.575 ;
        RECT 31.525 215.155 31.695 215.820 ;
        RECT 31.865 215.835 32.055 217.195 ;
        RECT 32.225 217.025 32.500 217.195 ;
        RECT 32.225 216.855 32.505 217.025 ;
        RECT 32.225 216.035 32.500 216.855 ;
        RECT 32.690 216.830 33.220 217.195 ;
        RECT 33.645 216.965 33.975 217.365 ;
        RECT 33.045 216.795 33.220 216.830 ;
        RECT 32.705 215.835 32.875 216.635 ;
        RECT 31.865 215.665 32.875 215.835 ;
        RECT 33.045 216.625 33.975 216.795 ;
        RECT 34.145 216.625 34.400 217.195 ;
        RECT 35.345 216.895 35.515 217.365 ;
        RECT 35.685 216.715 36.015 217.195 ;
        RECT 36.185 216.895 36.355 217.365 ;
        RECT 36.525 216.715 36.855 217.195 ;
        RECT 33.045 215.495 33.215 216.625 ;
        RECT 33.805 216.455 33.975 216.625 ;
        RECT 32.090 215.325 33.215 215.495 ;
        RECT 33.385 216.125 33.580 216.455 ;
        RECT 33.805 216.125 34.060 216.455 ;
        RECT 33.385 215.155 33.555 216.125 ;
        RECT 34.230 215.955 34.400 216.625 ;
        RECT 31.525 214.985 33.555 215.155 ;
        RECT 33.725 214.815 33.895 215.955 ;
        RECT 34.065 214.985 34.400 215.955 ;
        RECT 35.090 216.545 36.855 216.715 ;
        RECT 37.025 216.555 37.195 217.365 ;
        RECT 37.395 216.985 38.465 217.155 ;
        RECT 37.395 216.630 37.715 216.985 ;
        RECT 35.090 215.995 35.500 216.545 ;
        RECT 37.390 216.375 37.715 216.630 ;
        RECT 35.685 216.165 37.715 216.375 ;
        RECT 37.370 216.155 37.715 216.165 ;
        RECT 37.885 216.415 38.125 216.815 ;
        RECT 38.295 216.755 38.465 216.985 ;
        RECT 38.635 216.925 38.825 217.365 ;
        RECT 38.995 216.915 39.945 217.195 ;
        RECT 40.165 217.005 40.515 217.175 ;
        RECT 38.295 216.585 38.825 216.755 ;
        RECT 35.090 215.825 36.815 215.995 ;
        RECT 35.345 214.815 35.515 215.655 ;
        RECT 35.725 214.985 35.975 215.825 ;
        RECT 36.185 214.815 36.355 215.655 ;
        RECT 36.525 214.985 36.815 215.825 ;
        RECT 37.025 214.815 37.195 215.875 ;
        RECT 37.370 215.535 37.540 216.155 ;
        RECT 37.885 216.045 38.425 216.415 ;
        RECT 38.605 216.305 38.825 216.585 ;
        RECT 38.995 216.135 39.165 216.915 ;
        RECT 38.760 215.965 39.165 216.135 ;
        RECT 39.335 216.125 39.685 216.745 ;
        RECT 38.760 215.875 38.930 215.965 ;
        RECT 39.855 215.955 40.065 216.745 ;
        RECT 37.710 215.705 38.930 215.875 ;
        RECT 39.390 215.795 40.065 215.955 ;
        RECT 37.370 215.365 38.170 215.535 ;
        RECT 37.490 214.815 37.820 215.195 ;
        RECT 38.000 215.075 38.170 215.365 ;
        RECT 38.760 215.325 38.930 215.705 ;
        RECT 39.100 215.785 40.065 215.795 ;
        RECT 40.255 216.615 40.515 217.005 ;
        RECT 40.725 216.905 41.055 217.365 ;
        RECT 41.930 216.975 42.785 217.145 ;
        RECT 42.990 216.975 43.485 217.145 ;
        RECT 43.655 217.005 43.985 217.365 ;
        RECT 40.255 215.925 40.425 216.615 ;
        RECT 40.595 216.265 40.765 216.445 ;
        RECT 40.935 216.435 41.725 216.685 ;
        RECT 41.930 216.265 42.100 216.975 ;
        RECT 42.270 216.465 42.625 216.685 ;
        RECT 40.595 216.095 42.285 216.265 ;
        RECT 39.100 215.495 39.560 215.785 ;
        RECT 40.255 215.755 41.755 215.925 ;
        RECT 40.255 215.615 40.425 215.755 ;
        RECT 39.865 215.445 40.425 215.615 ;
        RECT 38.340 214.815 38.590 215.275 ;
        RECT 38.760 214.985 39.630 215.325 ;
        RECT 39.865 214.985 40.035 215.445 ;
        RECT 40.870 215.415 41.945 215.585 ;
        RECT 40.205 214.815 40.575 215.275 ;
        RECT 40.870 215.075 41.040 215.415 ;
        RECT 41.210 214.815 41.540 215.245 ;
        RECT 41.775 215.075 41.945 215.415 ;
        RECT 42.115 215.315 42.285 216.095 ;
        RECT 42.455 215.875 42.625 216.465 ;
        RECT 42.795 216.065 43.145 216.685 ;
        RECT 42.455 215.485 42.920 215.875 ;
        RECT 43.315 215.615 43.485 216.975 ;
        RECT 43.655 215.785 44.115 216.835 ;
        RECT 43.090 215.445 43.485 215.615 ;
        RECT 43.090 215.315 43.260 215.445 ;
        RECT 42.115 214.985 42.795 215.315 ;
        RECT 43.010 214.985 43.260 215.315 ;
        RECT 43.430 214.815 43.680 215.275 ;
        RECT 43.850 215.000 44.175 215.785 ;
        RECT 44.345 214.985 44.515 217.105 ;
        RECT 44.685 216.985 45.015 217.365 ;
        RECT 45.185 216.815 45.440 217.105 ;
        RECT 44.690 216.645 45.440 216.815 ;
        RECT 44.690 215.655 44.920 216.645 ;
        RECT 46.080 216.625 46.335 217.195 ;
        RECT 46.505 216.965 46.835 217.365 ;
        RECT 47.260 216.830 47.790 217.195 ;
        RECT 47.260 216.795 47.435 216.830 ;
        RECT 46.505 216.625 47.435 216.795 ;
        RECT 47.980 216.685 48.255 217.195 ;
        RECT 45.090 215.825 45.440 216.475 ;
        RECT 46.080 215.955 46.250 216.625 ;
        RECT 46.505 216.455 46.675 216.625 ;
        RECT 46.420 216.125 46.675 216.455 ;
        RECT 46.900 216.125 47.095 216.455 ;
        RECT 44.690 215.485 45.440 215.655 ;
        RECT 44.685 214.815 45.015 215.315 ;
        RECT 45.185 214.985 45.440 215.485 ;
        RECT 46.080 214.985 46.415 215.955 ;
        RECT 46.585 214.815 46.755 215.955 ;
        RECT 46.925 215.155 47.095 216.125 ;
        RECT 47.265 215.495 47.435 216.625 ;
        RECT 47.605 215.835 47.775 216.635 ;
        RECT 47.975 216.515 48.255 216.685 ;
        RECT 47.980 216.035 48.255 216.515 ;
        RECT 48.425 215.835 48.615 217.195 ;
        RECT 48.795 216.830 49.305 217.365 ;
        RECT 49.525 216.555 49.770 217.160 ;
        RECT 50.220 216.625 50.475 217.195 ;
        RECT 50.645 216.965 50.975 217.365 ;
        RECT 51.400 216.830 51.930 217.195 ;
        RECT 51.400 216.795 51.575 216.830 ;
        RECT 50.645 216.625 51.575 216.795 ;
        RECT 48.815 216.385 50.045 216.555 ;
        RECT 47.605 215.665 48.615 215.835 ;
        RECT 48.785 215.820 49.535 216.010 ;
        RECT 47.265 215.325 48.390 215.495 ;
        RECT 48.785 215.155 48.955 215.820 ;
        RECT 49.705 215.575 50.045 216.385 ;
        RECT 46.925 214.985 48.955 215.155 ;
        RECT 49.125 214.815 49.295 215.575 ;
        RECT 49.530 215.165 50.045 215.575 ;
        RECT 50.220 215.955 50.390 216.625 ;
        RECT 50.645 216.455 50.815 216.625 ;
        RECT 50.560 216.125 50.815 216.455 ;
        RECT 51.040 216.125 51.235 216.455 ;
        RECT 50.220 214.985 50.555 215.955 ;
        RECT 50.725 214.815 50.895 215.955 ;
        RECT 51.065 215.155 51.235 216.125 ;
        RECT 51.405 215.495 51.575 216.625 ;
        RECT 51.745 215.835 51.915 216.635 ;
        RECT 52.120 216.345 52.395 217.195 ;
        RECT 52.115 216.175 52.395 216.345 ;
        RECT 52.120 216.035 52.395 216.175 ;
        RECT 52.565 215.835 52.755 217.195 ;
        RECT 52.935 216.830 53.445 217.365 ;
        RECT 53.665 216.555 53.910 217.160 ;
        RECT 54.355 216.640 54.645 217.365 ;
        RECT 54.820 216.625 55.075 217.195 ;
        RECT 55.245 216.965 55.575 217.365 ;
        RECT 56.000 216.830 56.530 217.195 ;
        RECT 56.000 216.795 56.175 216.830 ;
        RECT 55.245 216.625 56.175 216.795 ;
        RECT 52.955 216.385 54.185 216.555 ;
        RECT 51.745 215.665 52.755 215.835 ;
        RECT 52.925 215.820 53.675 216.010 ;
        RECT 51.405 215.325 52.530 215.495 ;
        RECT 52.925 215.155 53.095 215.820 ;
        RECT 53.845 215.575 54.185 216.385 ;
        RECT 51.065 214.985 53.095 215.155 ;
        RECT 53.265 214.815 53.435 215.575 ;
        RECT 53.670 215.165 54.185 215.575 ;
        RECT 54.355 214.815 54.645 215.980 ;
        RECT 54.820 215.955 54.990 216.625 ;
        RECT 55.245 216.455 55.415 216.625 ;
        RECT 55.160 216.125 55.415 216.455 ;
        RECT 55.640 216.125 55.835 216.455 ;
        RECT 54.820 214.985 55.155 215.955 ;
        RECT 55.325 214.815 55.495 215.955 ;
        RECT 55.665 215.155 55.835 216.125 ;
        RECT 56.005 215.495 56.175 216.625 ;
        RECT 56.345 215.835 56.515 216.635 ;
        RECT 56.720 216.345 56.995 217.195 ;
        RECT 56.715 216.175 56.995 216.345 ;
        RECT 56.720 216.035 56.995 216.175 ;
        RECT 57.165 215.835 57.355 217.195 ;
        RECT 57.535 216.830 58.045 217.365 ;
        RECT 58.265 216.555 58.510 217.160 ;
        RECT 58.955 216.615 60.165 217.365 ;
        RECT 60.340 216.625 60.595 217.195 ;
        RECT 60.765 216.965 61.095 217.365 ;
        RECT 61.520 216.830 62.050 217.195 ;
        RECT 61.520 216.795 61.695 216.830 ;
        RECT 60.765 216.625 61.695 216.795 ;
        RECT 57.555 216.385 58.785 216.555 ;
        RECT 56.345 215.665 57.355 215.835 ;
        RECT 57.525 215.820 58.275 216.010 ;
        RECT 56.005 215.325 57.130 215.495 ;
        RECT 57.525 215.155 57.695 215.820 ;
        RECT 58.445 215.575 58.785 216.385 ;
        RECT 58.955 216.075 59.475 216.615 ;
        RECT 59.645 215.905 60.165 216.445 ;
        RECT 55.665 214.985 57.695 215.155 ;
        RECT 57.865 214.815 58.035 215.575 ;
        RECT 58.270 215.165 58.785 215.575 ;
        RECT 58.955 214.815 60.165 215.905 ;
        RECT 60.340 215.955 60.510 216.625 ;
        RECT 60.765 216.455 60.935 216.625 ;
        RECT 60.680 216.125 60.935 216.455 ;
        RECT 61.160 216.125 61.355 216.455 ;
        RECT 60.340 214.985 60.675 215.955 ;
        RECT 60.845 214.815 61.015 215.955 ;
        RECT 61.185 215.155 61.355 216.125 ;
        RECT 61.525 215.495 61.695 216.625 ;
        RECT 61.865 215.835 62.035 216.635 ;
        RECT 62.240 216.345 62.515 217.195 ;
        RECT 62.235 216.175 62.515 216.345 ;
        RECT 62.240 216.035 62.515 216.175 ;
        RECT 62.685 215.835 62.875 217.195 ;
        RECT 63.055 216.830 63.565 217.365 ;
        RECT 63.785 216.555 64.030 217.160 ;
        RECT 64.535 216.885 64.815 217.365 ;
        RECT 64.985 216.715 65.245 217.105 ;
        RECT 65.420 216.885 65.675 217.365 ;
        RECT 65.845 216.715 66.140 217.105 ;
        RECT 66.320 216.885 66.595 217.365 ;
        RECT 66.765 216.865 67.065 217.195 ;
        RECT 67.695 216.985 68.585 217.155 ;
        RECT 63.075 216.385 64.305 216.555 ;
        RECT 61.865 215.665 62.875 215.835 ;
        RECT 63.045 215.820 63.795 216.010 ;
        RECT 61.525 215.325 62.650 215.495 ;
        RECT 63.045 215.155 63.215 215.820 ;
        RECT 63.965 215.575 64.305 216.385 ;
        RECT 64.490 216.545 66.140 216.715 ;
        RECT 64.490 216.035 64.895 216.545 ;
        RECT 65.065 216.205 66.205 216.375 ;
        RECT 64.490 215.865 65.245 216.035 ;
        RECT 61.185 214.985 63.215 215.155 ;
        RECT 63.385 214.815 63.555 215.575 ;
        RECT 63.790 215.165 64.305 215.575 ;
        RECT 64.530 214.815 64.815 215.685 ;
        RECT 64.985 215.615 65.245 215.865 ;
        RECT 66.035 215.955 66.205 216.205 ;
        RECT 66.375 216.125 66.725 216.695 ;
        RECT 66.895 215.955 67.065 216.865 ;
        RECT 67.695 216.430 68.245 216.815 ;
        RECT 68.415 216.260 68.585 216.985 ;
        RECT 66.035 215.785 67.065 215.955 ;
        RECT 64.985 215.445 66.105 215.615 ;
        RECT 64.985 214.985 65.245 215.445 ;
        RECT 65.420 214.815 65.675 215.275 ;
        RECT 65.845 214.985 66.105 215.445 ;
        RECT 66.275 214.815 66.585 215.615 ;
        RECT 66.755 214.985 67.065 215.785 ;
        RECT 67.695 216.190 68.585 216.260 ;
        RECT 68.755 216.660 68.975 217.145 ;
        RECT 69.145 216.825 69.395 217.365 ;
        RECT 69.565 216.715 69.825 217.195 ;
        RECT 68.755 216.235 69.085 216.660 ;
        RECT 67.695 216.165 68.590 216.190 ;
        RECT 67.695 216.150 68.600 216.165 ;
        RECT 67.695 216.135 68.605 216.150 ;
        RECT 67.695 216.130 68.615 216.135 ;
        RECT 67.695 216.120 68.620 216.130 ;
        RECT 67.695 216.110 68.625 216.120 ;
        RECT 67.695 216.105 68.635 216.110 ;
        RECT 67.695 216.095 68.645 216.105 ;
        RECT 67.695 216.090 68.655 216.095 ;
        RECT 67.695 215.640 67.955 216.090 ;
        RECT 68.320 216.085 68.655 216.090 ;
        RECT 68.320 216.080 68.670 216.085 ;
        RECT 68.320 216.070 68.685 216.080 ;
        RECT 68.320 216.065 68.710 216.070 ;
        RECT 69.255 216.065 69.485 216.460 ;
        RECT 68.320 216.060 69.485 216.065 ;
        RECT 68.350 216.025 69.485 216.060 ;
        RECT 68.385 216.000 69.485 216.025 ;
        RECT 68.415 215.970 69.485 216.000 ;
        RECT 68.435 215.940 69.485 215.970 ;
        RECT 68.455 215.910 69.485 215.940 ;
        RECT 68.525 215.900 69.485 215.910 ;
        RECT 68.550 215.890 69.485 215.900 ;
        RECT 68.570 215.875 69.485 215.890 ;
        RECT 68.590 215.860 69.485 215.875 ;
        RECT 68.595 215.850 69.380 215.860 ;
        RECT 68.610 215.815 69.380 215.850 ;
        RECT 68.125 215.495 68.455 215.740 ;
        RECT 68.625 215.565 69.380 215.815 ;
        RECT 69.655 215.685 69.825 216.715 ;
        RECT 68.125 215.470 68.310 215.495 ;
        RECT 67.695 215.370 68.310 215.470 ;
        RECT 67.695 214.815 68.300 215.370 ;
        RECT 68.475 214.985 68.955 215.325 ;
        RECT 69.125 214.815 69.380 215.360 ;
        RECT 69.550 214.985 69.825 215.685 ;
        RECT 70.455 216.865 70.755 217.195 ;
        RECT 70.925 216.885 71.200 217.365 ;
        RECT 70.455 215.955 70.625 216.865 ;
        RECT 71.380 216.715 71.675 217.105 ;
        RECT 71.845 216.885 72.100 217.365 ;
        RECT 72.275 216.715 72.535 217.105 ;
        RECT 72.705 216.885 72.985 217.365 ;
        RECT 70.795 216.125 71.145 216.695 ;
        RECT 71.380 216.545 73.030 216.715 ;
        RECT 71.315 216.205 72.455 216.375 ;
        RECT 71.315 215.955 71.485 216.205 ;
        RECT 72.625 216.035 73.030 216.545 ;
        RECT 73.215 216.595 74.885 217.365 ;
        RECT 75.605 216.715 75.775 217.195 ;
        RECT 75.945 216.885 76.275 217.365 ;
        RECT 76.500 216.945 78.035 217.195 ;
        RECT 76.500 216.715 76.670 216.945 ;
        RECT 73.215 216.075 73.965 216.595 ;
        RECT 75.605 216.545 76.670 216.715 ;
        RECT 70.455 215.785 71.485 215.955 ;
        RECT 72.275 215.865 73.030 216.035 ;
        RECT 74.135 215.905 74.885 216.425 ;
        RECT 76.850 216.375 77.130 216.775 ;
        RECT 75.520 216.165 75.870 216.375 ;
        RECT 76.040 216.175 76.485 216.375 ;
        RECT 76.655 216.175 77.130 216.375 ;
        RECT 77.400 216.375 77.685 216.775 ;
        RECT 77.865 216.715 78.035 216.945 ;
        RECT 78.205 216.885 78.535 217.365 ;
        RECT 78.750 216.865 79.005 217.195 ;
        RECT 78.795 216.855 79.005 216.865 ;
        RECT 78.820 216.785 79.005 216.855 ;
        RECT 77.865 216.545 78.665 216.715 ;
        RECT 77.400 216.175 77.730 216.375 ;
        RECT 77.900 216.345 78.265 216.375 ;
        RECT 77.900 216.175 78.275 216.345 ;
        RECT 78.495 215.995 78.665 216.545 ;
        RECT 70.455 214.985 70.765 215.785 ;
        RECT 72.275 215.615 72.535 215.865 ;
        RECT 70.935 214.815 71.245 215.615 ;
        RECT 71.415 215.445 72.535 215.615 ;
        RECT 71.415 214.985 71.675 215.445 ;
        RECT 71.845 214.815 72.100 215.275 ;
        RECT 72.275 214.985 72.535 215.445 ;
        RECT 72.705 214.815 72.990 215.685 ;
        RECT 73.215 214.815 74.885 215.905 ;
        RECT 75.605 215.825 78.665 215.995 ;
        RECT 75.605 214.985 75.775 215.825 ;
        RECT 78.835 215.655 79.005 216.785 ;
        RECT 80.115 216.640 80.405 217.365 ;
        RECT 80.575 216.645 80.915 217.155 ;
        RECT 75.945 215.155 76.275 215.655 ;
        RECT 76.445 215.415 78.080 215.655 ;
        RECT 76.445 215.325 76.675 215.415 ;
        RECT 76.785 215.155 77.115 215.195 ;
        RECT 75.945 214.985 77.115 215.155 ;
        RECT 77.305 214.815 77.660 215.235 ;
        RECT 77.830 214.985 78.080 215.415 ;
        RECT 78.250 214.815 78.580 215.575 ;
        RECT 78.750 214.985 79.005 215.655 ;
        RECT 80.115 214.815 80.405 215.980 ;
        RECT 80.575 215.245 80.835 216.645 ;
        RECT 81.085 216.565 81.355 217.365 ;
        RECT 81.010 216.125 81.340 216.375 ;
        RECT 81.535 216.125 81.815 217.095 ;
        RECT 81.995 216.125 82.295 217.095 ;
        RECT 82.475 216.125 82.825 217.090 ;
        RECT 83.045 216.865 83.540 217.195 ;
        RECT 81.025 215.955 81.340 216.125 ;
        RECT 83.045 215.955 83.215 216.865 ;
        RECT 83.795 216.820 89.140 217.365 ;
        RECT 81.025 215.785 83.215 215.955 ;
        RECT 80.575 214.985 80.915 215.245 ;
        RECT 81.085 214.815 81.415 215.615 ;
        RECT 81.880 214.985 82.130 215.785 ;
        RECT 82.315 214.815 82.645 215.535 ;
        RECT 82.865 214.985 83.115 215.785 ;
        RECT 83.385 215.375 83.625 216.685 ;
        RECT 85.380 215.990 85.720 216.820 ;
        RECT 89.315 216.595 91.905 217.365 ;
        RECT 87.200 215.250 87.550 216.500 ;
        RECT 89.315 216.075 90.525 216.595 ;
        RECT 90.695 215.905 91.905 216.425 ;
        RECT 83.285 214.815 83.620 215.195 ;
        RECT 83.795 214.815 89.140 215.250 ;
        RECT 89.315 214.815 91.905 215.905 ;
        RECT 92.535 216.420 92.875 217.195 ;
        RECT 93.045 216.905 93.215 217.365 ;
        RECT 93.455 216.930 93.815 217.195 ;
        RECT 93.455 216.925 93.810 216.930 ;
        RECT 93.455 216.915 93.805 216.925 ;
        RECT 93.455 216.910 93.800 216.915 ;
        RECT 93.455 216.900 93.795 216.910 ;
        RECT 94.445 216.905 94.615 217.365 ;
        RECT 93.455 216.895 93.790 216.900 ;
        RECT 93.455 216.885 93.780 216.895 ;
        RECT 93.455 216.875 93.770 216.885 ;
        RECT 93.455 216.735 93.755 216.875 ;
        RECT 93.045 216.545 93.755 216.735 ;
        RECT 93.945 216.735 94.275 216.815 ;
        RECT 94.785 216.735 95.125 217.195 ;
        RECT 93.945 216.545 95.125 216.735 ;
        RECT 95.295 216.715 95.555 217.195 ;
        RECT 95.725 216.825 95.975 217.365 ;
        RECT 92.535 214.985 92.815 216.420 ;
        RECT 93.045 215.975 93.330 216.545 ;
        RECT 93.515 216.145 93.985 216.375 ;
        RECT 94.155 216.355 94.485 216.375 ;
        RECT 94.155 216.175 94.605 216.355 ;
        RECT 94.795 216.175 95.125 216.375 ;
        RECT 93.045 215.760 94.195 215.975 ;
        RECT 92.985 214.815 93.695 215.590 ;
        RECT 93.865 214.985 94.195 215.760 ;
        RECT 94.390 215.060 94.605 216.175 ;
        RECT 94.895 215.835 95.125 216.175 ;
        RECT 95.295 215.685 95.465 216.715 ;
        RECT 96.145 216.660 96.365 217.145 ;
        RECT 95.635 216.065 95.865 216.460 ;
        RECT 96.035 216.235 96.365 216.660 ;
        RECT 96.535 216.985 97.425 217.155 ;
        RECT 96.535 216.260 96.705 216.985 ;
        RECT 96.875 216.430 97.425 216.815 ;
        RECT 97.595 216.595 100.185 217.365 ;
        RECT 96.535 216.190 97.425 216.260 ;
        RECT 96.530 216.165 97.425 216.190 ;
        RECT 96.520 216.150 97.425 216.165 ;
        RECT 96.515 216.135 97.425 216.150 ;
        RECT 96.505 216.130 97.425 216.135 ;
        RECT 96.500 216.120 97.425 216.130 ;
        RECT 96.495 216.110 97.425 216.120 ;
        RECT 96.485 216.105 97.425 216.110 ;
        RECT 96.475 216.095 97.425 216.105 ;
        RECT 96.465 216.090 97.425 216.095 ;
        RECT 96.465 216.085 96.800 216.090 ;
        RECT 96.450 216.080 96.800 216.085 ;
        RECT 96.435 216.070 96.800 216.080 ;
        RECT 96.410 216.065 96.800 216.070 ;
        RECT 95.635 216.060 96.800 216.065 ;
        RECT 95.635 216.025 96.770 216.060 ;
        RECT 95.635 216.000 96.735 216.025 ;
        RECT 95.635 215.970 96.705 216.000 ;
        RECT 95.635 215.940 96.685 215.970 ;
        RECT 95.635 215.910 96.665 215.940 ;
        RECT 95.635 215.900 96.595 215.910 ;
        RECT 95.635 215.890 96.570 215.900 ;
        RECT 95.635 215.875 96.550 215.890 ;
        RECT 95.635 215.860 96.530 215.875 ;
        RECT 95.740 215.850 96.525 215.860 ;
        RECT 95.740 215.815 96.510 215.850 ;
        RECT 94.785 214.815 95.115 215.535 ;
        RECT 95.295 214.985 95.570 215.685 ;
        RECT 95.740 215.565 96.495 215.815 ;
        RECT 96.665 215.495 96.995 215.740 ;
        RECT 97.165 215.640 97.425 216.090 ;
        RECT 97.595 216.075 98.805 216.595 ;
        RECT 100.825 216.555 101.095 217.365 ;
        RECT 101.265 216.555 101.595 217.195 ;
        RECT 101.765 216.555 102.005 217.365 ;
        RECT 102.195 216.595 105.705 217.365 ;
        RECT 105.875 216.640 106.165 217.365 ;
        RECT 106.335 216.645 106.675 217.155 ;
        RECT 98.975 215.905 100.185 216.425 ;
        RECT 100.815 216.125 101.165 216.375 ;
        RECT 101.335 215.955 101.505 216.555 ;
        RECT 101.675 216.125 102.025 216.375 ;
        RECT 102.195 216.075 103.845 216.595 ;
        RECT 96.810 215.470 96.995 215.495 ;
        RECT 96.810 215.370 97.425 215.470 ;
        RECT 95.740 214.815 95.995 215.360 ;
        RECT 96.165 214.985 96.645 215.325 ;
        RECT 96.820 214.815 97.425 215.370 ;
        RECT 97.595 214.815 100.185 215.905 ;
        RECT 100.825 214.815 101.155 215.955 ;
        RECT 101.335 215.785 102.015 215.955 ;
        RECT 104.015 215.905 105.705 216.425 ;
        RECT 101.685 215.000 102.015 215.785 ;
        RECT 102.195 214.815 105.705 215.905 ;
        RECT 105.875 214.815 106.165 215.980 ;
        RECT 106.335 215.245 106.595 216.645 ;
        RECT 106.845 216.565 107.115 217.365 ;
        RECT 106.770 216.125 107.100 216.375 ;
        RECT 107.295 216.125 107.575 217.095 ;
        RECT 107.755 216.125 108.055 217.095 ;
        RECT 108.235 216.125 108.585 217.090 ;
        RECT 108.805 216.865 109.300 217.195 ;
        RECT 106.785 215.955 107.100 216.125 ;
        RECT 108.805 215.955 108.975 216.865 ;
        RECT 106.785 215.785 108.975 215.955 ;
        RECT 106.335 214.985 106.675 215.245 ;
        RECT 106.845 214.815 107.175 215.615 ;
        RECT 107.640 214.985 107.890 215.785 ;
        RECT 108.075 214.815 108.405 215.535 ;
        RECT 108.625 214.985 108.875 215.785 ;
        RECT 109.145 215.375 109.385 216.685 ;
        RECT 109.555 216.595 112.145 217.365 ;
        RECT 109.555 216.075 110.765 216.595 ;
        RECT 112.980 216.585 113.480 217.195 ;
        RECT 110.935 215.905 112.145 216.425 ;
        RECT 112.775 216.125 113.125 216.375 ;
        RECT 113.310 215.955 113.480 216.585 ;
        RECT 114.110 216.715 114.440 217.195 ;
        RECT 114.610 216.905 114.835 217.365 ;
        RECT 115.005 216.715 115.335 217.195 ;
        RECT 114.110 216.545 115.335 216.715 ;
        RECT 115.525 216.565 115.775 217.365 ;
        RECT 115.945 216.565 116.285 217.195 ;
        RECT 116.465 216.865 116.795 217.365 ;
        RECT 116.995 216.795 117.165 217.145 ;
        RECT 117.365 216.965 117.695 217.365 ;
        RECT 117.865 216.795 118.035 217.145 ;
        RECT 118.205 216.965 118.585 217.365 ;
        RECT 113.650 216.175 113.980 216.375 ;
        RECT 114.150 216.175 114.480 216.375 ;
        RECT 114.650 216.175 115.070 216.375 ;
        RECT 115.245 216.205 115.940 216.375 ;
        RECT 115.245 215.955 115.415 216.205 ;
        RECT 116.110 215.955 116.285 216.565 ;
        RECT 116.460 216.125 116.810 216.695 ;
        RECT 116.995 216.625 118.605 216.795 ;
        RECT 118.775 216.690 119.045 217.035 ;
        RECT 118.435 216.455 118.605 216.625 ;
        RECT 109.045 214.815 109.380 215.195 ;
        RECT 109.555 214.815 112.145 215.905 ;
        RECT 112.980 215.785 115.415 215.955 ;
        RECT 112.980 214.985 113.310 215.785 ;
        RECT 113.480 214.815 113.810 215.615 ;
        RECT 114.110 214.985 114.440 215.785 ;
        RECT 115.085 214.815 115.335 215.615 ;
        RECT 115.605 214.815 115.775 215.955 ;
        RECT 115.945 214.985 116.285 215.955 ;
        RECT 116.460 215.665 116.780 215.955 ;
        RECT 116.980 215.835 117.690 216.455 ;
        RECT 117.860 216.125 118.265 216.455 ;
        RECT 118.435 216.125 118.705 216.455 ;
        RECT 118.435 215.955 118.605 216.125 ;
        RECT 118.875 215.955 119.045 216.690 ;
        RECT 119.215 216.595 120.885 217.365 ;
        RECT 121.525 216.640 121.855 217.150 ;
        RECT 122.025 216.965 122.355 217.365 ;
        RECT 123.405 216.795 123.735 217.135 ;
        RECT 123.905 216.965 124.235 217.365 ;
        RECT 119.215 216.075 119.965 216.595 ;
        RECT 117.880 215.785 118.605 215.955 ;
        RECT 117.880 215.665 118.050 215.785 ;
        RECT 116.460 215.495 118.050 215.665 ;
        RECT 116.460 215.035 118.115 215.325 ;
        RECT 118.285 214.815 118.565 215.615 ;
        RECT 118.775 214.985 119.045 215.955 ;
        RECT 120.135 215.905 120.885 216.425 ;
        RECT 119.215 214.815 120.885 215.905 ;
        RECT 121.525 215.875 121.715 216.640 ;
        RECT 122.025 216.625 124.390 216.795 ;
        RECT 122.025 216.455 122.195 216.625 ;
        RECT 121.885 216.125 122.195 216.455 ;
        RECT 122.365 216.125 122.670 216.455 ;
        RECT 121.525 215.025 121.855 215.875 ;
        RECT 122.025 214.815 122.275 215.955 ;
        RECT 122.455 215.795 122.670 216.125 ;
        RECT 122.845 215.795 123.130 216.455 ;
        RECT 123.325 215.795 123.590 216.455 ;
        RECT 123.805 215.795 124.050 216.455 ;
        RECT 124.220 215.625 124.390 216.625 ;
        RECT 122.465 215.455 123.755 215.625 ;
        RECT 122.465 215.035 122.715 215.455 ;
        RECT 122.945 214.815 123.275 215.285 ;
        RECT 123.505 215.035 123.755 215.455 ;
        RECT 123.935 215.455 124.390 215.625 ;
        RECT 123.935 215.025 124.265 215.455 ;
        RECT 124.745 214.995 125.005 217.185 ;
        RECT 125.265 216.995 125.935 217.365 ;
        RECT 126.115 216.815 126.425 217.185 ;
        RECT 125.195 216.615 126.425 216.815 ;
        RECT 125.195 215.945 125.485 216.615 ;
        RECT 126.605 216.435 126.835 217.075 ;
        RECT 127.015 216.635 127.305 217.365 ;
        RECT 127.520 216.975 127.850 217.365 ;
        RECT 128.020 216.805 128.245 217.185 ;
        RECT 125.665 216.125 126.130 216.435 ;
        RECT 126.310 216.125 126.835 216.435 ;
        RECT 127.015 216.125 127.315 216.455 ;
        RECT 127.505 216.125 127.745 216.775 ;
        RECT 127.915 216.625 128.245 216.805 ;
        RECT 127.915 215.955 128.090 216.625 ;
        RECT 128.445 216.455 128.675 217.075 ;
        RECT 128.855 216.635 129.155 217.365 ;
        RECT 129.335 216.595 131.005 217.365 ;
        RECT 131.635 216.640 131.925 217.365 ;
        RECT 128.260 216.125 128.675 216.455 ;
        RECT 128.855 216.125 129.150 216.455 ;
        RECT 129.335 216.075 130.085 216.595 ;
        RECT 132.555 216.565 132.865 217.365 ;
        RECT 133.070 216.565 133.765 217.195 ;
        RECT 133.935 216.595 136.525 217.365 ;
        RECT 136.715 216.865 136.970 217.195 ;
        RECT 137.185 216.885 137.515 217.365 ;
        RECT 137.685 216.945 139.220 217.195 ;
        RECT 136.715 216.785 136.900 216.865 ;
        RECT 125.195 215.725 125.965 215.945 ;
        RECT 125.175 214.815 125.515 215.545 ;
        RECT 125.695 214.995 125.965 215.725 ;
        RECT 126.145 215.705 127.305 215.945 ;
        RECT 126.145 214.995 126.375 215.705 ;
        RECT 126.545 214.815 126.875 215.525 ;
        RECT 127.045 214.995 127.305 215.705 ;
        RECT 127.505 215.765 128.090 215.955 ;
        RECT 127.505 214.995 127.780 215.765 ;
        RECT 128.260 215.595 129.155 215.925 ;
        RECT 130.255 215.905 131.005 216.425 ;
        RECT 132.565 216.125 132.900 216.395 ;
        RECT 133.070 216.005 133.240 216.565 ;
        RECT 133.410 216.125 133.745 216.375 ;
        RECT 133.935 216.075 135.145 216.595 ;
        RECT 127.950 215.425 129.155 215.595 ;
        RECT 127.950 214.995 128.280 215.425 ;
        RECT 128.450 214.815 128.645 215.255 ;
        RECT 128.825 214.995 129.155 215.425 ;
        RECT 129.335 214.815 131.005 215.905 ;
        RECT 131.635 214.815 131.925 215.980 ;
        RECT 133.070 215.965 133.245 216.005 ;
        RECT 132.555 214.815 132.835 215.955 ;
        RECT 133.005 214.985 133.335 215.965 ;
        RECT 133.505 214.815 133.765 215.955 ;
        RECT 135.315 215.905 136.525 216.425 ;
        RECT 133.935 214.815 136.525 215.905 ;
        RECT 136.715 215.655 136.885 216.785 ;
        RECT 137.685 216.715 137.855 216.945 ;
        RECT 137.055 216.545 137.855 216.715 ;
        RECT 137.055 215.995 137.225 216.545 ;
        RECT 138.035 216.375 138.320 216.775 ;
        RECT 137.455 216.345 137.820 216.375 ;
        RECT 137.445 216.175 137.820 216.345 ;
        RECT 137.990 216.175 138.320 216.375 ;
        RECT 138.590 216.375 138.870 216.775 ;
        RECT 139.050 216.715 139.220 216.945 ;
        RECT 139.445 216.885 139.775 217.365 ;
        RECT 139.945 216.715 140.115 217.195 ;
        RECT 139.050 216.545 140.115 216.715 ;
        RECT 140.380 216.690 140.655 217.035 ;
        RECT 140.845 216.965 141.225 217.365 ;
        RECT 141.395 216.795 141.565 217.145 ;
        RECT 141.735 216.965 142.065 217.365 ;
        RECT 142.235 216.795 142.490 217.145 ;
        RECT 142.675 216.820 148.020 217.365 ;
        RECT 138.590 216.175 139.065 216.375 ;
        RECT 139.235 216.175 139.680 216.375 ;
        RECT 139.850 216.165 140.200 216.375 ;
        RECT 137.055 215.825 140.115 215.995 ;
        RECT 136.715 214.985 136.970 215.655 ;
        RECT 137.140 214.815 137.470 215.575 ;
        RECT 137.640 215.415 139.275 215.655 ;
        RECT 137.640 214.985 137.890 215.415 ;
        RECT 139.045 215.325 139.275 215.415 ;
        RECT 138.060 214.815 138.415 215.235 ;
        RECT 138.605 215.155 138.935 215.195 ;
        RECT 139.445 215.155 139.775 215.655 ;
        RECT 138.605 214.985 139.775 215.155 ;
        RECT 139.945 214.985 140.115 215.825 ;
        RECT 140.380 215.955 140.550 216.690 ;
        RECT 140.825 216.625 142.490 216.795 ;
        RECT 140.825 216.455 140.995 216.625 ;
        RECT 140.720 216.125 140.995 216.455 ;
        RECT 141.165 216.125 141.990 216.455 ;
        RECT 142.160 216.125 142.505 216.455 ;
        RECT 140.825 215.955 140.995 216.125 ;
        RECT 140.380 214.985 140.655 215.955 ;
        RECT 140.825 215.785 141.485 215.955 ;
        RECT 141.795 215.835 141.990 216.125 ;
        RECT 144.260 215.990 144.600 216.820 ;
        RECT 148.195 216.595 149.865 217.365 ;
        RECT 141.315 215.665 141.485 215.785 ;
        RECT 142.160 215.665 142.485 215.955 ;
        RECT 140.865 214.815 141.145 215.615 ;
        RECT 141.315 215.495 142.485 215.665 ;
        RECT 141.315 215.035 142.505 215.325 ;
        RECT 146.080 215.250 146.430 216.500 ;
        RECT 148.195 216.075 148.945 216.595 ;
        RECT 149.115 215.905 149.865 216.425 ;
        RECT 142.675 214.815 148.020 215.250 ;
        RECT 148.195 214.815 149.865 215.905 ;
        RECT 150.495 216.420 150.835 217.195 ;
        RECT 151.005 216.905 151.175 217.365 ;
        RECT 151.415 216.930 151.775 217.195 ;
        RECT 151.415 216.925 151.770 216.930 ;
        RECT 151.415 216.915 151.765 216.925 ;
        RECT 151.415 216.910 151.760 216.915 ;
        RECT 151.415 216.900 151.755 216.910 ;
        RECT 152.405 216.905 152.575 217.365 ;
        RECT 151.415 216.895 151.750 216.900 ;
        RECT 151.415 216.885 151.740 216.895 ;
        RECT 151.415 216.875 151.730 216.885 ;
        RECT 151.415 216.735 151.715 216.875 ;
        RECT 151.005 216.545 151.715 216.735 ;
        RECT 151.905 216.735 152.235 216.815 ;
        RECT 152.745 216.735 153.085 217.195 ;
        RECT 151.905 216.545 153.085 216.735 ;
        RECT 153.255 216.865 153.555 217.195 ;
        RECT 153.725 216.885 154.000 217.365 ;
        RECT 150.495 214.985 150.775 216.420 ;
        RECT 151.005 215.975 151.290 216.545 ;
        RECT 151.475 216.145 151.945 216.375 ;
        RECT 152.115 216.355 152.445 216.375 ;
        RECT 152.115 216.175 152.565 216.355 ;
        RECT 152.755 216.175 153.085 216.375 ;
        RECT 151.005 215.760 152.155 215.975 ;
        RECT 150.945 214.815 151.655 215.590 ;
        RECT 151.825 214.985 152.155 215.760 ;
        RECT 152.350 215.060 152.565 216.175 ;
        RECT 152.855 215.835 153.085 216.175 ;
        RECT 153.255 215.955 153.425 216.865 ;
        RECT 154.180 216.715 154.475 217.105 ;
        RECT 154.645 216.885 154.900 217.365 ;
        RECT 155.075 216.715 155.335 217.105 ;
        RECT 155.505 216.885 155.785 217.365 ;
        RECT 153.595 216.125 153.945 216.695 ;
        RECT 154.180 216.545 155.830 216.715 ;
        RECT 156.935 216.615 158.145 217.365 ;
        RECT 154.115 216.205 155.255 216.375 ;
        RECT 154.115 215.955 154.285 216.205 ;
        RECT 155.425 216.035 155.830 216.545 ;
        RECT 153.255 215.785 154.285 215.955 ;
        RECT 155.075 215.865 155.830 216.035 ;
        RECT 156.935 215.905 157.455 216.445 ;
        RECT 157.625 216.075 158.145 216.615 ;
        RECT 152.745 214.815 153.075 215.535 ;
        RECT 153.255 214.985 153.565 215.785 ;
        RECT 155.075 215.615 155.335 215.865 ;
        RECT 153.735 214.815 154.045 215.615 ;
        RECT 154.215 215.445 155.335 215.615 ;
        RECT 154.215 214.985 154.475 215.445 ;
        RECT 154.645 214.815 154.900 215.275 ;
        RECT 155.075 214.985 155.335 215.445 ;
        RECT 155.505 214.815 155.790 215.685 ;
        RECT 156.935 214.815 158.145 215.905 ;
        RECT 2.750 214.645 158.230 214.815 ;
        RECT 2.835 213.555 4.045 214.645 ;
        RECT 2.835 212.845 3.355 213.385 ;
        RECT 3.525 213.015 4.045 213.555 ;
        RECT 4.765 213.715 4.935 214.475 ;
        RECT 5.115 213.885 5.445 214.645 ;
        RECT 4.765 213.545 5.430 213.715 ;
        RECT 5.615 213.570 5.885 214.475 ;
        RECT 5.260 213.400 5.430 213.545 ;
        RECT 4.695 212.995 5.025 213.365 ;
        RECT 5.260 213.070 5.545 213.400 ;
        RECT 2.835 212.095 4.045 212.845 ;
        RECT 5.260 212.815 5.430 213.070 ;
        RECT 4.765 212.645 5.430 212.815 ;
        RECT 5.715 212.770 5.885 213.570 ;
        RECT 4.765 212.265 4.935 212.645 ;
        RECT 5.115 212.095 5.445 212.475 ;
        RECT 5.625 212.265 5.885 212.770 ;
        RECT 6.060 213.505 6.395 214.475 ;
        RECT 6.565 213.505 6.735 214.645 ;
        RECT 6.905 214.305 8.935 214.475 ;
        RECT 6.060 212.835 6.230 213.505 ;
        RECT 6.905 213.335 7.075 214.305 ;
        RECT 6.400 213.005 6.655 213.335 ;
        RECT 6.880 213.005 7.075 213.335 ;
        RECT 7.245 213.965 8.370 214.135 ;
        RECT 6.485 212.835 6.655 213.005 ;
        RECT 7.245 212.835 7.415 213.965 ;
        RECT 6.060 212.265 6.315 212.835 ;
        RECT 6.485 212.665 7.415 212.835 ;
        RECT 7.585 213.625 8.595 213.795 ;
        RECT 7.585 212.825 7.755 213.625 ;
        RECT 7.960 213.285 8.235 213.425 ;
        RECT 7.955 213.115 8.235 213.285 ;
        RECT 7.240 212.630 7.415 212.665 ;
        RECT 6.485 212.095 6.815 212.495 ;
        RECT 7.240 212.265 7.770 212.630 ;
        RECT 7.960 212.265 8.235 213.115 ;
        RECT 8.405 212.265 8.595 213.625 ;
        RECT 8.765 213.640 8.935 214.305 ;
        RECT 9.105 213.885 9.275 214.645 ;
        RECT 9.510 213.885 10.025 214.295 ;
        RECT 8.765 213.450 9.515 213.640 ;
        RECT 9.685 213.075 10.025 213.885 ;
        RECT 8.795 212.905 10.025 213.075 ;
        RECT 10.200 213.505 10.535 214.475 ;
        RECT 10.705 213.505 10.875 214.645 ;
        RECT 11.045 214.305 13.075 214.475 ;
        RECT 8.775 212.095 9.285 212.630 ;
        RECT 9.505 212.300 9.750 212.905 ;
        RECT 10.200 212.835 10.370 213.505 ;
        RECT 11.045 213.335 11.215 214.305 ;
        RECT 10.540 213.005 10.795 213.335 ;
        RECT 11.020 213.005 11.215 213.335 ;
        RECT 11.385 213.965 12.510 214.135 ;
        RECT 10.625 212.835 10.795 213.005 ;
        RECT 11.385 212.835 11.555 213.965 ;
        RECT 10.200 212.265 10.455 212.835 ;
        RECT 10.625 212.665 11.555 212.835 ;
        RECT 11.725 213.625 12.735 213.795 ;
        RECT 11.725 212.825 11.895 213.625 ;
        RECT 12.100 212.945 12.375 213.425 ;
        RECT 12.095 212.775 12.375 212.945 ;
        RECT 11.380 212.630 11.555 212.665 ;
        RECT 10.625 212.095 10.955 212.495 ;
        RECT 11.380 212.265 11.910 212.630 ;
        RECT 12.100 212.265 12.375 212.775 ;
        RECT 12.545 212.265 12.735 213.625 ;
        RECT 12.905 213.640 13.075 214.305 ;
        RECT 13.245 213.885 13.415 214.645 ;
        RECT 13.650 213.885 14.165 214.295 ;
        RECT 12.905 213.450 13.655 213.640 ;
        RECT 13.825 213.075 14.165 213.885 ;
        RECT 12.935 212.905 14.165 213.075 ;
        RECT 14.335 213.570 14.605 214.475 ;
        RECT 14.775 213.885 15.105 214.645 ;
        RECT 15.285 213.715 15.455 214.475 ;
        RECT 12.915 212.095 13.425 212.630 ;
        RECT 13.645 212.300 13.890 212.905 ;
        RECT 14.335 212.770 14.505 213.570 ;
        RECT 14.790 213.545 15.455 213.715 ;
        RECT 14.790 213.400 14.960 213.545 ;
        RECT 15.715 213.480 16.005 214.645 ;
        RECT 16.180 213.975 16.435 214.475 ;
        RECT 16.605 214.145 16.935 214.645 ;
        RECT 16.180 213.805 16.930 213.975 ;
        RECT 14.675 213.070 14.960 213.400 ;
        RECT 14.790 212.815 14.960 213.070 ;
        RECT 15.195 212.995 15.525 213.365 ;
        RECT 16.180 212.985 16.530 213.635 ;
        RECT 14.335 212.265 14.595 212.770 ;
        RECT 14.790 212.645 15.455 212.815 ;
        RECT 14.775 212.095 15.105 212.475 ;
        RECT 15.285 212.265 15.455 212.645 ;
        RECT 15.715 212.095 16.005 212.820 ;
        RECT 16.700 212.815 16.930 213.805 ;
        RECT 16.180 212.645 16.930 212.815 ;
        RECT 16.180 212.355 16.435 212.645 ;
        RECT 16.605 212.095 16.935 212.475 ;
        RECT 17.105 212.355 17.275 214.475 ;
        RECT 17.445 213.675 17.770 214.460 ;
        RECT 17.940 214.185 18.190 214.645 ;
        RECT 18.360 214.145 18.610 214.475 ;
        RECT 18.825 214.145 19.505 214.475 ;
        RECT 18.360 214.015 18.530 214.145 ;
        RECT 18.135 213.845 18.530 214.015 ;
        RECT 17.505 212.625 17.965 213.675 ;
        RECT 18.135 212.485 18.305 213.845 ;
        RECT 18.700 213.585 19.165 213.975 ;
        RECT 18.475 212.775 18.825 213.395 ;
        RECT 18.995 212.995 19.165 213.585 ;
        RECT 19.335 213.365 19.505 214.145 ;
        RECT 19.675 214.045 19.845 214.385 ;
        RECT 20.080 214.215 20.410 214.645 ;
        RECT 20.580 214.045 20.750 214.385 ;
        RECT 21.045 214.185 21.415 214.645 ;
        RECT 19.675 213.875 20.750 214.045 ;
        RECT 21.585 214.015 21.755 214.475 ;
        RECT 21.990 214.135 22.860 214.475 ;
        RECT 23.030 214.185 23.280 214.645 ;
        RECT 21.195 213.845 21.755 214.015 ;
        RECT 21.195 213.705 21.365 213.845 ;
        RECT 19.865 213.535 21.365 213.705 ;
        RECT 22.060 213.675 22.520 213.965 ;
        RECT 19.335 213.195 21.025 213.365 ;
        RECT 18.995 212.775 19.350 212.995 ;
        RECT 19.520 212.485 19.690 213.195 ;
        RECT 19.895 212.775 20.685 213.025 ;
        RECT 20.855 213.015 21.025 213.195 ;
        RECT 21.195 212.845 21.365 213.535 ;
        RECT 17.635 212.095 17.965 212.455 ;
        RECT 18.135 212.315 18.630 212.485 ;
        RECT 18.835 212.315 19.690 212.485 ;
        RECT 20.565 212.095 20.895 212.555 ;
        RECT 21.105 212.455 21.365 212.845 ;
        RECT 21.555 213.665 22.520 213.675 ;
        RECT 22.690 213.755 22.860 214.135 ;
        RECT 23.450 214.095 23.620 214.385 ;
        RECT 23.800 214.265 24.130 214.645 ;
        RECT 23.450 213.925 24.250 214.095 ;
        RECT 21.555 213.505 22.230 213.665 ;
        RECT 22.690 213.585 23.910 213.755 ;
        RECT 21.555 212.715 21.765 213.505 ;
        RECT 22.690 213.495 22.860 213.585 ;
        RECT 21.935 212.715 22.285 213.335 ;
        RECT 22.455 213.325 22.860 213.495 ;
        RECT 22.455 212.545 22.625 213.325 ;
        RECT 22.795 212.875 23.015 213.155 ;
        RECT 23.195 213.045 23.735 213.415 ;
        RECT 24.080 213.305 24.250 213.925 ;
        RECT 24.425 213.585 24.595 214.645 ;
        RECT 24.805 213.635 25.095 214.475 ;
        RECT 25.265 213.805 25.435 214.645 ;
        RECT 25.645 213.635 25.895 214.475 ;
        RECT 26.105 213.805 26.275 214.645 ;
        RECT 27.985 213.805 28.155 214.645 ;
        RECT 28.365 213.635 28.615 214.475 ;
        RECT 28.825 213.805 28.995 214.645 ;
        RECT 29.165 213.635 29.455 214.475 ;
        RECT 24.805 213.465 26.530 213.635 ;
        RECT 22.795 212.705 23.325 212.875 ;
        RECT 21.105 212.285 21.455 212.455 ;
        RECT 21.675 212.265 22.625 212.545 ;
        RECT 22.795 212.095 22.985 212.535 ;
        RECT 23.155 212.475 23.325 212.705 ;
        RECT 23.495 212.645 23.735 213.045 ;
        RECT 23.905 213.295 24.250 213.305 ;
        RECT 23.905 213.085 25.935 213.295 ;
        RECT 23.905 212.830 24.230 213.085 ;
        RECT 26.120 212.915 26.530 213.465 ;
        RECT 23.905 212.475 24.225 212.830 ;
        RECT 23.155 212.305 24.225 212.475 ;
        RECT 24.425 212.095 24.595 212.905 ;
        RECT 24.765 212.745 26.530 212.915 ;
        RECT 27.730 213.465 29.455 213.635 ;
        RECT 29.665 213.585 29.835 214.645 ;
        RECT 30.130 214.265 30.460 214.645 ;
        RECT 30.640 214.095 30.810 214.385 ;
        RECT 30.980 214.185 31.230 214.645 ;
        RECT 30.010 213.925 30.810 214.095 ;
        RECT 31.400 214.135 32.270 214.475 ;
        RECT 27.730 212.915 28.140 213.465 ;
        RECT 30.010 213.305 30.180 213.925 ;
        RECT 31.400 213.755 31.570 214.135 ;
        RECT 32.505 214.015 32.675 214.475 ;
        RECT 32.845 214.185 33.215 214.645 ;
        RECT 33.510 214.045 33.680 214.385 ;
        RECT 33.850 214.215 34.180 214.645 ;
        RECT 34.415 214.045 34.585 214.385 ;
        RECT 30.350 213.585 31.570 213.755 ;
        RECT 31.740 213.675 32.200 213.965 ;
        RECT 32.505 213.845 33.065 214.015 ;
        RECT 33.510 213.875 34.585 214.045 ;
        RECT 34.755 214.145 35.435 214.475 ;
        RECT 35.650 214.145 35.900 214.475 ;
        RECT 36.070 214.185 36.320 214.645 ;
        RECT 32.895 213.705 33.065 213.845 ;
        RECT 31.740 213.665 32.705 213.675 ;
        RECT 31.400 213.495 31.570 213.585 ;
        RECT 32.030 213.505 32.705 213.665 ;
        RECT 30.010 213.295 30.355 213.305 ;
        RECT 28.325 213.085 30.355 213.295 ;
        RECT 27.730 212.745 29.495 212.915 ;
        RECT 24.765 212.265 25.095 212.745 ;
        RECT 25.265 212.095 25.435 212.565 ;
        RECT 25.605 212.265 25.935 212.745 ;
        RECT 26.105 212.095 26.275 212.565 ;
        RECT 27.985 212.095 28.155 212.565 ;
        RECT 28.325 212.265 28.655 212.745 ;
        RECT 28.825 212.095 28.995 212.565 ;
        RECT 29.165 212.265 29.495 212.745 ;
        RECT 29.665 212.095 29.835 212.905 ;
        RECT 30.030 212.830 30.355 213.085 ;
        RECT 30.035 212.475 30.355 212.830 ;
        RECT 30.525 213.045 31.065 213.415 ;
        RECT 31.400 213.325 31.805 213.495 ;
        RECT 30.525 212.645 30.765 213.045 ;
        RECT 31.245 212.875 31.465 213.155 ;
        RECT 30.935 212.705 31.465 212.875 ;
        RECT 30.935 212.475 31.105 212.705 ;
        RECT 31.635 212.545 31.805 213.325 ;
        RECT 31.975 212.715 32.325 213.335 ;
        RECT 32.495 212.715 32.705 213.505 ;
        RECT 32.895 213.535 34.395 213.705 ;
        RECT 32.895 212.845 33.065 213.535 ;
        RECT 34.755 213.365 34.925 214.145 ;
        RECT 35.730 214.015 35.900 214.145 ;
        RECT 33.235 213.195 34.925 213.365 ;
        RECT 35.095 213.585 35.560 213.975 ;
        RECT 35.730 213.845 36.125 214.015 ;
        RECT 33.235 213.015 33.405 213.195 ;
        RECT 30.035 212.305 31.105 212.475 ;
        RECT 31.275 212.095 31.465 212.535 ;
        RECT 31.635 212.265 32.585 212.545 ;
        RECT 32.895 212.455 33.155 212.845 ;
        RECT 33.575 212.775 34.365 213.025 ;
        RECT 32.805 212.285 33.155 212.455 ;
        RECT 33.365 212.095 33.695 212.555 ;
        RECT 34.570 212.485 34.740 213.195 ;
        RECT 35.095 212.995 35.265 213.585 ;
        RECT 34.910 212.775 35.265 212.995 ;
        RECT 35.435 212.775 35.785 213.395 ;
        RECT 35.955 212.485 36.125 213.845 ;
        RECT 36.490 213.675 36.815 214.460 ;
        RECT 36.295 212.625 36.755 213.675 ;
        RECT 34.570 212.315 35.425 212.485 ;
        RECT 35.630 212.315 36.125 212.485 ;
        RECT 36.295 212.095 36.625 212.455 ;
        RECT 36.985 212.355 37.155 214.475 ;
        RECT 37.325 214.145 37.655 214.645 ;
        RECT 37.825 213.975 38.080 214.475 ;
        RECT 37.330 213.805 38.080 213.975 ;
        RECT 37.330 212.815 37.560 213.805 ;
        RECT 38.770 213.775 39.055 214.645 ;
        RECT 39.225 214.015 39.485 214.475 ;
        RECT 39.660 214.185 39.915 214.645 ;
        RECT 40.085 214.015 40.345 214.475 ;
        RECT 39.225 213.845 40.345 214.015 ;
        RECT 40.515 213.845 40.825 214.645 ;
        RECT 37.730 212.985 38.080 213.635 ;
        RECT 39.225 213.595 39.485 213.845 ;
        RECT 40.995 213.675 41.305 214.475 ;
        RECT 38.730 213.425 39.485 213.595 ;
        RECT 40.275 213.505 41.305 213.675 ;
        RECT 38.730 212.915 39.135 213.425 ;
        RECT 40.275 213.255 40.445 213.505 ;
        RECT 39.305 213.085 40.445 213.255 ;
        RECT 37.330 212.645 38.080 212.815 ;
        RECT 38.730 212.745 40.380 212.915 ;
        RECT 40.615 212.765 40.965 213.335 ;
        RECT 37.325 212.095 37.655 212.475 ;
        RECT 37.825 212.355 38.080 212.645 ;
        RECT 38.775 212.095 39.055 212.575 ;
        RECT 39.225 212.355 39.485 212.745 ;
        RECT 39.660 212.095 39.915 212.575 ;
        RECT 40.085 212.355 40.380 212.745 ;
        RECT 41.135 212.595 41.305 213.505 ;
        RECT 41.475 213.480 41.765 214.645 ;
        RECT 41.990 213.775 42.275 214.645 ;
        RECT 42.445 214.015 42.705 214.475 ;
        RECT 42.880 214.185 43.135 214.645 ;
        RECT 43.305 214.015 43.565 214.475 ;
        RECT 42.445 213.845 43.565 214.015 ;
        RECT 43.735 213.845 44.045 214.645 ;
        RECT 42.445 213.595 42.705 213.845 ;
        RECT 44.215 213.675 44.525 214.475 ;
        RECT 41.950 213.425 42.705 213.595 ;
        RECT 43.495 213.505 44.525 213.675 ;
        RECT 41.950 212.915 42.355 213.425 ;
        RECT 43.495 213.255 43.665 213.505 ;
        RECT 42.525 213.085 43.665 213.255 ;
        RECT 40.560 212.095 40.835 212.575 ;
        RECT 41.005 212.265 41.305 212.595 ;
        RECT 41.475 212.095 41.765 212.820 ;
        RECT 41.950 212.745 43.600 212.915 ;
        RECT 43.835 212.765 44.185 213.335 ;
        RECT 41.995 212.095 42.275 212.575 ;
        RECT 42.445 212.355 42.705 212.745 ;
        RECT 42.880 212.095 43.135 212.575 ;
        RECT 43.305 212.355 43.600 212.745 ;
        RECT 44.355 212.595 44.525 213.505 ;
        RECT 43.780 212.095 44.055 212.575 ;
        RECT 44.225 212.265 44.525 212.595 ;
        RECT 44.700 213.505 45.035 214.475 ;
        RECT 45.205 213.505 45.375 214.645 ;
        RECT 45.545 214.305 47.575 214.475 ;
        RECT 44.700 212.835 44.870 213.505 ;
        RECT 45.545 213.335 45.715 214.305 ;
        RECT 45.040 213.005 45.295 213.335 ;
        RECT 45.520 213.005 45.715 213.335 ;
        RECT 45.885 213.965 47.010 214.135 ;
        RECT 45.125 212.835 45.295 213.005 ;
        RECT 45.885 212.835 46.055 213.965 ;
        RECT 44.700 212.265 44.955 212.835 ;
        RECT 45.125 212.665 46.055 212.835 ;
        RECT 46.225 213.625 47.235 213.795 ;
        RECT 46.225 212.825 46.395 213.625 ;
        RECT 46.600 212.945 46.875 213.425 ;
        RECT 46.595 212.775 46.875 212.945 ;
        RECT 45.880 212.630 46.055 212.665 ;
        RECT 45.125 212.095 45.455 212.495 ;
        RECT 45.880 212.265 46.410 212.630 ;
        RECT 46.600 212.265 46.875 212.775 ;
        RECT 47.045 212.265 47.235 213.625 ;
        RECT 47.405 213.640 47.575 214.305 ;
        RECT 47.745 213.885 47.915 214.645 ;
        RECT 48.150 213.885 48.665 214.295 ;
        RECT 47.405 213.450 48.155 213.640 ;
        RECT 48.325 213.075 48.665 213.885 ;
        RECT 47.435 212.905 48.665 213.075 ;
        RECT 48.835 213.885 49.350 214.295 ;
        RECT 49.585 213.885 49.755 214.645 ;
        RECT 49.925 214.305 51.955 214.475 ;
        RECT 48.835 213.075 49.175 213.885 ;
        RECT 49.925 213.640 50.095 214.305 ;
        RECT 50.490 213.965 51.615 214.135 ;
        RECT 49.345 213.450 50.095 213.640 ;
        RECT 50.265 213.625 51.275 213.795 ;
        RECT 48.835 212.905 50.065 213.075 ;
        RECT 47.415 212.095 47.925 212.630 ;
        RECT 48.145 212.300 48.390 212.905 ;
        RECT 49.110 212.300 49.355 212.905 ;
        RECT 49.575 212.095 50.085 212.630 ;
        RECT 50.265 212.265 50.455 213.625 ;
        RECT 50.625 212.605 50.900 213.425 ;
        RECT 51.105 212.825 51.275 213.625 ;
        RECT 51.445 212.835 51.615 213.965 ;
        RECT 51.785 213.335 51.955 214.305 ;
        RECT 52.125 213.505 52.295 214.645 ;
        RECT 52.465 213.505 52.800 214.475 ;
        RECT 53.950 213.775 54.235 214.645 ;
        RECT 54.405 214.015 54.665 214.475 ;
        RECT 54.840 214.185 55.095 214.645 ;
        RECT 55.265 214.015 55.525 214.475 ;
        RECT 54.405 213.845 55.525 214.015 ;
        RECT 55.695 213.845 56.005 214.645 ;
        RECT 54.405 213.595 54.665 213.845 ;
        RECT 56.175 213.675 56.485 214.475 ;
        RECT 51.785 213.005 51.980 213.335 ;
        RECT 52.205 213.005 52.460 213.335 ;
        RECT 52.205 212.835 52.375 213.005 ;
        RECT 52.630 212.835 52.800 213.505 ;
        RECT 51.445 212.665 52.375 212.835 ;
        RECT 51.445 212.630 51.620 212.665 ;
        RECT 50.625 212.435 50.905 212.605 ;
        RECT 50.625 212.265 50.900 212.435 ;
        RECT 51.090 212.265 51.620 212.630 ;
        RECT 52.045 212.095 52.375 212.495 ;
        RECT 52.545 212.265 52.800 212.835 ;
        RECT 53.910 213.425 54.665 213.595 ;
        RECT 55.455 213.505 56.485 213.675 ;
        RECT 57.030 213.665 57.285 214.335 ;
        RECT 57.465 213.845 57.750 214.645 ;
        RECT 57.930 213.925 58.260 214.435 ;
        RECT 57.030 213.625 57.210 213.665 ;
        RECT 53.910 212.915 54.315 213.425 ;
        RECT 55.455 213.255 55.625 213.505 ;
        RECT 54.485 213.085 55.625 213.255 ;
        RECT 53.910 212.745 55.560 212.915 ;
        RECT 55.795 212.765 56.145 213.335 ;
        RECT 53.955 212.095 54.235 212.575 ;
        RECT 54.405 212.355 54.665 212.745 ;
        RECT 54.840 212.095 55.095 212.575 ;
        RECT 55.265 212.355 55.560 212.745 ;
        RECT 56.315 212.595 56.485 213.505 ;
        RECT 56.945 213.455 57.210 213.625 ;
        RECT 55.740 212.095 56.015 212.575 ;
        RECT 56.185 212.265 56.485 212.595 ;
        RECT 57.030 212.805 57.210 213.455 ;
        RECT 57.930 213.335 58.180 213.925 ;
        RECT 58.530 213.775 58.700 214.385 ;
        RECT 58.870 213.955 59.200 214.645 ;
        RECT 59.430 214.095 59.670 214.385 ;
        RECT 59.870 214.265 60.290 214.645 ;
        RECT 60.470 214.175 61.100 214.425 ;
        RECT 61.570 214.265 61.900 214.645 ;
        RECT 60.470 214.095 60.640 214.175 ;
        RECT 62.070 214.095 62.240 214.385 ;
        RECT 62.420 214.265 62.800 214.645 ;
        RECT 63.040 214.260 63.870 214.430 ;
        RECT 59.430 213.925 60.640 214.095 ;
        RECT 57.380 213.005 58.180 213.335 ;
        RECT 57.030 212.275 57.285 212.805 ;
        RECT 57.465 212.095 57.750 212.555 ;
        RECT 57.930 212.355 58.180 213.005 ;
        RECT 58.380 213.755 58.700 213.775 ;
        RECT 58.380 213.585 60.300 213.755 ;
        RECT 58.380 212.690 58.570 213.585 ;
        RECT 60.470 213.415 60.640 213.925 ;
        RECT 60.810 213.665 61.330 213.975 ;
        RECT 58.740 213.245 60.640 213.415 ;
        RECT 58.740 213.185 59.070 213.245 ;
        RECT 59.220 213.015 59.550 213.075 ;
        RECT 58.890 212.745 59.550 213.015 ;
        RECT 58.380 212.360 58.700 212.690 ;
        RECT 58.880 212.095 59.540 212.575 ;
        RECT 59.740 212.485 59.910 213.245 ;
        RECT 60.810 213.075 60.990 213.485 ;
        RECT 60.080 212.905 60.410 213.025 ;
        RECT 61.160 212.905 61.330 213.665 ;
        RECT 60.080 212.735 61.330 212.905 ;
        RECT 61.500 213.845 62.870 214.095 ;
        RECT 61.500 213.075 61.690 213.845 ;
        RECT 62.620 213.585 62.870 213.845 ;
        RECT 61.860 213.415 62.110 213.575 ;
        RECT 63.040 213.415 63.210 214.260 ;
        RECT 64.105 213.975 64.275 214.475 ;
        RECT 64.445 214.145 64.775 214.645 ;
        RECT 63.380 213.585 63.880 213.965 ;
        RECT 64.105 213.805 64.800 213.975 ;
        RECT 61.860 213.245 63.210 213.415 ;
        RECT 62.790 213.205 63.210 213.245 ;
        RECT 61.500 212.735 61.920 213.075 ;
        RECT 62.210 212.745 62.620 213.075 ;
        RECT 59.740 212.315 60.590 212.485 ;
        RECT 61.150 212.095 61.470 212.555 ;
        RECT 61.670 212.305 61.920 212.735 ;
        RECT 62.210 212.095 62.620 212.535 ;
        RECT 62.790 212.475 62.960 213.205 ;
        RECT 63.130 212.655 63.480 213.025 ;
        RECT 63.660 212.715 63.880 213.585 ;
        RECT 64.050 213.015 64.460 213.635 ;
        RECT 64.630 212.835 64.800 213.805 ;
        RECT 64.105 212.645 64.800 212.835 ;
        RECT 62.790 212.275 63.805 212.475 ;
        RECT 64.105 212.315 64.275 212.645 ;
        RECT 64.445 212.095 64.775 212.475 ;
        RECT 64.990 212.355 65.215 214.475 ;
        RECT 65.385 214.145 65.715 214.645 ;
        RECT 65.885 213.975 66.055 214.475 ;
        RECT 65.390 213.805 66.055 213.975 ;
        RECT 65.390 212.815 65.620 213.805 ;
        RECT 65.790 212.985 66.140 213.635 ;
        RECT 67.235 213.480 67.525 214.645 ;
        RECT 67.735 213.505 67.965 214.645 ;
        RECT 68.135 213.495 68.465 214.475 ;
        RECT 68.635 213.505 68.845 214.645 ;
        RECT 69.075 213.555 70.285 214.645 ;
        RECT 67.715 213.085 68.045 213.335 ;
        RECT 65.390 212.645 66.055 212.815 ;
        RECT 65.385 212.095 65.715 212.475 ;
        RECT 65.885 212.355 66.055 212.645 ;
        RECT 67.235 212.095 67.525 212.820 ;
        RECT 67.735 212.095 67.965 212.915 ;
        RECT 68.215 212.895 68.465 213.495 ;
        RECT 68.135 212.265 68.465 212.895 ;
        RECT 68.635 212.095 68.845 212.915 ;
        RECT 69.075 212.845 69.595 213.385 ;
        RECT 69.765 213.015 70.285 213.555 ;
        RECT 70.455 214.175 70.795 214.435 ;
        RECT 70.965 214.185 71.215 214.645 ;
        RECT 69.075 212.095 70.285 212.845 ;
        RECT 70.455 212.570 70.715 214.175 ;
        RECT 71.405 214.005 71.735 214.435 ;
        RECT 70.885 213.835 71.735 214.005 ;
        RECT 71.905 213.975 72.075 214.475 ;
        RECT 72.285 214.185 72.535 214.645 ;
        RECT 72.745 213.975 72.915 214.475 ;
        RECT 73.215 214.185 73.465 214.645 ;
        RECT 73.705 213.975 73.875 214.475 ;
        RECT 70.885 212.915 71.055 213.835 ;
        RECT 71.905 213.805 73.875 213.975 ;
        RECT 71.375 213.085 71.705 213.645 ;
        RECT 71.905 213.335 72.205 213.630 ;
        RECT 71.905 213.285 72.285 213.335 ;
        RECT 71.895 213.115 72.285 213.285 ;
        RECT 71.905 213.005 72.285 213.115 ;
        RECT 70.885 212.820 71.705 212.915 ;
        RECT 70.885 212.745 71.900 212.820 ;
        RECT 70.455 212.310 70.795 212.570 ;
        RECT 70.965 212.095 71.295 212.575 ;
        RECT 71.485 212.310 71.900 212.745 ;
        RECT 72.595 212.610 72.815 213.335 ;
        RECT 73.075 213.005 73.455 213.635 ;
        RECT 73.685 213.005 73.940 213.635 ;
        RECT 74.135 213.505 74.395 214.645 ;
        RECT 74.565 213.495 74.895 214.475 ;
        RECT 75.065 213.505 75.345 214.645 ;
        RECT 75.515 213.555 77.185 214.645 ;
        RECT 74.155 213.085 74.490 213.335 ;
        RECT 72.070 212.425 73.020 212.610 ;
        RECT 73.250 212.405 73.455 213.005 ;
        RECT 74.660 212.895 74.830 213.495 ;
        RECT 75.000 213.065 75.335 213.335 ;
        RECT 73.625 212.095 73.965 212.820 ;
        RECT 74.135 212.265 74.830 212.895 ;
        RECT 75.035 212.095 75.345 212.895 ;
        RECT 75.515 212.865 76.265 213.385 ;
        RECT 76.435 213.035 77.185 213.555 ;
        RECT 77.355 213.505 77.615 214.645 ;
        RECT 77.785 213.495 78.115 214.475 ;
        RECT 78.285 213.505 78.565 214.645 ;
        RECT 78.740 214.265 79.075 214.645 ;
        RECT 77.375 213.085 77.710 213.335 ;
        RECT 77.880 212.895 78.050 213.495 ;
        RECT 78.220 213.065 78.555 213.335 ;
        RECT 75.515 212.095 77.185 212.865 ;
        RECT 77.355 212.265 78.050 212.895 ;
        RECT 78.255 212.095 78.565 212.895 ;
        RECT 78.735 212.775 78.975 214.085 ;
        RECT 79.245 213.675 79.495 214.475 ;
        RECT 79.715 213.925 80.045 214.645 ;
        RECT 80.230 213.675 80.480 214.475 ;
        RECT 80.945 213.845 81.275 214.645 ;
        RECT 81.445 214.215 81.785 214.475 ;
        RECT 79.145 213.505 81.335 213.675 ;
        RECT 79.145 212.595 79.315 213.505 ;
        RECT 81.020 213.335 81.335 213.505 ;
        RECT 78.820 212.265 79.315 212.595 ;
        RECT 79.535 212.370 79.885 213.335 ;
        RECT 80.065 212.365 80.365 213.335 ;
        RECT 80.545 212.365 80.825 213.335 ;
        RECT 81.020 213.085 81.350 213.335 ;
        RECT 81.005 212.095 81.275 212.895 ;
        RECT 81.525 212.815 81.785 214.215 ;
        RECT 81.965 213.505 82.295 214.645 ;
        RECT 82.825 213.675 83.155 214.460 ;
        RECT 82.475 213.505 83.155 213.675 ;
        RECT 83.795 213.505 84.055 214.645 ;
        RECT 81.955 213.085 82.305 213.335 ;
        RECT 82.475 212.905 82.645 213.505 ;
        RECT 84.225 213.495 84.555 214.475 ;
        RECT 84.725 213.505 85.005 214.645 ;
        RECT 85.185 213.585 85.515 214.435 ;
        RECT 82.815 213.085 83.165 213.335 ;
        RECT 83.815 213.085 84.150 213.335 ;
        RECT 81.445 212.305 81.785 212.815 ;
        RECT 81.965 212.095 82.235 212.905 ;
        RECT 82.405 212.265 82.735 212.905 ;
        RECT 82.905 212.095 83.145 212.905 ;
        RECT 84.320 212.895 84.490 213.495 ;
        RECT 84.660 213.065 84.995 213.335 ;
        RECT 83.795 212.265 84.490 212.895 ;
        RECT 84.695 212.095 85.005 212.895 ;
        RECT 85.185 212.820 85.375 213.585 ;
        RECT 85.685 213.505 85.935 214.645 ;
        RECT 86.125 214.005 86.375 214.425 ;
        RECT 86.605 214.175 86.935 214.645 ;
        RECT 87.165 214.005 87.415 214.425 ;
        RECT 86.125 213.835 87.415 214.005 ;
        RECT 87.595 214.005 87.925 214.435 ;
        RECT 87.595 213.835 88.050 214.005 ;
        RECT 86.115 213.335 86.330 213.665 ;
        RECT 85.545 213.005 85.855 213.335 ;
        RECT 86.025 213.005 86.330 213.335 ;
        RECT 86.505 213.005 86.790 213.665 ;
        RECT 86.985 213.005 87.250 213.665 ;
        RECT 87.465 213.005 87.710 213.665 ;
        RECT 85.685 212.835 85.855 213.005 ;
        RECT 87.880 212.835 88.050 213.835 ;
        RECT 85.185 212.310 85.515 212.820 ;
        RECT 85.685 212.665 88.050 212.835 ;
        RECT 88.395 213.775 88.670 214.475 ;
        RECT 88.840 214.100 89.095 214.645 ;
        RECT 89.265 214.135 89.745 214.475 ;
        RECT 89.920 214.090 90.525 214.645 ;
        RECT 89.910 213.990 90.525 214.090 ;
        RECT 89.910 213.965 90.095 213.990 ;
        RECT 88.395 212.745 88.565 213.775 ;
        RECT 88.840 213.645 89.595 213.895 ;
        RECT 89.765 213.720 90.095 213.965 ;
        RECT 88.840 213.610 89.610 213.645 ;
        RECT 88.840 213.600 89.625 213.610 ;
        RECT 88.735 213.585 89.630 213.600 ;
        RECT 88.735 213.570 89.650 213.585 ;
        RECT 88.735 213.560 89.670 213.570 ;
        RECT 88.735 213.550 89.695 213.560 ;
        RECT 88.735 213.520 89.765 213.550 ;
        RECT 88.735 213.490 89.785 213.520 ;
        RECT 88.735 213.460 89.805 213.490 ;
        RECT 88.735 213.435 89.835 213.460 ;
        RECT 88.735 213.400 89.870 213.435 ;
        RECT 88.735 213.395 89.900 213.400 ;
        RECT 88.735 213.000 88.965 213.395 ;
        RECT 89.510 213.390 89.900 213.395 ;
        RECT 89.535 213.380 89.900 213.390 ;
        RECT 89.550 213.375 89.900 213.380 ;
        RECT 89.565 213.370 89.900 213.375 ;
        RECT 90.265 213.370 90.525 213.820 ;
        RECT 90.695 213.555 92.365 214.645 ;
        RECT 89.565 213.365 90.525 213.370 ;
        RECT 89.575 213.355 90.525 213.365 ;
        RECT 89.585 213.350 90.525 213.355 ;
        RECT 89.595 213.340 90.525 213.350 ;
        RECT 89.600 213.330 90.525 213.340 ;
        RECT 89.605 213.325 90.525 213.330 ;
        RECT 89.615 213.310 90.525 213.325 ;
        RECT 89.620 213.295 90.525 213.310 ;
        RECT 89.630 213.270 90.525 213.295 ;
        RECT 89.135 212.800 89.465 213.225 ;
        RECT 85.685 212.095 86.015 212.495 ;
        RECT 87.065 212.325 87.395 212.665 ;
        RECT 87.565 212.095 87.895 212.495 ;
        RECT 88.395 212.265 88.655 212.745 ;
        RECT 88.825 212.095 89.075 212.635 ;
        RECT 89.245 212.315 89.465 212.800 ;
        RECT 89.635 213.200 90.525 213.270 ;
        RECT 89.635 212.475 89.805 213.200 ;
        RECT 89.975 212.645 90.525 213.030 ;
        RECT 90.695 212.865 91.445 213.385 ;
        RECT 91.615 213.035 92.365 213.555 ;
        RECT 92.995 213.480 93.285 214.645 ;
        RECT 93.455 214.210 98.800 214.645 ;
        RECT 89.635 212.305 90.525 212.475 ;
        RECT 90.695 212.095 92.365 212.865 ;
        RECT 92.995 212.095 93.285 212.820 ;
        RECT 95.040 212.640 95.380 213.470 ;
        RECT 96.860 212.960 97.210 214.210 ;
        RECT 99.895 213.845 100.335 214.475 ;
        RECT 99.895 212.835 100.205 213.845 ;
        RECT 100.510 213.795 100.825 214.645 ;
        RECT 100.995 214.305 102.425 214.475 ;
        RECT 100.995 213.625 101.165 214.305 ;
        RECT 100.375 213.455 101.165 213.625 ;
        RECT 100.375 213.005 100.545 213.455 ;
        RECT 101.335 213.335 101.535 214.135 ;
        RECT 100.715 213.005 101.105 213.285 ;
        RECT 101.290 213.005 101.535 213.335 ;
        RECT 101.735 213.005 101.985 214.135 ;
        RECT 102.175 213.675 102.425 214.305 ;
        RECT 102.605 213.845 102.935 214.645 ;
        RECT 102.175 213.505 102.945 213.675 ;
        RECT 103.115 213.555 104.325 214.645 ;
        RECT 102.200 213.005 102.605 213.335 ;
        RECT 102.775 212.835 102.945 213.505 ;
        RECT 93.455 212.095 98.800 212.640 ;
        RECT 99.895 212.275 100.335 212.835 ;
        RECT 100.505 212.095 100.955 212.835 ;
        RECT 101.125 212.665 102.285 212.835 ;
        RECT 101.125 212.265 101.295 212.665 ;
        RECT 101.465 212.095 101.885 212.495 ;
        RECT 102.055 212.265 102.285 212.665 ;
        RECT 102.455 212.265 102.945 212.835 ;
        RECT 103.115 212.845 103.635 213.385 ;
        RECT 103.805 213.015 104.325 213.555 ;
        RECT 104.495 213.505 104.835 214.475 ;
        RECT 105.005 213.505 105.175 214.645 ;
        RECT 105.445 213.845 105.695 214.645 ;
        RECT 106.340 213.675 106.670 214.475 ;
        RECT 106.970 213.845 107.300 214.645 ;
        RECT 107.470 213.675 107.800 214.475 ;
        RECT 105.365 213.505 107.800 213.675 ;
        RECT 108.175 213.555 110.765 214.645 ;
        RECT 104.495 212.945 104.670 213.505 ;
        RECT 105.365 213.255 105.535 213.505 ;
        RECT 104.840 213.085 105.535 213.255 ;
        RECT 105.710 213.085 106.130 213.285 ;
        RECT 106.300 213.085 106.630 213.285 ;
        RECT 106.800 213.085 107.130 213.285 ;
        RECT 104.495 212.895 104.725 212.945 ;
        RECT 103.115 212.095 104.325 212.845 ;
        RECT 104.495 212.265 104.835 212.895 ;
        RECT 105.005 212.095 105.255 212.895 ;
        RECT 105.445 212.745 106.670 212.915 ;
        RECT 105.445 212.265 105.775 212.745 ;
        RECT 105.945 212.095 106.170 212.555 ;
        RECT 106.340 212.265 106.670 212.745 ;
        RECT 107.300 212.875 107.470 213.505 ;
        RECT 107.655 213.085 108.005 213.335 ;
        RECT 107.300 212.265 107.800 212.875 ;
        RECT 108.175 212.865 109.385 213.385 ;
        RECT 109.555 213.035 110.765 213.555 ;
        RECT 111.100 213.735 111.350 214.465 ;
        RECT 111.520 213.915 111.850 214.645 ;
        RECT 112.020 213.735 112.205 214.465 ;
        RECT 111.100 213.535 112.205 213.735 ;
        RECT 112.375 213.335 112.605 214.465 ;
        RECT 112.785 213.795 113.510 214.465 ;
        RECT 108.175 212.095 110.765 212.865 ;
        RECT 110.945 212.775 111.285 213.335 ;
        RECT 111.455 213.005 112.095 213.335 ;
        RECT 112.275 213.005 112.605 213.335 ;
        RECT 112.785 213.005 113.085 213.625 ;
        RECT 110.935 212.095 111.275 212.605 ;
        RECT 111.455 212.275 111.705 213.005 ;
        RECT 113.295 212.825 113.510 213.795 ;
        RECT 113.695 213.555 117.205 214.645 ;
        RECT 117.375 213.555 118.585 214.645 ;
        RECT 112.030 212.635 113.510 212.825 ;
        RECT 113.695 212.865 115.345 213.385 ;
        RECT 115.515 213.035 117.205 213.555 ;
        RECT 112.030 212.275 112.215 212.635 ;
        RECT 112.395 212.095 112.725 212.465 ;
        RECT 112.905 212.275 113.130 212.635 ;
        RECT 113.695 212.095 117.205 212.865 ;
        RECT 117.375 212.845 117.895 213.385 ;
        RECT 118.065 213.015 118.585 213.555 ;
        RECT 118.755 213.480 119.045 214.645 ;
        RECT 119.215 213.555 122.725 214.645 ;
        RECT 119.215 212.865 120.865 213.385 ;
        RECT 121.035 213.035 122.725 213.555 ;
        RECT 122.900 213.505 123.220 214.645 ;
        RECT 123.400 213.335 123.595 214.385 ;
        RECT 123.775 213.795 124.105 214.475 ;
        RECT 124.305 213.845 124.560 214.645 ;
        RECT 124.735 214.210 130.080 214.645 ;
        RECT 123.775 213.515 124.125 213.795 ;
        RECT 122.960 213.005 123.220 213.335 ;
        RECT 123.400 213.005 123.785 213.335 ;
        RECT 123.955 213.135 124.125 213.515 ;
        RECT 124.315 213.305 124.560 213.665 ;
        RECT 123.955 212.965 124.475 213.135 ;
        RECT 117.375 212.095 118.585 212.845 ;
        RECT 118.755 212.095 119.045 212.820 ;
        RECT 119.215 212.095 122.725 212.865 ;
        RECT 122.900 212.625 124.115 212.795 ;
        RECT 122.900 212.275 123.190 212.625 ;
        RECT 123.385 212.095 123.715 212.455 ;
        RECT 123.885 212.320 124.115 212.625 ;
        RECT 124.305 212.400 124.475 212.965 ;
        RECT 126.320 212.640 126.660 213.470 ;
        RECT 128.140 212.960 128.490 214.210 ;
        RECT 130.255 213.555 133.765 214.645 ;
        RECT 130.255 212.865 131.905 213.385 ;
        RECT 132.075 213.035 133.765 213.555 ;
        RECT 134.420 213.420 134.675 214.645 ;
        RECT 134.845 213.805 135.100 214.475 ;
        RECT 135.270 214.245 135.600 214.645 ;
        RECT 136.470 214.245 136.875 214.645 ;
        RECT 137.145 214.065 137.495 214.435 ;
        RECT 135.410 213.895 137.495 214.065 ;
        RECT 124.735 212.095 130.080 212.640 ;
        RECT 130.255 212.095 133.765 212.865 ;
        RECT 134.420 212.095 134.675 212.920 ;
        RECT 134.845 212.835 135.015 213.805 ;
        RECT 135.410 213.625 135.580 213.895 ;
        RECT 135.185 213.455 135.580 213.625 ;
        RECT 135.750 213.505 136.770 213.725 ;
        RECT 135.185 213.005 135.355 213.455 ;
        RECT 136.505 213.365 136.770 213.505 ;
        RECT 136.940 213.505 137.495 213.895 ;
        RECT 135.525 213.085 135.995 213.285 ;
        RECT 136.165 212.915 136.335 213.110 ;
        RECT 134.845 212.265 135.180 212.835 ;
        RECT 135.825 212.780 136.335 212.915 ;
        RECT 135.375 212.095 135.545 212.760 ;
        RECT 135.825 212.745 136.330 212.780 ;
        RECT 135.825 212.390 136.045 212.745 ;
        RECT 136.505 212.575 136.675 213.365 ;
        RECT 136.940 213.255 137.110 213.505 ;
        RECT 137.665 213.335 137.835 214.435 ;
        RECT 138.040 213.825 138.355 214.645 ;
        RECT 138.535 214.210 143.880 214.645 ;
        RECT 136.920 213.085 137.110 213.255 ;
        RECT 137.280 213.085 137.835 213.335 ;
        RECT 138.010 213.085 138.355 213.655 ;
        RECT 136.920 212.700 137.090 213.085 ;
        RECT 136.215 212.405 136.675 212.575 ;
        RECT 136.845 212.330 137.090 212.700 ;
        RECT 137.265 212.735 138.355 212.915 ;
        RECT 137.265 212.330 137.495 212.735 ;
        RECT 137.685 212.095 137.855 212.565 ;
        RECT 138.025 212.330 138.355 212.735 ;
        RECT 140.120 212.640 140.460 213.470 ;
        RECT 141.940 212.960 142.290 214.210 ;
        RECT 144.515 213.480 144.805 214.645 ;
        RECT 144.985 213.505 145.315 214.645 ;
        RECT 145.490 213.755 145.660 214.315 ;
        RECT 145.830 213.925 146.090 214.645 ;
        RECT 146.260 214.185 146.590 214.355 ;
        RECT 146.260 213.755 146.430 214.185 ;
        RECT 146.840 214.015 147.120 214.365 ;
        RECT 145.490 213.585 146.430 213.755 ;
        RECT 146.600 213.845 147.120 214.015 ;
        RECT 144.980 212.985 145.310 213.335 ;
        RECT 145.490 213.005 145.915 213.335 ;
        RECT 146.085 213.005 146.345 213.335 ;
        RECT 146.600 213.005 146.825 213.845 ;
        RECT 147.300 213.675 147.540 214.345 ;
        RECT 146.995 213.505 147.540 213.675 ;
        RECT 148.195 213.675 148.505 214.475 ;
        RECT 148.675 213.845 148.985 214.645 ;
        RECT 149.155 214.015 149.415 214.475 ;
        RECT 149.585 214.185 149.840 214.645 ;
        RECT 150.015 214.015 150.275 214.475 ;
        RECT 149.155 213.845 150.275 214.015 ;
        RECT 148.195 213.505 149.225 213.675 ;
        RECT 138.535 212.095 143.880 212.640 ;
        RECT 144.515 212.095 144.805 212.820 ;
        RECT 144.985 212.095 145.315 212.815 ;
        RECT 145.490 212.275 145.685 213.005 ;
        RECT 146.085 212.670 146.255 213.005 ;
        RECT 146.995 212.835 147.165 213.505 ;
        RECT 147.335 213.005 147.575 213.335 ;
        RECT 145.855 212.275 146.255 212.670 ;
        RECT 146.425 212.665 147.540 212.835 ;
        RECT 146.425 212.265 146.595 212.665 ;
        RECT 146.795 212.095 147.125 212.495 ;
        RECT 147.295 212.305 147.540 212.665 ;
        RECT 148.195 212.595 148.365 213.505 ;
        RECT 148.535 212.765 148.885 213.335 ;
        RECT 149.055 213.255 149.225 213.505 ;
        RECT 150.015 213.595 150.275 213.845 ;
        RECT 150.445 213.775 150.730 214.645 ;
        RECT 150.015 213.425 150.770 213.595 ;
        RECT 150.955 213.555 152.165 214.645 ;
        RECT 152.375 214.305 153.515 214.475 ;
        RECT 152.375 213.845 152.675 214.305 ;
        RECT 152.845 213.675 153.175 214.135 ;
        RECT 149.055 213.085 150.195 213.255 ;
        RECT 150.365 212.915 150.770 213.425 ;
        RECT 149.120 212.745 150.770 212.915 ;
        RECT 150.955 212.845 151.475 213.385 ;
        RECT 151.645 213.015 152.165 213.555 ;
        RECT 152.415 213.455 153.175 213.675 ;
        RECT 153.345 213.675 153.515 214.305 ;
        RECT 153.685 213.845 154.015 214.645 ;
        RECT 154.185 213.675 154.460 214.475 ;
        RECT 153.345 213.465 154.460 213.675 ;
        RECT 155.095 213.505 155.355 214.645 ;
        RECT 155.525 213.495 155.855 214.475 ;
        RECT 156.025 213.505 156.305 214.645 ;
        RECT 156.935 213.555 158.145 214.645 ;
        RECT 152.415 212.915 152.630 213.455 ;
        RECT 152.800 213.085 153.570 213.285 ;
        RECT 153.740 213.085 154.460 213.285 ;
        RECT 155.115 213.085 155.450 213.335 ;
        RECT 148.195 212.265 148.495 212.595 ;
        RECT 148.665 212.095 148.940 212.575 ;
        RECT 149.120 212.355 149.415 212.745 ;
        RECT 149.585 212.095 149.840 212.575 ;
        RECT 150.015 212.355 150.275 212.745 ;
        RECT 150.445 212.095 150.725 212.575 ;
        RECT 150.955 212.095 152.165 212.845 ;
        RECT 152.415 212.745 154.015 212.915 ;
        RECT 152.845 212.735 154.015 212.745 ;
        RECT 152.385 212.095 152.675 212.565 ;
        RECT 152.845 212.265 153.175 212.735 ;
        RECT 153.345 212.095 153.515 212.565 ;
        RECT 153.685 212.265 154.015 212.735 ;
        RECT 154.185 212.095 154.460 212.915 ;
        RECT 155.620 212.895 155.790 213.495 ;
        RECT 155.960 213.065 156.295 213.335 ;
        RECT 156.935 213.015 157.455 213.555 ;
        RECT 155.095 212.265 155.790 212.895 ;
        RECT 155.995 212.095 156.305 212.895 ;
        RECT 157.625 212.845 158.145 213.385 ;
        RECT 156.935 212.095 158.145 212.845 ;
        RECT 2.750 211.925 158.230 212.095 ;
        RECT 2.835 211.175 4.045 211.925 ;
        RECT 4.680 211.375 4.935 211.665 ;
        RECT 5.105 211.545 5.435 211.925 ;
        RECT 4.680 211.205 5.430 211.375 ;
        RECT 2.835 210.635 3.355 211.175 ;
        RECT 3.525 210.465 4.045 211.005 ;
        RECT 2.835 209.375 4.045 210.465 ;
        RECT 4.680 210.385 5.030 211.035 ;
        RECT 5.200 210.215 5.430 211.205 ;
        RECT 4.680 210.045 5.430 210.215 ;
        RECT 4.680 209.545 4.935 210.045 ;
        RECT 5.105 209.375 5.435 209.875 ;
        RECT 5.605 209.545 5.775 211.665 ;
        RECT 6.135 211.565 6.465 211.925 ;
        RECT 6.635 211.535 7.130 211.705 ;
        RECT 7.335 211.535 8.190 211.705 ;
        RECT 6.005 210.345 6.465 211.395 ;
        RECT 5.945 209.560 6.270 210.345 ;
        RECT 6.635 210.175 6.805 211.535 ;
        RECT 6.975 210.625 7.325 211.245 ;
        RECT 7.495 211.025 7.850 211.245 ;
        RECT 7.495 210.435 7.665 211.025 ;
        RECT 8.020 210.825 8.190 211.535 ;
        RECT 9.065 211.465 9.395 211.925 ;
        RECT 9.605 211.565 9.955 211.735 ;
        RECT 8.395 210.995 9.185 211.245 ;
        RECT 9.605 211.175 9.865 211.565 ;
        RECT 10.175 211.475 11.125 211.755 ;
        RECT 11.295 211.485 11.485 211.925 ;
        RECT 11.655 211.545 12.725 211.715 ;
        RECT 9.355 210.825 9.525 211.005 ;
        RECT 6.635 210.005 7.030 210.175 ;
        RECT 7.200 210.045 7.665 210.435 ;
        RECT 7.835 210.655 9.525 210.825 ;
        RECT 6.860 209.875 7.030 210.005 ;
        RECT 7.835 209.875 8.005 210.655 ;
        RECT 9.695 210.485 9.865 211.175 ;
        RECT 8.365 210.315 9.865 210.485 ;
        RECT 10.055 210.515 10.265 211.305 ;
        RECT 10.435 210.685 10.785 211.305 ;
        RECT 10.955 210.695 11.125 211.475 ;
        RECT 11.655 211.315 11.825 211.545 ;
        RECT 11.295 211.145 11.825 211.315 ;
        RECT 11.295 210.865 11.515 211.145 ;
        RECT 11.995 210.975 12.235 211.375 ;
        RECT 10.955 210.525 11.360 210.695 ;
        RECT 11.695 210.605 12.235 210.975 ;
        RECT 12.405 211.190 12.725 211.545 ;
        RECT 12.405 210.935 12.730 211.190 ;
        RECT 12.925 211.115 13.095 211.925 ;
        RECT 13.265 211.275 13.595 211.755 ;
        RECT 13.765 211.455 13.935 211.925 ;
        RECT 14.105 211.275 14.435 211.755 ;
        RECT 14.605 211.455 14.775 211.925 ;
        RECT 13.265 211.105 15.030 211.275 ;
        RECT 12.405 210.725 14.435 210.935 ;
        RECT 12.405 210.715 12.750 210.725 ;
        RECT 10.055 210.355 10.730 210.515 ;
        RECT 11.190 210.435 11.360 210.525 ;
        RECT 10.055 210.345 11.020 210.355 ;
        RECT 9.695 210.175 9.865 210.315 ;
        RECT 6.440 209.375 6.690 209.835 ;
        RECT 6.860 209.545 7.110 209.875 ;
        RECT 7.325 209.545 8.005 209.875 ;
        RECT 8.175 209.975 9.250 210.145 ;
        RECT 9.695 210.005 10.255 210.175 ;
        RECT 10.560 210.055 11.020 210.345 ;
        RECT 11.190 210.265 12.410 210.435 ;
        RECT 8.175 209.635 8.345 209.975 ;
        RECT 8.580 209.375 8.910 209.805 ;
        RECT 9.080 209.635 9.250 209.975 ;
        RECT 9.545 209.375 9.915 209.835 ;
        RECT 10.085 209.545 10.255 210.005 ;
        RECT 11.190 209.885 11.360 210.265 ;
        RECT 12.580 210.095 12.750 210.715 ;
        RECT 14.620 210.555 15.030 211.105 ;
        RECT 15.255 211.155 17.845 211.925 ;
        RECT 18.105 211.375 18.275 211.665 ;
        RECT 18.445 211.545 18.775 211.925 ;
        RECT 18.105 211.205 18.770 211.375 ;
        RECT 15.255 210.635 16.465 211.155 ;
        RECT 10.490 209.545 11.360 209.885 ;
        RECT 11.950 209.925 12.750 210.095 ;
        RECT 11.530 209.375 11.780 209.835 ;
        RECT 11.950 209.635 12.120 209.925 ;
        RECT 12.300 209.375 12.630 209.755 ;
        RECT 12.925 209.375 13.095 210.435 ;
        RECT 13.305 210.385 15.030 210.555 ;
        RECT 16.635 210.465 17.845 210.985 ;
        RECT 13.305 209.545 13.595 210.385 ;
        RECT 13.765 209.375 13.935 210.215 ;
        RECT 14.145 209.545 14.395 210.385 ;
        RECT 14.605 209.375 14.775 210.215 ;
        RECT 15.255 209.375 17.845 210.465 ;
        RECT 18.020 210.385 18.370 211.035 ;
        RECT 18.540 210.215 18.770 211.205 ;
        RECT 18.105 210.045 18.770 210.215 ;
        RECT 18.105 209.545 18.275 210.045 ;
        RECT 18.445 209.375 18.775 209.875 ;
        RECT 18.945 209.545 19.170 211.665 ;
        RECT 19.385 211.545 19.715 211.925 ;
        RECT 19.885 211.375 20.055 211.705 ;
        RECT 20.355 211.545 21.370 211.745 ;
        RECT 19.360 211.185 20.055 211.375 ;
        RECT 19.360 210.215 19.530 211.185 ;
        RECT 19.700 210.385 20.110 211.005 ;
        RECT 20.280 210.435 20.500 211.305 ;
        RECT 20.680 210.995 21.030 211.365 ;
        RECT 21.200 210.815 21.370 211.545 ;
        RECT 21.540 211.485 21.950 211.925 ;
        RECT 22.240 211.285 22.490 211.715 ;
        RECT 22.690 211.465 23.010 211.925 ;
        RECT 23.570 211.535 24.420 211.705 ;
        RECT 21.540 210.945 21.950 211.275 ;
        RECT 22.240 210.945 22.660 211.285 ;
        RECT 20.950 210.775 21.370 210.815 ;
        RECT 20.950 210.605 22.300 210.775 ;
        RECT 19.360 210.045 20.055 210.215 ;
        RECT 20.280 210.055 20.780 210.435 ;
        RECT 19.385 209.375 19.715 209.875 ;
        RECT 19.885 209.545 20.055 210.045 ;
        RECT 20.950 209.760 21.120 210.605 ;
        RECT 22.050 210.445 22.300 210.605 ;
        RECT 21.290 210.175 21.540 210.435 ;
        RECT 22.470 210.175 22.660 210.945 ;
        RECT 21.290 209.925 22.660 210.175 ;
        RECT 22.830 211.115 24.080 211.285 ;
        RECT 22.830 210.355 23.000 211.115 ;
        RECT 23.750 210.995 24.080 211.115 ;
        RECT 23.170 210.535 23.350 210.945 ;
        RECT 24.250 210.775 24.420 211.535 ;
        RECT 24.620 211.445 25.280 211.925 ;
        RECT 25.460 211.330 25.780 211.660 ;
        RECT 24.610 211.005 25.270 211.275 ;
        RECT 24.610 210.945 24.940 211.005 ;
        RECT 25.090 210.775 25.420 210.835 ;
        RECT 23.520 210.605 25.420 210.775 ;
        RECT 22.830 210.045 23.350 210.355 ;
        RECT 23.520 210.095 23.690 210.605 ;
        RECT 25.590 210.435 25.780 211.330 ;
        RECT 23.860 210.265 25.780 210.435 ;
        RECT 25.460 210.245 25.780 210.265 ;
        RECT 25.980 211.015 26.230 211.665 ;
        RECT 26.410 211.465 26.695 211.925 ;
        RECT 26.875 211.215 27.130 211.745 ;
        RECT 25.980 210.685 26.780 211.015 ;
        RECT 23.520 209.925 24.730 210.095 ;
        RECT 20.290 209.590 21.120 209.760 ;
        RECT 21.360 209.375 21.740 209.755 ;
        RECT 21.920 209.635 22.090 209.925 ;
        RECT 23.520 209.845 23.690 209.925 ;
        RECT 22.260 209.375 22.590 209.755 ;
        RECT 23.060 209.595 23.690 209.845 ;
        RECT 23.870 209.375 24.290 209.755 ;
        RECT 24.490 209.635 24.730 209.925 ;
        RECT 24.960 209.375 25.290 210.065 ;
        RECT 25.460 209.635 25.630 210.245 ;
        RECT 25.980 210.095 26.230 210.685 ;
        RECT 26.950 210.355 27.130 211.215 ;
        RECT 28.595 211.200 28.885 211.925 ;
        RECT 29.520 211.375 29.775 211.665 ;
        RECT 29.945 211.545 30.275 211.925 ;
        RECT 29.520 211.205 30.270 211.375 ;
        RECT 25.900 209.585 26.230 210.095 ;
        RECT 26.410 209.375 26.695 210.175 ;
        RECT 26.875 209.885 27.130 210.355 ;
        RECT 26.875 209.715 27.215 209.885 ;
        RECT 26.875 209.685 27.130 209.715 ;
        RECT 28.595 209.375 28.885 210.540 ;
        RECT 29.520 210.385 29.870 211.035 ;
        RECT 30.040 210.215 30.270 211.205 ;
        RECT 29.520 210.045 30.270 210.215 ;
        RECT 29.520 209.545 29.775 210.045 ;
        RECT 29.945 209.375 30.275 209.875 ;
        RECT 30.445 209.545 30.615 211.665 ;
        RECT 30.975 211.565 31.305 211.925 ;
        RECT 31.475 211.535 31.970 211.705 ;
        RECT 32.175 211.535 33.030 211.705 ;
        RECT 30.845 210.345 31.305 211.395 ;
        RECT 30.785 209.560 31.110 210.345 ;
        RECT 31.475 210.175 31.645 211.535 ;
        RECT 31.815 210.625 32.165 211.245 ;
        RECT 32.335 211.025 32.690 211.245 ;
        RECT 32.335 210.435 32.505 211.025 ;
        RECT 32.860 210.825 33.030 211.535 ;
        RECT 33.905 211.465 34.235 211.925 ;
        RECT 34.445 211.565 34.795 211.735 ;
        RECT 33.235 210.995 34.025 211.245 ;
        RECT 34.445 211.175 34.705 211.565 ;
        RECT 35.015 211.475 35.965 211.755 ;
        RECT 36.135 211.485 36.325 211.925 ;
        RECT 36.495 211.545 37.565 211.715 ;
        RECT 34.195 210.825 34.365 211.005 ;
        RECT 31.475 210.005 31.870 210.175 ;
        RECT 32.040 210.045 32.505 210.435 ;
        RECT 32.675 210.655 34.365 210.825 ;
        RECT 31.700 209.875 31.870 210.005 ;
        RECT 32.675 209.875 32.845 210.655 ;
        RECT 34.535 210.485 34.705 211.175 ;
        RECT 33.205 210.315 34.705 210.485 ;
        RECT 34.895 210.515 35.105 211.305 ;
        RECT 35.275 210.685 35.625 211.305 ;
        RECT 35.795 210.695 35.965 211.475 ;
        RECT 36.495 211.315 36.665 211.545 ;
        RECT 36.135 211.145 36.665 211.315 ;
        RECT 36.135 210.865 36.355 211.145 ;
        RECT 36.835 210.975 37.075 211.375 ;
        RECT 35.795 210.525 36.200 210.695 ;
        RECT 36.535 210.605 37.075 210.975 ;
        RECT 37.245 211.190 37.565 211.545 ;
        RECT 37.245 210.935 37.570 211.190 ;
        RECT 37.765 211.115 37.935 211.925 ;
        RECT 38.105 211.275 38.435 211.755 ;
        RECT 38.605 211.455 38.775 211.925 ;
        RECT 38.945 211.275 39.275 211.755 ;
        RECT 39.445 211.455 39.615 211.925 ;
        RECT 40.100 211.375 40.355 211.665 ;
        RECT 40.525 211.545 40.855 211.925 ;
        RECT 38.105 211.105 39.870 211.275 ;
        RECT 40.100 211.205 40.850 211.375 ;
        RECT 37.245 210.725 39.275 210.935 ;
        RECT 37.245 210.715 37.590 210.725 ;
        RECT 34.895 210.355 35.570 210.515 ;
        RECT 36.030 210.435 36.200 210.525 ;
        RECT 34.895 210.345 35.860 210.355 ;
        RECT 34.535 210.175 34.705 210.315 ;
        RECT 31.280 209.375 31.530 209.835 ;
        RECT 31.700 209.545 31.950 209.875 ;
        RECT 32.165 209.545 32.845 209.875 ;
        RECT 33.015 209.975 34.090 210.145 ;
        RECT 34.535 210.005 35.095 210.175 ;
        RECT 35.400 210.055 35.860 210.345 ;
        RECT 36.030 210.265 37.250 210.435 ;
        RECT 33.015 209.635 33.185 209.975 ;
        RECT 33.420 209.375 33.750 209.805 ;
        RECT 33.920 209.635 34.090 209.975 ;
        RECT 34.385 209.375 34.755 209.835 ;
        RECT 34.925 209.545 35.095 210.005 ;
        RECT 36.030 209.885 36.200 210.265 ;
        RECT 37.420 210.095 37.590 210.715 ;
        RECT 39.460 210.555 39.870 211.105 ;
        RECT 35.330 209.545 36.200 209.885 ;
        RECT 36.790 209.925 37.590 210.095 ;
        RECT 36.370 209.375 36.620 209.835 ;
        RECT 36.790 209.635 36.960 209.925 ;
        RECT 37.140 209.375 37.470 209.755 ;
        RECT 37.765 209.375 37.935 210.435 ;
        RECT 38.145 210.385 39.870 210.555 ;
        RECT 40.100 210.385 40.450 211.035 ;
        RECT 38.145 209.545 38.435 210.385 ;
        RECT 38.605 209.375 38.775 210.215 ;
        RECT 38.985 209.545 39.235 210.385 ;
        RECT 40.620 210.215 40.850 211.205 ;
        RECT 39.445 209.375 39.615 210.215 ;
        RECT 40.100 210.045 40.850 210.215 ;
        RECT 40.100 209.545 40.355 210.045 ;
        RECT 40.525 209.375 40.855 209.875 ;
        RECT 41.025 209.545 41.195 211.665 ;
        RECT 41.555 211.565 41.885 211.925 ;
        RECT 42.055 211.535 42.550 211.705 ;
        RECT 42.755 211.535 43.610 211.705 ;
        RECT 41.425 210.345 41.885 211.395 ;
        RECT 41.365 209.560 41.690 210.345 ;
        RECT 42.055 210.175 42.225 211.535 ;
        RECT 42.395 210.625 42.745 211.245 ;
        RECT 42.915 211.025 43.270 211.245 ;
        RECT 42.915 210.435 43.085 211.025 ;
        RECT 43.440 210.825 43.610 211.535 ;
        RECT 44.485 211.465 44.815 211.925 ;
        RECT 45.025 211.565 45.375 211.735 ;
        RECT 43.815 210.995 44.605 211.245 ;
        RECT 45.025 211.175 45.285 211.565 ;
        RECT 45.595 211.475 46.545 211.755 ;
        RECT 46.715 211.485 46.905 211.925 ;
        RECT 47.075 211.545 48.145 211.715 ;
        RECT 44.775 210.825 44.945 211.005 ;
        RECT 42.055 210.005 42.450 210.175 ;
        RECT 42.620 210.045 43.085 210.435 ;
        RECT 43.255 210.655 44.945 210.825 ;
        RECT 42.280 209.875 42.450 210.005 ;
        RECT 43.255 209.875 43.425 210.655 ;
        RECT 45.115 210.485 45.285 211.175 ;
        RECT 43.785 210.315 45.285 210.485 ;
        RECT 45.475 210.515 45.685 211.305 ;
        RECT 45.855 210.685 46.205 211.305 ;
        RECT 46.375 210.695 46.545 211.475 ;
        RECT 47.075 211.315 47.245 211.545 ;
        RECT 46.715 211.145 47.245 211.315 ;
        RECT 46.715 210.865 46.935 211.145 ;
        RECT 47.415 210.975 47.655 211.375 ;
        RECT 46.375 210.525 46.780 210.695 ;
        RECT 47.115 210.605 47.655 210.975 ;
        RECT 47.825 211.190 48.145 211.545 ;
        RECT 48.390 211.465 48.695 211.925 ;
        RECT 48.865 211.215 49.120 211.745 ;
        RECT 47.825 211.015 48.150 211.190 ;
        RECT 47.825 210.715 48.740 211.015 ;
        RECT 48.000 210.685 48.740 210.715 ;
        RECT 45.475 210.355 46.150 210.515 ;
        RECT 46.610 210.435 46.780 210.525 ;
        RECT 45.475 210.345 46.440 210.355 ;
        RECT 45.115 210.175 45.285 210.315 ;
        RECT 41.860 209.375 42.110 209.835 ;
        RECT 42.280 209.545 42.530 209.875 ;
        RECT 42.745 209.545 43.425 209.875 ;
        RECT 43.595 209.975 44.670 210.145 ;
        RECT 45.115 210.005 45.675 210.175 ;
        RECT 45.980 210.055 46.440 210.345 ;
        RECT 46.610 210.265 47.830 210.435 ;
        RECT 43.595 209.635 43.765 209.975 ;
        RECT 44.000 209.375 44.330 209.805 ;
        RECT 44.500 209.635 44.670 209.975 ;
        RECT 44.965 209.375 45.335 209.835 ;
        RECT 45.505 209.545 45.675 210.005 ;
        RECT 46.610 209.885 46.780 210.265 ;
        RECT 48.000 210.095 48.170 210.685 ;
        RECT 48.910 210.565 49.120 211.215 ;
        RECT 49.760 211.085 50.020 211.925 ;
        RECT 50.195 211.180 50.450 211.755 ;
        RECT 50.620 211.545 50.950 211.925 ;
        RECT 51.165 211.375 51.335 211.755 ;
        RECT 51.655 211.445 51.935 211.925 ;
        RECT 50.620 211.205 51.335 211.375 ;
        RECT 52.105 211.275 52.365 211.665 ;
        RECT 52.540 211.445 52.795 211.925 ;
        RECT 52.965 211.275 53.260 211.665 ;
        RECT 53.440 211.445 53.715 211.925 ;
        RECT 53.885 211.425 54.185 211.755 ;
        RECT 45.910 209.545 46.780 209.885 ;
        RECT 47.370 209.925 48.170 210.095 ;
        RECT 46.950 209.375 47.200 209.835 ;
        RECT 47.370 209.635 47.540 209.925 ;
        RECT 47.720 209.375 48.050 209.755 ;
        RECT 48.390 209.375 48.695 210.515 ;
        RECT 48.865 209.685 49.120 210.565 ;
        RECT 49.760 209.375 50.020 210.525 ;
        RECT 50.195 210.450 50.365 211.180 ;
        RECT 50.620 211.015 50.790 211.205 ;
        RECT 51.610 211.105 53.260 211.275 ;
        RECT 50.535 210.685 50.790 211.015 ;
        RECT 50.620 210.475 50.790 210.685 ;
        RECT 51.070 210.655 51.425 211.025 ;
        RECT 51.610 210.595 52.015 211.105 ;
        RECT 52.185 210.765 53.325 210.935 ;
        RECT 50.195 209.545 50.450 210.450 ;
        RECT 50.620 210.305 51.335 210.475 ;
        RECT 51.610 210.425 52.365 210.595 ;
        RECT 50.620 209.375 50.950 210.135 ;
        RECT 51.165 209.545 51.335 210.305 ;
        RECT 51.650 209.375 51.935 210.245 ;
        RECT 52.105 210.175 52.365 210.425 ;
        RECT 53.155 210.515 53.325 210.765 ;
        RECT 53.495 210.685 53.845 211.255 ;
        RECT 54.015 210.515 54.185 211.425 ;
        RECT 54.355 211.200 54.645 211.925 ;
        RECT 54.820 211.185 55.075 211.755 ;
        RECT 55.245 211.525 55.575 211.925 ;
        RECT 56.000 211.390 56.530 211.755 ;
        RECT 56.000 211.355 56.175 211.390 ;
        RECT 55.245 211.185 56.175 211.355 ;
        RECT 53.155 210.345 54.185 210.515 ;
        RECT 52.105 210.005 53.225 210.175 ;
        RECT 52.105 209.545 52.365 210.005 ;
        RECT 52.540 209.375 52.795 209.835 ;
        RECT 52.965 209.545 53.225 210.005 ;
        RECT 53.395 209.375 53.705 210.175 ;
        RECT 53.875 209.545 54.185 210.345 ;
        RECT 54.355 209.375 54.645 210.540 ;
        RECT 54.820 210.515 54.990 211.185 ;
        RECT 55.245 211.015 55.415 211.185 ;
        RECT 55.160 210.685 55.415 211.015 ;
        RECT 55.640 210.685 55.835 211.015 ;
        RECT 54.820 209.545 55.155 210.515 ;
        RECT 55.325 209.375 55.495 210.515 ;
        RECT 55.665 209.715 55.835 210.685 ;
        RECT 56.005 210.055 56.175 211.185 ;
        RECT 56.345 210.395 56.515 211.195 ;
        RECT 56.720 210.905 56.995 211.755 ;
        RECT 56.715 210.735 56.995 210.905 ;
        RECT 56.720 210.595 56.995 210.735 ;
        RECT 57.165 210.395 57.355 211.755 ;
        RECT 57.535 211.390 58.045 211.925 ;
        RECT 58.265 211.115 58.510 211.720 ;
        RECT 59.475 211.445 59.755 211.925 ;
        RECT 59.925 211.275 60.185 211.665 ;
        RECT 60.360 211.445 60.615 211.925 ;
        RECT 60.785 211.275 61.080 211.665 ;
        RECT 61.260 211.445 61.535 211.925 ;
        RECT 61.705 211.425 62.005 211.755 ;
        RECT 57.555 210.945 58.785 211.115 ;
        RECT 56.345 210.225 57.355 210.395 ;
        RECT 57.525 210.380 58.275 210.570 ;
        RECT 56.005 209.885 57.130 210.055 ;
        RECT 57.525 209.715 57.695 210.380 ;
        RECT 58.445 210.135 58.785 210.945 ;
        RECT 59.430 211.105 61.080 211.275 ;
        RECT 59.430 210.595 59.835 211.105 ;
        RECT 60.005 210.765 61.145 210.935 ;
        RECT 59.430 210.425 60.185 210.595 ;
        RECT 55.665 209.545 57.695 209.715 ;
        RECT 57.865 209.375 58.035 210.135 ;
        RECT 58.270 209.725 58.785 210.135 ;
        RECT 59.470 209.375 59.755 210.245 ;
        RECT 59.925 210.175 60.185 210.425 ;
        RECT 60.975 210.515 61.145 210.765 ;
        RECT 61.315 210.685 61.665 211.255 ;
        RECT 61.835 210.515 62.005 211.425 ;
        RECT 62.215 211.105 62.445 211.925 ;
        RECT 62.615 211.125 62.945 211.755 ;
        RECT 62.195 210.685 62.525 210.935 ;
        RECT 62.695 210.525 62.945 211.125 ;
        RECT 63.115 211.105 63.325 211.925 ;
        RECT 63.555 211.380 68.900 211.925 ;
        RECT 69.075 211.380 74.420 211.925 ;
        RECT 74.595 211.380 79.940 211.925 ;
        RECT 65.140 210.550 65.480 211.380 ;
        RECT 60.975 210.345 62.005 210.515 ;
        RECT 59.925 210.005 61.045 210.175 ;
        RECT 59.925 209.545 60.185 210.005 ;
        RECT 60.360 209.375 60.615 209.835 ;
        RECT 60.785 209.545 61.045 210.005 ;
        RECT 61.215 209.375 61.525 210.175 ;
        RECT 61.695 209.545 62.005 210.345 ;
        RECT 62.215 209.375 62.445 210.515 ;
        RECT 62.615 209.545 62.945 210.525 ;
        RECT 63.115 209.375 63.325 210.515 ;
        RECT 66.960 209.810 67.310 211.060 ;
        RECT 70.660 210.550 71.000 211.380 ;
        RECT 72.480 209.810 72.830 211.060 ;
        RECT 76.180 210.550 76.520 211.380 ;
        RECT 80.115 211.200 80.405 211.925 ;
        RECT 80.575 211.380 85.920 211.925 ;
        RECT 78.000 209.810 78.350 211.060 ;
        RECT 82.160 210.550 82.500 211.380 ;
        RECT 86.095 211.155 87.765 211.925 ;
        RECT 87.950 211.355 88.205 211.705 ;
        RECT 88.375 211.525 88.705 211.925 ;
        RECT 88.875 211.355 89.045 211.705 ;
        RECT 89.215 211.525 89.595 211.925 ;
        RECT 87.950 211.185 89.615 211.355 ;
        RECT 89.785 211.250 90.060 211.595 ;
        RECT 63.555 209.375 68.900 209.810 ;
        RECT 69.075 209.375 74.420 209.810 ;
        RECT 74.595 209.375 79.940 209.810 ;
        RECT 80.115 209.375 80.405 210.540 ;
        RECT 83.980 209.810 84.330 211.060 ;
        RECT 86.095 210.635 86.845 211.155 ;
        RECT 89.445 211.015 89.615 211.185 ;
        RECT 87.015 210.465 87.765 210.985 ;
        RECT 87.935 210.685 88.280 211.015 ;
        RECT 88.450 210.685 89.275 211.015 ;
        RECT 89.445 210.685 89.720 211.015 ;
        RECT 80.575 209.375 85.920 209.810 ;
        RECT 86.095 209.375 87.765 210.465 ;
        RECT 87.955 210.225 88.280 210.515 ;
        RECT 88.450 210.395 88.645 210.685 ;
        RECT 89.445 210.515 89.615 210.685 ;
        RECT 89.890 210.515 90.060 211.250 ;
        RECT 90.235 211.295 90.575 211.755 ;
        RECT 90.745 211.465 90.915 211.925 ;
        RECT 91.545 211.490 91.905 211.755 ;
        RECT 91.550 211.485 91.905 211.490 ;
        RECT 91.555 211.475 91.905 211.485 ;
        RECT 91.560 211.470 91.905 211.475 ;
        RECT 91.565 211.460 91.905 211.470 ;
        RECT 92.145 211.465 92.315 211.925 ;
        RECT 91.570 211.455 91.905 211.460 ;
        RECT 91.580 211.445 91.905 211.455 ;
        RECT 91.590 211.435 91.905 211.445 ;
        RECT 91.085 211.295 91.415 211.375 ;
        RECT 90.235 211.105 91.415 211.295 ;
        RECT 91.605 211.295 91.905 211.435 ;
        RECT 91.605 211.105 92.315 211.295 ;
        RECT 88.955 210.345 89.615 210.515 ;
        RECT 88.955 210.225 89.125 210.345 ;
        RECT 87.955 210.055 89.125 210.225 ;
        RECT 87.935 209.595 89.125 209.885 ;
        RECT 89.295 209.375 89.575 210.175 ;
        RECT 89.785 209.545 90.060 210.515 ;
        RECT 90.235 210.735 90.565 210.935 ;
        RECT 90.875 210.915 91.205 210.935 ;
        RECT 90.755 210.735 91.205 210.915 ;
        RECT 90.235 210.395 90.465 210.735 ;
        RECT 90.245 209.375 90.575 210.095 ;
        RECT 90.755 209.620 90.970 210.735 ;
        RECT 91.375 210.705 91.845 210.935 ;
        RECT 92.030 210.535 92.315 211.105 ;
        RECT 92.485 210.980 92.825 211.755 ;
        RECT 93.200 211.145 93.700 211.755 ;
        RECT 91.165 210.320 92.315 210.535 ;
        RECT 91.165 209.545 91.495 210.320 ;
        RECT 91.665 209.375 92.375 210.150 ;
        RECT 92.545 209.545 92.825 210.980 ;
        RECT 92.995 210.685 93.345 210.935 ;
        RECT 93.530 210.515 93.700 211.145 ;
        RECT 94.330 211.275 94.660 211.755 ;
        RECT 94.830 211.465 95.055 211.925 ;
        RECT 95.225 211.275 95.555 211.755 ;
        RECT 94.330 211.105 95.555 211.275 ;
        RECT 95.745 211.125 95.995 211.925 ;
        RECT 96.165 211.125 96.505 211.755 ;
        RECT 93.870 210.735 94.200 210.935 ;
        RECT 94.370 210.735 94.700 210.935 ;
        RECT 94.870 210.735 95.290 210.935 ;
        RECT 95.465 210.765 96.160 210.935 ;
        RECT 95.465 210.515 95.635 210.765 ;
        RECT 96.330 210.515 96.505 211.125 ;
        RECT 93.200 210.345 95.635 210.515 ;
        RECT 93.200 209.545 93.530 210.345 ;
        RECT 93.700 209.375 94.030 210.175 ;
        RECT 94.330 209.545 94.660 210.345 ;
        RECT 95.305 209.375 95.555 210.175 ;
        RECT 95.825 209.375 95.995 210.515 ;
        RECT 96.165 209.545 96.505 210.515 ;
        RECT 96.675 211.125 97.015 211.755 ;
        RECT 97.305 211.465 97.475 211.925 ;
        RECT 97.745 211.295 98.075 211.740 ;
        RECT 96.675 210.555 96.945 211.125 ;
        RECT 97.325 211.105 98.075 211.295 ;
        RECT 98.245 211.275 98.415 211.595 ;
        RECT 98.640 211.465 98.970 211.925 ;
        RECT 99.170 211.275 99.500 211.755 ;
        RECT 99.715 211.465 100.045 211.925 ;
        RECT 100.215 211.275 100.545 211.755 ;
        RECT 98.245 211.105 100.545 211.275 ;
        RECT 100.815 211.155 104.325 211.925 ;
        RECT 104.495 211.175 105.705 211.925 ;
        RECT 105.875 211.200 106.165 211.925 ;
        RECT 97.325 210.935 97.695 211.105 ;
        RECT 97.115 210.725 97.695 210.935 ;
        RECT 97.865 210.725 98.285 210.935 ;
        RECT 97.435 210.555 97.695 210.725 ;
        RECT 96.675 209.545 97.200 210.555 ;
        RECT 97.435 210.265 98.185 210.555 ;
        RECT 97.435 209.375 97.765 210.095 ;
        RECT 97.935 209.545 98.185 210.265 ;
        RECT 98.455 209.620 98.785 210.935 ;
        RECT 98.995 209.620 99.325 210.935 ;
        RECT 99.495 209.620 99.865 210.935 ;
        RECT 100.075 210.685 100.585 210.935 ;
        RECT 100.815 210.635 102.465 211.155 ;
        RECT 100.195 209.375 100.525 210.495 ;
        RECT 102.635 210.465 104.325 210.985 ;
        RECT 104.495 210.635 105.015 211.175 ;
        RECT 106.335 211.155 109.845 211.925 ;
        RECT 110.345 211.525 110.675 211.925 ;
        RECT 110.845 211.355 111.175 211.695 ;
        RECT 112.225 211.525 112.555 211.925 ;
        RECT 110.190 211.185 112.555 211.355 ;
        RECT 112.725 211.200 113.055 211.710 ;
        RECT 105.185 210.465 105.705 211.005 ;
        RECT 106.335 210.635 107.985 211.155 ;
        RECT 100.815 209.375 104.325 210.465 ;
        RECT 104.495 209.375 105.705 210.465 ;
        RECT 105.875 209.375 106.165 210.540 ;
        RECT 108.155 210.465 109.845 210.985 ;
        RECT 106.335 209.375 109.845 210.465 ;
        RECT 110.190 210.185 110.360 211.185 ;
        RECT 112.385 211.015 112.555 211.185 ;
        RECT 110.530 210.355 110.775 211.015 ;
        RECT 110.990 210.355 111.255 211.015 ;
        RECT 111.450 210.355 111.735 211.015 ;
        RECT 111.910 210.685 112.215 211.015 ;
        RECT 112.385 210.685 112.695 211.015 ;
        RECT 111.910 210.355 112.125 210.685 ;
        RECT 112.865 210.565 113.055 211.200 ;
        RECT 113.320 211.355 113.495 211.755 ;
        RECT 113.665 211.545 113.995 211.925 ;
        RECT 114.240 211.425 114.470 211.755 ;
        RECT 113.320 211.185 113.950 211.355 ;
        RECT 113.780 211.015 113.950 211.185 ;
        RECT 110.190 210.015 110.645 210.185 ;
        RECT 110.315 209.585 110.645 210.015 ;
        RECT 110.825 210.015 112.115 210.185 ;
        RECT 110.825 209.595 111.075 210.015 ;
        RECT 111.305 209.375 111.635 209.845 ;
        RECT 111.865 209.595 112.115 210.015 ;
        RECT 112.305 209.375 112.555 210.515 ;
        RECT 112.835 210.435 113.055 210.565 ;
        RECT 112.725 209.585 113.055 210.435 ;
        RECT 113.235 210.335 113.600 211.015 ;
        RECT 113.780 210.685 114.130 211.015 ;
        RECT 113.780 210.165 113.950 210.685 ;
        RECT 113.320 209.995 113.950 210.165 ;
        RECT 114.300 210.135 114.470 211.425 ;
        RECT 114.670 210.315 114.950 211.590 ;
        RECT 115.175 211.245 115.445 211.590 ;
        RECT 115.905 211.545 116.235 211.925 ;
        RECT 116.405 211.670 116.740 211.715 ;
        RECT 115.135 211.075 115.445 211.245 ;
        RECT 115.175 210.315 115.445 211.075 ;
        RECT 115.635 210.315 115.975 211.345 ;
        RECT 116.405 211.205 116.745 211.670 ;
        RECT 116.915 211.425 117.255 211.925 ;
        RECT 116.145 210.685 116.405 211.015 ;
        RECT 116.145 210.135 116.315 210.685 ;
        RECT 116.575 210.515 116.745 211.205 ;
        RECT 116.915 210.685 117.255 211.255 ;
        RECT 117.425 211.015 117.670 211.705 ;
        RECT 117.865 211.425 118.195 211.925 ;
        RECT 118.395 211.355 118.565 211.705 ;
        RECT 118.740 211.525 119.070 211.925 ;
        RECT 119.240 211.355 119.410 211.705 ;
        RECT 119.580 211.525 119.960 211.925 ;
        RECT 118.395 211.185 119.980 211.355 ;
        RECT 120.150 211.250 120.425 211.595 ;
        RECT 119.810 211.015 119.980 211.185 ;
        RECT 117.425 210.685 118.080 211.015 ;
        RECT 113.320 209.545 113.495 209.995 ;
        RECT 114.300 209.965 116.315 210.135 ;
        RECT 113.665 209.375 113.995 209.815 ;
        RECT 114.300 209.545 114.470 209.965 ;
        RECT 114.705 209.375 115.375 209.785 ;
        RECT 115.590 209.545 115.760 209.965 ;
        RECT 115.960 209.375 116.290 209.785 ;
        RECT 116.485 209.545 116.745 210.515 ;
        RECT 116.915 209.375 117.255 210.450 ;
        RECT 117.425 210.090 117.665 210.685 ;
        RECT 117.860 210.225 118.180 210.515 ;
        RECT 118.350 210.395 119.090 211.015 ;
        RECT 119.260 210.685 119.640 211.015 ;
        RECT 119.810 210.685 120.085 211.015 ;
        RECT 119.810 210.515 119.980 210.685 ;
        RECT 120.255 210.515 120.425 211.250 ;
        RECT 119.320 210.345 119.980 210.515 ;
        RECT 119.320 210.225 119.490 210.345 ;
        RECT 117.860 210.055 119.490 210.225 ;
        RECT 117.440 209.595 119.490 209.885 ;
        RECT 119.660 209.375 119.940 210.175 ;
        RECT 120.150 209.545 120.425 210.515 ;
        RECT 120.605 209.555 120.865 211.745 ;
        RECT 121.125 211.555 121.795 211.925 ;
        RECT 121.975 211.375 122.285 211.745 ;
        RECT 121.055 211.175 122.285 211.375 ;
        RECT 121.055 210.505 121.345 211.175 ;
        RECT 122.465 210.995 122.695 211.635 ;
        RECT 122.875 211.195 123.165 211.925 ;
        RECT 123.815 211.125 124.510 211.755 ;
        RECT 124.715 211.125 125.025 211.925 ;
        RECT 125.245 211.455 125.535 211.925 ;
        RECT 125.705 211.285 126.035 211.755 ;
        RECT 126.205 211.455 126.375 211.925 ;
        RECT 126.545 211.285 126.875 211.755 ;
        RECT 125.705 211.275 126.875 211.285 ;
        RECT 121.525 210.685 121.990 210.995 ;
        RECT 122.170 210.685 122.695 210.995 ;
        RECT 122.875 210.685 123.175 211.015 ;
        RECT 123.835 210.685 124.170 210.935 ;
        RECT 124.340 210.565 124.510 211.125 ;
        RECT 125.275 211.105 126.875 211.275 ;
        RECT 127.045 211.105 127.320 211.925 ;
        RECT 127.495 211.155 131.005 211.925 ;
        RECT 131.635 211.200 131.925 211.925 ;
        RECT 132.095 211.185 132.680 211.755 ;
        RECT 132.930 211.355 133.260 211.700 ;
        RECT 133.475 211.525 133.850 211.925 ;
        RECT 134.030 211.355 134.325 211.700 ;
        RECT 132.930 211.185 134.325 211.355 ;
        RECT 134.495 211.185 135.165 211.925 ;
        RECT 124.680 210.685 125.015 210.955 ;
        RECT 124.335 210.525 124.510 210.565 ;
        RECT 125.275 210.565 125.490 211.105 ;
        RECT 125.660 210.735 126.430 210.935 ;
        RECT 126.600 210.735 127.320 210.935 ;
        RECT 127.495 210.635 129.145 211.155 ;
        RECT 121.055 210.285 121.825 210.505 ;
        RECT 121.035 209.375 121.375 210.105 ;
        RECT 121.555 209.555 121.825 210.285 ;
        RECT 122.005 210.265 123.165 210.505 ;
        RECT 122.005 209.555 122.235 210.265 ;
        RECT 122.405 209.375 122.735 210.085 ;
        RECT 122.905 209.555 123.165 210.265 ;
        RECT 123.815 209.375 124.075 210.515 ;
        RECT 124.245 209.545 124.575 210.525 ;
        RECT 124.745 209.375 125.025 210.515 ;
        RECT 125.275 210.345 126.035 210.565 ;
        RECT 125.235 209.715 125.535 210.175 ;
        RECT 125.705 209.885 126.035 210.345 ;
        RECT 126.205 210.345 127.320 210.555 ;
        RECT 129.315 210.465 131.005 210.985 ;
        RECT 132.095 210.685 132.340 211.015 ;
        RECT 126.205 209.715 126.375 210.345 ;
        RECT 125.235 209.545 126.375 209.715 ;
        RECT 126.545 209.375 126.875 210.175 ;
        RECT 127.045 209.545 127.320 210.345 ;
        RECT 127.495 209.375 131.005 210.465 ;
        RECT 131.635 209.375 131.925 210.540 ;
        RECT 132.510 210.515 132.680 211.185 ;
        RECT 132.850 210.685 133.250 211.015 ;
        RECT 133.420 210.685 133.710 211.015 ;
        RECT 132.095 210.345 133.305 210.515 ;
        RECT 132.095 209.545 132.385 210.345 ;
        RECT 132.555 209.375 132.790 210.175 ;
        RECT 132.975 209.715 133.305 210.345 ;
        RECT 133.475 209.940 133.710 210.685 ;
        RECT 133.900 210.685 134.240 211.015 ;
        RECT 134.410 210.685 134.745 211.015 ;
        RECT 133.900 209.940 134.170 210.685 ;
        RECT 134.915 210.515 135.085 211.015 ;
        RECT 135.335 210.940 135.605 211.755 ;
        RECT 134.340 210.345 135.085 210.515 ;
        RECT 134.340 209.715 134.510 210.345 ;
        RECT 132.975 209.545 134.510 209.715 ;
        RECT 134.680 209.375 135.085 210.175 ;
        RECT 135.255 209.545 135.605 210.940 ;
        RECT 135.775 211.155 138.365 211.925 ;
        RECT 138.535 211.185 138.975 211.745 ;
        RECT 139.145 211.185 139.595 211.925 ;
        RECT 139.765 211.355 139.935 211.755 ;
        RECT 140.105 211.525 140.525 211.925 ;
        RECT 140.695 211.355 140.925 211.755 ;
        RECT 139.765 211.185 140.925 211.355 ;
        RECT 141.095 211.185 141.585 211.755 ;
        RECT 141.755 211.380 147.100 211.925 ;
        RECT 135.775 210.635 136.985 211.155 ;
        RECT 137.155 210.465 138.365 210.985 ;
        RECT 135.775 209.375 138.365 210.465 ;
        RECT 138.535 210.175 138.845 211.185 ;
        RECT 139.015 210.565 139.185 211.015 ;
        RECT 139.355 210.735 139.745 211.015 ;
        RECT 139.930 210.685 140.175 211.015 ;
        RECT 139.015 210.395 139.805 210.565 ;
        RECT 138.535 209.545 138.975 210.175 ;
        RECT 139.150 209.375 139.465 210.225 ;
        RECT 139.635 209.715 139.805 210.395 ;
        RECT 139.975 209.885 140.175 210.685 ;
        RECT 140.375 209.885 140.625 211.015 ;
        RECT 140.840 210.685 141.245 211.015 ;
        RECT 141.415 210.515 141.585 211.185 ;
        RECT 143.340 210.550 143.680 211.380 ;
        RECT 147.275 211.155 150.785 211.925 ;
        RECT 151.415 211.295 151.755 211.755 ;
        RECT 151.925 211.465 152.095 211.925 ;
        RECT 152.265 211.545 153.435 211.755 ;
        RECT 152.265 211.295 152.515 211.545 ;
        RECT 153.105 211.525 153.435 211.545 ;
        RECT 140.815 210.345 141.585 210.515 ;
        RECT 140.815 209.715 141.065 210.345 ;
        RECT 139.635 209.545 141.065 209.715 ;
        RECT 141.245 209.375 141.575 210.175 ;
        RECT 145.160 209.810 145.510 211.060 ;
        RECT 147.275 210.635 148.925 211.155 ;
        RECT 151.415 211.125 152.515 211.295 ;
        RECT 152.685 211.105 153.545 211.355 ;
        RECT 149.095 210.465 150.785 210.985 ;
        RECT 151.415 210.685 152.175 210.935 ;
        RECT 152.345 210.685 153.095 210.935 ;
        RECT 153.265 210.515 153.545 211.105 ;
        RECT 153.715 211.155 156.305 211.925 ;
        RECT 156.935 211.175 158.145 211.925 ;
        RECT 153.715 210.635 154.925 211.155 ;
        RECT 141.755 209.375 147.100 209.810 ;
        RECT 147.275 209.375 150.785 210.465 ;
        RECT 151.415 209.375 151.675 210.515 ;
        RECT 151.845 210.345 153.545 210.515 ;
        RECT 155.095 210.465 156.305 210.985 ;
        RECT 151.845 209.545 152.175 210.345 ;
        RECT 152.345 209.375 152.515 210.175 ;
        RECT 152.685 209.545 153.015 210.345 ;
        RECT 153.185 209.375 153.440 210.175 ;
        RECT 153.715 209.375 156.305 210.465 ;
        RECT 156.935 210.465 157.455 211.005 ;
        RECT 157.625 210.635 158.145 211.175 ;
        RECT 156.935 209.375 158.145 210.465 ;
        RECT 2.750 209.205 158.230 209.375 ;
        RECT 2.835 208.115 4.045 209.205 ;
        RECT 4.220 208.535 4.475 209.035 ;
        RECT 4.645 208.705 4.975 209.205 ;
        RECT 4.220 208.365 4.970 208.535 ;
        RECT 2.835 207.405 3.355 207.945 ;
        RECT 3.525 207.575 4.045 208.115 ;
        RECT 4.220 207.545 4.570 208.195 ;
        RECT 2.835 206.655 4.045 207.405 ;
        RECT 4.740 207.375 4.970 208.365 ;
        RECT 4.220 207.205 4.970 207.375 ;
        RECT 4.220 206.915 4.475 207.205 ;
        RECT 4.645 206.655 4.975 207.035 ;
        RECT 5.145 206.915 5.315 209.035 ;
        RECT 5.485 208.235 5.810 209.020 ;
        RECT 5.980 208.745 6.230 209.205 ;
        RECT 6.400 208.705 6.650 209.035 ;
        RECT 6.865 208.705 7.545 209.035 ;
        RECT 6.400 208.575 6.570 208.705 ;
        RECT 6.175 208.405 6.570 208.575 ;
        RECT 5.545 207.185 6.005 208.235 ;
        RECT 6.175 207.045 6.345 208.405 ;
        RECT 6.740 208.145 7.205 208.535 ;
        RECT 6.515 207.335 6.865 207.955 ;
        RECT 7.035 207.555 7.205 208.145 ;
        RECT 7.375 207.925 7.545 208.705 ;
        RECT 7.715 208.605 7.885 208.945 ;
        RECT 8.120 208.775 8.450 209.205 ;
        RECT 8.620 208.605 8.790 208.945 ;
        RECT 9.085 208.745 9.455 209.205 ;
        RECT 7.715 208.435 8.790 208.605 ;
        RECT 9.625 208.575 9.795 209.035 ;
        RECT 10.030 208.695 10.900 209.035 ;
        RECT 11.070 208.745 11.320 209.205 ;
        RECT 9.235 208.405 9.795 208.575 ;
        RECT 9.235 208.265 9.405 208.405 ;
        RECT 7.905 208.095 9.405 208.265 ;
        RECT 10.100 208.235 10.560 208.525 ;
        RECT 7.375 207.755 9.065 207.925 ;
        RECT 7.035 207.335 7.390 207.555 ;
        RECT 7.560 207.045 7.730 207.755 ;
        RECT 7.935 207.335 8.725 207.585 ;
        RECT 8.895 207.575 9.065 207.755 ;
        RECT 9.235 207.405 9.405 208.095 ;
        RECT 5.675 206.655 6.005 207.015 ;
        RECT 6.175 206.875 6.670 207.045 ;
        RECT 6.875 206.875 7.730 207.045 ;
        RECT 8.605 206.655 8.935 207.115 ;
        RECT 9.145 207.015 9.405 207.405 ;
        RECT 9.595 208.225 10.560 208.235 ;
        RECT 10.730 208.315 10.900 208.695 ;
        RECT 11.490 208.655 11.660 208.945 ;
        RECT 11.840 208.825 12.170 209.205 ;
        RECT 11.490 208.485 12.290 208.655 ;
        RECT 9.595 208.065 10.270 208.225 ;
        RECT 10.730 208.145 11.950 208.315 ;
        RECT 9.595 207.275 9.805 208.065 ;
        RECT 10.730 208.055 10.900 208.145 ;
        RECT 9.975 207.275 10.325 207.895 ;
        RECT 10.495 207.885 10.900 208.055 ;
        RECT 10.495 207.105 10.665 207.885 ;
        RECT 10.835 207.435 11.055 207.715 ;
        RECT 11.235 207.605 11.775 207.975 ;
        RECT 12.120 207.895 12.290 208.485 ;
        RECT 12.510 208.065 12.815 209.205 ;
        RECT 12.985 208.015 13.240 208.895 ;
        RECT 14.425 208.275 14.595 209.035 ;
        RECT 14.775 208.445 15.105 209.205 ;
        RECT 14.425 208.105 15.090 208.275 ;
        RECT 15.275 208.130 15.545 209.035 ;
        RECT 12.120 207.865 12.860 207.895 ;
        RECT 10.835 207.265 11.365 207.435 ;
        RECT 9.145 206.845 9.495 207.015 ;
        RECT 9.715 206.825 10.665 207.105 ;
        RECT 10.835 206.655 11.025 207.095 ;
        RECT 11.195 207.035 11.365 207.265 ;
        RECT 11.535 207.205 11.775 207.605 ;
        RECT 11.945 207.565 12.860 207.865 ;
        RECT 11.945 207.390 12.270 207.565 ;
        RECT 11.945 207.035 12.265 207.390 ;
        RECT 13.030 207.365 13.240 208.015 ;
        RECT 14.920 207.960 15.090 208.105 ;
        RECT 14.355 207.555 14.685 207.925 ;
        RECT 14.920 207.630 15.205 207.960 ;
        RECT 14.920 207.375 15.090 207.630 ;
        RECT 11.195 206.865 12.265 207.035 ;
        RECT 12.510 206.655 12.815 207.115 ;
        RECT 12.985 206.835 13.240 207.365 ;
        RECT 14.425 207.205 15.090 207.375 ;
        RECT 15.375 207.330 15.545 208.130 ;
        RECT 15.715 208.040 16.005 209.205 ;
        RECT 16.175 208.650 16.780 209.205 ;
        RECT 16.955 208.695 17.435 209.035 ;
        RECT 17.605 208.660 17.860 209.205 ;
        RECT 16.175 208.550 16.790 208.650 ;
        RECT 16.605 208.525 16.790 208.550 ;
        RECT 16.175 207.930 16.435 208.380 ;
        RECT 16.605 208.280 16.935 208.525 ;
        RECT 17.105 208.205 17.860 208.455 ;
        RECT 18.030 208.335 18.305 209.035 ;
        RECT 17.090 208.170 17.860 208.205 ;
        RECT 17.075 208.160 17.860 208.170 ;
        RECT 17.070 208.145 17.965 208.160 ;
        RECT 17.050 208.130 17.965 208.145 ;
        RECT 17.030 208.120 17.965 208.130 ;
        RECT 17.005 208.110 17.965 208.120 ;
        RECT 16.935 208.080 17.965 208.110 ;
        RECT 16.915 208.050 17.965 208.080 ;
        RECT 16.895 208.020 17.965 208.050 ;
        RECT 16.865 207.995 17.965 208.020 ;
        RECT 16.830 207.960 17.965 207.995 ;
        RECT 16.800 207.955 17.965 207.960 ;
        RECT 16.800 207.950 17.190 207.955 ;
        RECT 16.800 207.940 17.165 207.950 ;
        RECT 16.800 207.935 17.150 207.940 ;
        RECT 16.800 207.930 17.135 207.935 ;
        RECT 16.175 207.925 17.135 207.930 ;
        RECT 16.175 207.915 17.125 207.925 ;
        RECT 16.175 207.910 17.115 207.915 ;
        RECT 16.175 207.900 17.105 207.910 ;
        RECT 16.175 207.890 17.100 207.900 ;
        RECT 16.175 207.885 17.095 207.890 ;
        RECT 16.175 207.870 17.085 207.885 ;
        RECT 16.175 207.855 17.080 207.870 ;
        RECT 16.175 207.830 17.070 207.855 ;
        RECT 16.175 207.760 17.065 207.830 ;
        RECT 14.425 206.825 14.595 207.205 ;
        RECT 14.775 206.655 15.105 207.035 ;
        RECT 15.285 206.825 15.545 207.330 ;
        RECT 15.715 206.655 16.005 207.380 ;
        RECT 16.175 207.205 16.725 207.590 ;
        RECT 16.895 207.035 17.065 207.760 ;
        RECT 16.175 206.865 17.065 207.035 ;
        RECT 17.235 207.360 17.565 207.785 ;
        RECT 17.735 207.560 17.965 207.955 ;
        RECT 17.235 206.875 17.455 207.360 ;
        RECT 18.135 207.305 18.305 208.335 ;
        RECT 17.625 206.655 17.875 207.195 ;
        RECT 18.045 206.825 18.305 207.305 ;
        RECT 18.480 208.065 18.815 209.035 ;
        RECT 18.985 208.065 19.155 209.205 ;
        RECT 19.325 208.865 21.355 209.035 ;
        RECT 18.480 207.395 18.650 208.065 ;
        RECT 19.325 207.895 19.495 208.865 ;
        RECT 18.820 207.565 19.075 207.895 ;
        RECT 19.300 207.565 19.495 207.895 ;
        RECT 19.665 208.525 20.790 208.695 ;
        RECT 18.905 207.395 19.075 207.565 ;
        RECT 19.665 207.395 19.835 208.525 ;
        RECT 18.480 206.825 18.735 207.395 ;
        RECT 18.905 207.225 19.835 207.395 ;
        RECT 20.005 208.185 21.015 208.355 ;
        RECT 20.005 207.385 20.175 208.185 ;
        RECT 19.660 207.190 19.835 207.225 ;
        RECT 18.905 206.655 19.235 207.055 ;
        RECT 19.660 206.825 20.190 207.190 ;
        RECT 20.380 207.165 20.655 207.985 ;
        RECT 20.375 206.995 20.655 207.165 ;
        RECT 20.380 206.825 20.655 206.995 ;
        RECT 20.825 206.825 21.015 208.185 ;
        RECT 21.185 208.200 21.355 208.865 ;
        RECT 21.525 208.445 21.695 209.205 ;
        RECT 21.930 208.445 22.445 208.855 ;
        RECT 21.185 208.010 21.935 208.200 ;
        RECT 22.105 207.635 22.445 208.445 ;
        RECT 21.215 207.465 22.445 207.635 ;
        RECT 22.615 208.445 23.130 208.855 ;
        RECT 23.365 208.445 23.535 209.205 ;
        RECT 23.705 208.865 25.735 209.035 ;
        RECT 22.615 207.635 22.955 208.445 ;
        RECT 23.705 208.200 23.875 208.865 ;
        RECT 24.270 208.525 25.395 208.695 ;
        RECT 23.125 208.010 23.875 208.200 ;
        RECT 24.045 208.185 25.055 208.355 ;
        RECT 22.615 207.465 23.845 207.635 ;
        RECT 21.195 206.655 21.705 207.190 ;
        RECT 21.925 206.860 22.170 207.465 ;
        RECT 22.890 206.860 23.135 207.465 ;
        RECT 23.355 206.655 23.865 207.190 ;
        RECT 24.045 206.825 24.235 208.185 ;
        RECT 24.405 207.165 24.680 207.985 ;
        RECT 24.885 207.385 25.055 208.185 ;
        RECT 25.225 207.395 25.395 208.525 ;
        RECT 25.565 207.895 25.735 208.865 ;
        RECT 25.905 208.065 26.075 209.205 ;
        RECT 26.245 208.065 26.580 209.035 ;
        RECT 25.565 207.565 25.760 207.895 ;
        RECT 25.985 207.565 26.240 207.895 ;
        RECT 25.985 207.395 26.155 207.565 ;
        RECT 26.410 207.395 26.580 208.065 ;
        RECT 26.755 208.445 27.270 208.855 ;
        RECT 27.505 208.445 27.675 209.205 ;
        RECT 27.845 208.865 29.875 209.035 ;
        RECT 26.755 207.635 27.095 208.445 ;
        RECT 27.845 208.200 28.015 208.865 ;
        RECT 28.410 208.525 29.535 208.695 ;
        RECT 27.265 208.010 28.015 208.200 ;
        RECT 28.185 208.185 29.195 208.355 ;
        RECT 26.755 207.465 27.985 207.635 ;
        RECT 25.225 207.225 26.155 207.395 ;
        RECT 25.225 207.190 25.400 207.225 ;
        RECT 24.405 206.995 24.685 207.165 ;
        RECT 24.405 206.825 24.680 206.995 ;
        RECT 24.870 206.825 25.400 207.190 ;
        RECT 25.825 206.655 26.155 207.055 ;
        RECT 26.325 206.825 26.580 207.395 ;
        RECT 27.030 206.860 27.275 207.465 ;
        RECT 27.495 206.655 28.005 207.190 ;
        RECT 28.185 206.825 28.375 208.185 ;
        RECT 28.545 207.165 28.820 207.985 ;
        RECT 29.025 207.385 29.195 208.185 ;
        RECT 29.365 207.395 29.535 208.525 ;
        RECT 29.705 207.895 29.875 208.865 ;
        RECT 30.045 208.065 30.215 209.205 ;
        RECT 30.385 208.065 30.720 209.035 ;
        RECT 29.705 207.565 29.900 207.895 ;
        RECT 30.125 207.565 30.380 207.895 ;
        RECT 30.125 207.395 30.295 207.565 ;
        RECT 30.550 207.395 30.720 208.065 ;
        RECT 29.365 207.225 30.295 207.395 ;
        RECT 29.365 207.190 29.540 207.225 ;
        RECT 28.545 206.995 28.825 207.165 ;
        RECT 28.545 206.825 28.820 206.995 ;
        RECT 29.010 206.825 29.540 207.190 ;
        RECT 29.965 206.655 30.295 207.055 ;
        RECT 30.465 206.825 30.720 207.395 ;
        RECT 31.360 208.065 31.695 209.035 ;
        RECT 31.865 208.065 32.035 209.205 ;
        RECT 32.205 208.865 34.235 209.035 ;
        RECT 31.360 207.395 31.530 208.065 ;
        RECT 32.205 207.895 32.375 208.865 ;
        RECT 31.700 207.565 31.955 207.895 ;
        RECT 32.180 207.565 32.375 207.895 ;
        RECT 32.545 208.525 33.670 208.695 ;
        RECT 31.785 207.395 31.955 207.565 ;
        RECT 32.545 207.395 32.715 208.525 ;
        RECT 31.360 206.825 31.615 207.395 ;
        RECT 31.785 207.225 32.715 207.395 ;
        RECT 32.885 208.185 33.895 208.355 ;
        RECT 32.885 207.385 33.055 208.185 ;
        RECT 33.260 207.505 33.535 207.985 ;
        RECT 33.255 207.335 33.535 207.505 ;
        RECT 32.540 207.190 32.715 207.225 ;
        RECT 31.785 206.655 32.115 207.055 ;
        RECT 32.540 206.825 33.070 207.190 ;
        RECT 33.260 206.825 33.535 207.335 ;
        RECT 33.705 206.825 33.895 208.185 ;
        RECT 34.065 208.200 34.235 208.865 ;
        RECT 34.405 208.445 34.575 209.205 ;
        RECT 34.810 208.445 35.325 208.855 ;
        RECT 34.065 208.010 34.815 208.200 ;
        RECT 34.985 207.635 35.325 208.445 ;
        RECT 36.010 208.335 36.295 209.205 ;
        RECT 36.465 208.575 36.725 209.035 ;
        RECT 36.900 208.745 37.155 209.205 ;
        RECT 37.325 208.575 37.585 209.035 ;
        RECT 36.465 208.405 37.585 208.575 ;
        RECT 37.755 208.405 38.065 209.205 ;
        RECT 36.465 208.155 36.725 208.405 ;
        RECT 38.235 208.235 38.545 209.035 ;
        RECT 38.770 208.335 39.055 209.205 ;
        RECT 39.225 208.575 39.485 209.035 ;
        RECT 39.660 208.745 39.915 209.205 ;
        RECT 40.085 208.575 40.345 209.035 ;
        RECT 39.225 208.405 40.345 208.575 ;
        RECT 40.515 208.405 40.825 209.205 ;
        RECT 34.095 207.465 35.325 207.635 ;
        RECT 35.970 207.985 36.725 208.155 ;
        RECT 37.515 208.065 38.545 208.235 ;
        RECT 39.225 208.155 39.485 208.405 ;
        RECT 39.695 208.355 39.865 208.405 ;
        RECT 40.995 208.235 41.305 209.035 ;
        RECT 35.970 207.475 36.375 207.985 ;
        RECT 37.515 207.815 37.685 208.065 ;
        RECT 36.545 207.645 37.685 207.815 ;
        RECT 34.075 206.655 34.585 207.190 ;
        RECT 34.805 206.860 35.050 207.465 ;
        RECT 35.970 207.305 37.620 207.475 ;
        RECT 37.855 207.325 38.205 207.895 ;
        RECT 36.015 206.655 36.295 207.135 ;
        RECT 36.465 206.915 36.725 207.305 ;
        RECT 36.900 206.655 37.155 207.135 ;
        RECT 37.325 206.915 37.620 207.305 ;
        RECT 38.375 207.155 38.545 208.065 ;
        RECT 38.730 207.985 39.485 208.155 ;
        RECT 40.275 208.065 41.305 208.235 ;
        RECT 38.730 207.475 39.135 207.985 ;
        RECT 40.275 207.815 40.445 208.065 ;
        RECT 39.305 207.645 40.445 207.815 ;
        RECT 38.730 207.305 40.380 207.475 ;
        RECT 40.615 207.325 40.965 207.895 ;
        RECT 37.800 206.655 38.075 207.135 ;
        RECT 38.245 206.825 38.545 207.155 ;
        RECT 38.775 206.655 39.055 207.135 ;
        RECT 39.225 206.915 39.485 207.305 ;
        RECT 39.660 206.655 39.915 207.135 ;
        RECT 40.085 206.915 40.380 207.305 ;
        RECT 41.135 207.155 41.305 208.065 ;
        RECT 41.475 208.040 41.765 209.205 ;
        RECT 41.935 208.445 42.450 208.855 ;
        RECT 42.685 208.445 42.855 209.205 ;
        RECT 43.025 208.865 45.055 209.035 ;
        RECT 41.935 207.635 42.275 208.445 ;
        RECT 43.025 208.200 43.195 208.865 ;
        RECT 43.590 208.525 44.715 208.695 ;
        RECT 42.445 208.010 43.195 208.200 ;
        RECT 43.365 208.185 44.375 208.355 ;
        RECT 41.935 207.465 43.165 207.635 ;
        RECT 40.560 206.655 40.835 207.135 ;
        RECT 41.005 206.825 41.305 207.155 ;
        RECT 41.475 206.655 41.765 207.380 ;
        RECT 42.210 206.860 42.455 207.465 ;
        RECT 42.675 206.655 43.185 207.190 ;
        RECT 43.365 206.825 43.555 208.185 ;
        RECT 43.725 207.845 44.000 207.985 ;
        RECT 43.725 207.675 44.005 207.845 ;
        RECT 43.725 206.825 44.000 207.675 ;
        RECT 44.205 207.385 44.375 208.185 ;
        RECT 44.545 207.395 44.715 208.525 ;
        RECT 44.885 207.895 45.055 208.865 ;
        RECT 45.225 208.065 45.395 209.205 ;
        RECT 45.565 208.065 45.900 209.035 ;
        RECT 44.885 207.565 45.080 207.895 ;
        RECT 45.305 207.565 45.560 207.895 ;
        RECT 45.305 207.395 45.475 207.565 ;
        RECT 45.730 207.395 45.900 208.065 ;
        RECT 44.545 207.225 45.475 207.395 ;
        RECT 44.545 207.190 44.720 207.225 ;
        RECT 44.190 206.825 44.720 207.190 ;
        RECT 45.145 206.655 45.475 207.055 ;
        RECT 45.645 206.825 45.900 207.395 ;
        RECT 46.075 208.235 46.385 209.035 ;
        RECT 46.555 208.405 46.865 209.205 ;
        RECT 47.035 208.575 47.295 209.035 ;
        RECT 47.465 208.745 47.720 209.205 ;
        RECT 47.895 208.575 48.155 209.035 ;
        RECT 47.035 208.405 48.155 208.575 ;
        RECT 46.075 208.065 47.105 208.235 ;
        RECT 46.075 207.155 46.245 208.065 ;
        RECT 46.415 207.325 46.765 207.895 ;
        RECT 46.935 207.815 47.105 208.065 ;
        RECT 47.895 208.155 48.155 208.405 ;
        RECT 48.325 208.335 48.610 209.205 ;
        RECT 48.835 208.235 49.145 209.035 ;
        RECT 49.315 208.405 49.625 209.205 ;
        RECT 49.795 208.575 50.055 209.035 ;
        RECT 50.225 208.745 50.480 209.205 ;
        RECT 50.655 208.575 50.915 209.035 ;
        RECT 49.795 208.405 50.915 208.575 ;
        RECT 47.895 207.985 48.650 208.155 ;
        RECT 46.935 207.645 48.075 207.815 ;
        RECT 48.245 207.475 48.650 207.985 ;
        RECT 47.000 207.305 48.650 207.475 ;
        RECT 48.835 208.065 49.865 208.235 ;
        RECT 46.075 206.825 46.375 207.155 ;
        RECT 46.545 206.655 46.820 207.135 ;
        RECT 47.000 206.915 47.295 207.305 ;
        RECT 47.465 206.655 47.720 207.135 ;
        RECT 47.895 206.915 48.155 207.305 ;
        RECT 48.835 207.155 49.005 208.065 ;
        RECT 49.175 207.325 49.525 207.895 ;
        RECT 49.695 207.815 49.865 208.065 ;
        RECT 50.655 208.155 50.915 208.405 ;
        RECT 51.085 208.335 51.370 209.205 ;
        RECT 52.110 208.335 52.395 209.205 ;
        RECT 52.565 208.575 52.825 209.035 ;
        RECT 53.000 208.745 53.255 209.205 ;
        RECT 53.425 208.575 53.685 209.035 ;
        RECT 52.565 208.405 53.685 208.575 ;
        RECT 53.855 208.405 54.165 209.205 ;
        RECT 52.565 208.155 52.825 208.405 ;
        RECT 54.335 208.235 54.645 209.035 ;
        RECT 50.655 207.985 51.410 208.155 ;
        RECT 49.695 207.645 50.835 207.815 ;
        RECT 51.005 207.475 51.410 207.985 ;
        RECT 49.760 207.305 51.410 207.475 ;
        RECT 52.070 207.985 52.825 208.155 ;
        RECT 53.615 208.065 54.645 208.235 ;
        RECT 54.815 208.115 56.025 209.205 ;
        RECT 52.070 207.475 52.475 207.985 ;
        RECT 53.615 207.815 53.785 208.065 ;
        RECT 52.645 207.645 53.785 207.815 ;
        RECT 52.070 207.305 53.720 207.475 ;
        RECT 53.955 207.325 54.305 207.895 ;
        RECT 48.325 206.655 48.605 207.135 ;
        RECT 48.835 206.825 49.135 207.155 ;
        RECT 49.305 206.655 49.580 207.135 ;
        RECT 49.760 206.915 50.055 207.305 ;
        RECT 50.225 206.655 50.480 207.135 ;
        RECT 50.655 206.915 50.915 207.305 ;
        RECT 51.085 206.655 51.365 207.135 ;
        RECT 52.115 206.655 52.395 207.135 ;
        RECT 52.565 206.915 52.825 207.305 ;
        RECT 53.000 206.655 53.255 207.135 ;
        RECT 53.425 206.915 53.720 207.305 ;
        RECT 54.475 207.155 54.645 208.065 ;
        RECT 53.900 206.655 54.175 207.135 ;
        RECT 54.345 206.825 54.645 207.155 ;
        RECT 54.815 207.405 55.335 207.945 ;
        RECT 55.505 207.575 56.025 208.115 ;
        RECT 56.200 208.485 56.535 208.995 ;
        RECT 54.815 206.655 56.025 207.405 ;
        RECT 56.200 207.130 56.455 208.485 ;
        RECT 56.785 208.405 57.115 209.205 ;
        RECT 57.360 208.615 57.645 209.035 ;
        RECT 57.900 208.785 58.230 209.205 ;
        RECT 58.455 208.865 59.615 209.035 ;
        RECT 58.455 208.615 58.785 208.865 ;
        RECT 57.360 208.445 58.785 208.615 ;
        RECT 59.015 208.235 59.185 208.695 ;
        RECT 59.445 208.365 59.615 208.865 ;
        RECT 56.815 208.065 59.185 208.235 ;
        RECT 56.815 207.895 56.985 208.065 ;
        RECT 59.435 207.895 59.640 208.185 ;
        RECT 59.875 208.115 61.085 209.205 ;
        RECT 56.680 207.565 56.985 207.895 ;
        RECT 57.180 207.845 57.430 207.895 ;
        RECT 57.640 207.845 57.910 207.895 ;
        RECT 57.175 207.675 57.430 207.845 ;
        RECT 57.635 207.675 57.910 207.845 ;
        RECT 57.180 207.565 57.430 207.675 ;
        RECT 56.815 207.395 56.985 207.565 ;
        RECT 56.815 207.225 57.375 207.395 ;
        RECT 57.640 207.235 57.910 207.675 ;
        RECT 58.100 207.505 58.390 207.895 ;
        RECT 58.095 207.335 58.390 207.505 ;
        RECT 58.100 207.235 58.390 207.335 ;
        RECT 58.560 207.230 58.980 207.895 ;
        RECT 59.290 207.845 59.640 207.895 ;
        RECT 59.290 207.675 59.645 207.845 ;
        RECT 59.290 207.565 59.640 207.675 ;
        RECT 59.875 207.405 60.395 207.945 ;
        RECT 60.565 207.575 61.085 208.115 ;
        RECT 56.200 206.870 56.535 207.130 ;
        RECT 57.205 207.055 57.375 207.225 ;
        RECT 56.705 206.655 57.035 207.055 ;
        RECT 57.205 206.885 58.820 207.055 ;
        RECT 59.365 206.655 59.695 207.375 ;
        RECT 59.875 206.655 61.085 207.405 ;
        RECT 61.265 206.835 61.525 209.025 ;
        RECT 61.695 208.475 62.035 209.205 ;
        RECT 62.215 208.295 62.485 209.025 ;
        RECT 61.715 208.075 62.485 208.295 ;
        RECT 62.665 208.315 62.895 209.025 ;
        RECT 63.065 208.495 63.395 209.205 ;
        RECT 63.565 208.315 63.825 209.025 ;
        RECT 62.665 208.075 63.825 208.315 ;
        RECT 61.715 207.405 62.005 208.075 ;
        RECT 64.945 208.065 65.275 209.205 ;
        RECT 65.805 208.235 66.135 209.020 ;
        RECT 65.455 208.065 66.135 208.235 ;
        RECT 62.185 207.585 62.650 207.895 ;
        RECT 62.830 207.585 63.355 207.895 ;
        RECT 61.715 207.205 62.945 207.405 ;
        RECT 61.785 206.655 62.455 207.025 ;
        RECT 62.635 206.835 62.945 207.205 ;
        RECT 63.125 206.945 63.355 207.585 ;
        RECT 63.535 207.565 63.835 207.895 ;
        RECT 64.935 207.645 65.285 207.895 ;
        RECT 65.455 207.465 65.625 208.065 ;
        RECT 67.235 208.040 67.525 209.205 ;
        RECT 67.695 208.115 68.905 209.205 ;
        RECT 65.795 207.645 66.145 207.895 ;
        RECT 63.535 206.655 63.825 207.385 ;
        RECT 64.945 206.655 65.215 207.465 ;
        RECT 65.385 206.825 65.715 207.465 ;
        RECT 65.885 206.655 66.125 207.465 ;
        RECT 67.695 207.405 68.215 207.945 ;
        RECT 68.385 207.575 68.905 208.115 ;
        RECT 69.075 208.605 69.335 209.025 ;
        RECT 69.505 208.775 69.835 209.205 ;
        RECT 70.500 208.775 71.245 208.945 ;
        RECT 71.470 208.865 72.110 209.025 ;
        RECT 69.075 208.435 70.905 208.605 ;
        RECT 67.235 206.655 67.525 207.380 ;
        RECT 67.695 206.655 68.905 207.405 ;
        RECT 69.075 207.395 69.245 208.435 ;
        RECT 69.415 207.565 69.765 208.265 ;
        RECT 69.980 208.095 70.565 208.265 ;
        RECT 69.935 207.565 70.225 207.895 ;
        RECT 70.395 207.815 70.565 208.095 ;
        RECT 70.735 208.155 70.905 208.435 ;
        RECT 71.075 208.525 71.245 208.775 ;
        RECT 71.435 208.695 72.110 208.865 ;
        RECT 71.075 208.355 72.110 208.525 ;
        RECT 72.280 208.405 72.560 209.205 ;
        RECT 71.940 208.235 72.110 208.355 ;
        RECT 70.735 207.985 71.385 208.155 ;
        RECT 71.940 208.065 72.600 208.235 ;
        RECT 72.770 208.065 73.045 209.035 ;
        RECT 70.395 207.645 70.820 207.815 ;
        RECT 70.395 207.395 70.565 207.645 ;
        RECT 71.215 207.565 71.385 207.985 ;
        RECT 72.430 207.895 72.600 208.065 ;
        RECT 71.605 207.565 72.260 207.895 ;
        RECT 72.430 207.565 72.705 207.895 ;
        RECT 72.430 207.395 72.600 207.565 ;
        RECT 69.075 207.020 69.390 207.395 ;
        RECT 69.645 206.655 69.815 207.395 ;
        RECT 70.065 207.225 70.565 207.395 ;
        RECT 71.005 207.225 72.600 207.395 ;
        RECT 72.875 207.330 73.045 208.065 ;
        RECT 70.065 207.020 70.235 207.225 ;
        RECT 70.460 206.655 70.835 207.055 ;
        RECT 71.005 206.875 71.175 207.225 ;
        RECT 71.360 206.655 71.690 207.055 ;
        RECT 71.860 206.875 72.030 207.225 ;
        RECT 72.200 206.655 72.580 207.055 ;
        RECT 72.770 206.985 73.045 207.330 ;
        RECT 73.225 208.145 73.555 208.995 ;
        RECT 73.225 207.380 73.415 208.145 ;
        RECT 73.725 208.065 73.975 209.205 ;
        RECT 74.165 208.565 74.415 208.985 ;
        RECT 74.645 208.735 74.975 209.205 ;
        RECT 75.205 208.565 75.455 208.985 ;
        RECT 74.165 208.395 75.455 208.565 ;
        RECT 75.635 208.565 75.965 208.995 ;
        RECT 75.635 208.395 76.090 208.565 ;
        RECT 74.155 207.895 74.370 208.225 ;
        RECT 73.585 207.565 73.895 207.895 ;
        RECT 74.065 207.565 74.370 207.895 ;
        RECT 74.545 207.565 74.830 208.225 ;
        RECT 75.025 207.565 75.290 208.225 ;
        RECT 75.505 207.565 75.750 208.225 ;
        RECT 73.725 207.395 73.895 207.565 ;
        RECT 75.920 207.395 76.090 208.395 ;
        RECT 73.225 206.870 73.555 207.380 ;
        RECT 73.725 207.225 76.090 207.395 ;
        RECT 76.445 208.145 76.775 208.995 ;
        RECT 76.445 207.380 76.635 208.145 ;
        RECT 76.945 208.065 77.195 209.205 ;
        RECT 77.385 208.565 77.635 208.985 ;
        RECT 77.865 208.735 78.195 209.205 ;
        RECT 78.425 208.565 78.675 208.985 ;
        RECT 77.385 208.395 78.675 208.565 ;
        RECT 78.855 208.565 79.185 208.995 ;
        RECT 78.855 208.395 79.310 208.565 ;
        RECT 77.375 207.895 77.590 208.225 ;
        RECT 76.805 207.565 77.115 207.895 ;
        RECT 77.285 207.565 77.590 207.895 ;
        RECT 77.765 207.565 78.050 208.225 ;
        RECT 78.245 207.565 78.510 208.225 ;
        RECT 78.725 207.565 78.970 208.225 ;
        RECT 76.945 207.395 77.115 207.565 ;
        RECT 79.140 207.395 79.310 208.395 ;
        RECT 79.655 208.115 80.865 209.205 ;
        RECT 73.725 206.655 74.055 207.055 ;
        RECT 75.105 206.885 75.435 207.225 ;
        RECT 75.605 206.655 75.935 207.055 ;
        RECT 76.445 206.870 76.775 207.380 ;
        RECT 76.945 207.225 79.310 207.395 ;
        RECT 79.655 207.405 80.175 207.945 ;
        RECT 80.345 207.575 80.865 208.115 ;
        RECT 81.045 208.145 81.375 208.995 ;
        RECT 76.945 206.655 77.275 207.055 ;
        RECT 78.325 206.885 78.655 207.225 ;
        RECT 78.825 206.655 79.155 207.055 ;
        RECT 79.655 206.655 80.865 207.405 ;
        RECT 81.045 207.380 81.235 208.145 ;
        RECT 81.545 208.065 81.795 209.205 ;
        RECT 81.985 208.565 82.235 208.985 ;
        RECT 82.465 208.735 82.795 209.205 ;
        RECT 83.025 208.565 83.275 208.985 ;
        RECT 81.985 208.395 83.275 208.565 ;
        RECT 83.455 208.565 83.785 208.995 ;
        RECT 83.455 208.395 83.910 208.565 ;
        RECT 81.975 207.895 82.190 208.225 ;
        RECT 81.405 207.565 81.715 207.895 ;
        RECT 81.885 207.565 82.190 207.895 ;
        RECT 82.365 207.565 82.650 208.225 ;
        RECT 82.845 207.565 83.110 208.225 ;
        RECT 83.325 207.565 83.570 208.225 ;
        RECT 81.545 207.395 81.715 207.565 ;
        RECT 83.740 207.395 83.910 208.395 ;
        RECT 84.805 208.235 84.975 209.035 ;
        RECT 85.735 208.575 85.985 209.035 ;
        RECT 86.185 208.825 86.855 209.205 ;
        RECT 87.045 208.575 87.295 209.035 ;
        RECT 87.470 208.745 87.715 209.205 ;
        RECT 85.735 208.405 87.295 208.575 ;
        RECT 87.885 208.355 88.225 208.995 ;
        RECT 84.805 208.065 87.745 208.235 ;
        RECT 87.575 207.895 87.745 208.065 ;
        RECT 84.775 207.565 84.960 207.895 ;
        RECT 85.215 207.565 85.690 207.895 ;
        RECT 86.000 207.565 86.345 207.895 ;
        RECT 81.045 206.870 81.375 207.380 ;
        RECT 81.545 207.225 83.910 207.395 ;
        RECT 84.805 207.225 85.985 207.395 ;
        RECT 86.155 207.335 86.345 207.565 ;
        RECT 86.605 207.320 86.800 207.895 ;
        RECT 87.070 207.565 87.405 207.895 ;
        RECT 87.575 207.565 87.885 207.895 ;
        RECT 87.575 207.395 87.745 207.565 ;
        RECT 81.545 206.655 81.875 207.055 ;
        RECT 82.925 206.885 83.255 207.225 ;
        RECT 83.425 206.655 83.755 207.055 ;
        RECT 84.805 206.825 84.975 207.225 ;
        RECT 85.215 206.655 85.545 207.055 ;
        RECT 85.815 206.995 85.985 207.225 ;
        RECT 87.050 207.225 87.745 207.395 ;
        RECT 88.055 207.240 88.225 208.355 ;
        RECT 88.395 208.115 91.905 209.205 ;
        RECT 87.050 206.995 87.220 207.225 ;
        RECT 85.815 206.825 87.220 206.995 ;
        RECT 87.390 206.655 87.720 207.035 ;
        RECT 87.915 206.825 88.225 207.240 ;
        RECT 88.395 207.425 90.045 207.945 ;
        RECT 90.215 207.595 91.905 208.115 ;
        RECT 92.995 208.040 93.285 209.205 ;
        RECT 93.915 208.650 94.520 209.205 ;
        RECT 94.695 208.695 95.175 209.035 ;
        RECT 95.345 208.660 95.600 209.205 ;
        RECT 93.915 208.550 94.530 208.650 ;
        RECT 94.345 208.525 94.530 208.550 ;
        RECT 93.915 207.930 94.175 208.380 ;
        RECT 94.345 208.280 94.675 208.525 ;
        RECT 94.845 208.205 95.600 208.455 ;
        RECT 95.770 208.335 96.045 209.035 ;
        RECT 94.830 208.170 95.600 208.205 ;
        RECT 94.815 208.160 95.600 208.170 ;
        RECT 94.810 208.145 95.705 208.160 ;
        RECT 94.790 208.130 95.705 208.145 ;
        RECT 94.770 208.120 95.705 208.130 ;
        RECT 94.745 208.110 95.705 208.120 ;
        RECT 94.675 208.080 95.705 208.110 ;
        RECT 94.655 208.050 95.705 208.080 ;
        RECT 94.635 208.020 95.705 208.050 ;
        RECT 94.605 207.995 95.705 208.020 ;
        RECT 94.570 207.960 95.705 207.995 ;
        RECT 94.540 207.955 95.705 207.960 ;
        RECT 94.540 207.950 94.930 207.955 ;
        RECT 94.540 207.940 94.905 207.950 ;
        RECT 94.540 207.935 94.890 207.940 ;
        RECT 94.540 207.930 94.875 207.935 ;
        RECT 93.915 207.925 94.875 207.930 ;
        RECT 93.915 207.915 94.865 207.925 ;
        RECT 93.915 207.910 94.855 207.915 ;
        RECT 93.915 207.900 94.845 207.910 ;
        RECT 93.915 207.890 94.840 207.900 ;
        RECT 93.915 207.885 94.835 207.890 ;
        RECT 93.915 207.870 94.825 207.885 ;
        RECT 93.915 207.855 94.820 207.870 ;
        RECT 93.915 207.830 94.810 207.855 ;
        RECT 93.915 207.760 94.805 207.830 ;
        RECT 88.395 206.655 91.905 207.425 ;
        RECT 92.995 206.655 93.285 207.380 ;
        RECT 93.915 207.205 94.465 207.590 ;
        RECT 94.635 207.035 94.805 207.760 ;
        RECT 93.915 206.865 94.805 207.035 ;
        RECT 94.975 207.360 95.305 207.785 ;
        RECT 95.475 207.560 95.705 207.955 ;
        RECT 94.975 206.875 95.195 207.360 ;
        RECT 95.875 207.305 96.045 208.335 ;
        RECT 96.215 208.065 96.495 209.205 ;
        RECT 96.665 208.055 96.995 209.035 ;
        RECT 97.165 208.065 97.425 209.205 ;
        RECT 97.595 208.115 100.185 209.205 ;
        RECT 96.225 207.625 96.560 207.895 ;
        RECT 96.730 207.455 96.900 208.055 ;
        RECT 97.070 207.645 97.405 207.895 ;
        RECT 95.365 206.655 95.615 207.195 ;
        RECT 95.785 206.825 96.045 207.305 ;
        RECT 96.215 206.655 96.525 207.455 ;
        RECT 96.730 206.825 97.425 207.455 ;
        RECT 97.595 207.425 98.805 207.945 ;
        RECT 98.975 207.595 100.185 208.115 ;
        RECT 100.365 208.145 100.695 208.995 ;
        RECT 97.595 206.655 100.185 207.425 ;
        RECT 100.365 207.380 100.555 208.145 ;
        RECT 100.865 208.065 101.115 209.205 ;
        RECT 101.305 208.565 101.555 208.985 ;
        RECT 101.785 208.735 102.115 209.205 ;
        RECT 102.345 208.565 102.595 208.985 ;
        RECT 101.305 208.395 102.595 208.565 ;
        RECT 102.775 208.565 103.105 208.995 ;
        RECT 102.775 208.395 103.230 208.565 ;
        RECT 101.295 207.895 101.510 208.225 ;
        RECT 100.725 207.565 101.035 207.895 ;
        RECT 101.205 207.565 101.510 207.895 ;
        RECT 101.685 207.565 101.970 208.225 ;
        RECT 102.165 207.565 102.430 208.225 ;
        RECT 102.645 207.565 102.890 208.225 ;
        RECT 100.865 207.395 101.035 207.565 ;
        RECT 103.060 207.395 103.230 208.395 ;
        RECT 103.665 208.235 103.835 209.035 ;
        RECT 104.595 208.575 104.845 209.035 ;
        RECT 105.045 208.825 105.715 209.205 ;
        RECT 105.905 208.575 106.155 209.035 ;
        RECT 106.330 208.745 106.575 209.205 ;
        RECT 104.595 208.405 106.155 208.575 ;
        RECT 106.745 208.355 107.085 208.995 ;
        RECT 103.665 208.065 106.605 208.235 ;
        RECT 106.435 207.895 106.605 208.065 ;
        RECT 103.635 207.565 103.820 207.895 ;
        RECT 104.075 207.565 104.550 207.895 ;
        RECT 104.860 207.565 105.205 207.895 ;
        RECT 100.365 206.870 100.695 207.380 ;
        RECT 100.865 207.225 103.230 207.395 ;
        RECT 103.665 207.225 104.845 207.395 ;
        RECT 105.015 207.335 105.205 207.565 ;
        RECT 105.465 207.320 105.660 207.895 ;
        RECT 105.930 207.565 106.265 207.895 ;
        RECT 106.435 207.565 106.745 207.895 ;
        RECT 106.435 207.395 106.605 207.565 ;
        RECT 100.865 206.655 101.195 207.055 ;
        RECT 102.245 206.885 102.575 207.225 ;
        RECT 102.745 206.655 103.075 207.055 ;
        RECT 103.665 206.825 103.835 207.225 ;
        RECT 104.075 206.655 104.405 207.055 ;
        RECT 104.675 206.995 104.845 207.225 ;
        RECT 105.910 207.225 106.605 207.395 ;
        RECT 106.915 207.240 107.085 208.355 ;
        RECT 105.910 206.995 106.080 207.225 ;
        RECT 104.675 206.825 106.080 206.995 ;
        RECT 106.250 206.655 106.580 207.035 ;
        RECT 106.775 206.825 107.085 207.240 ;
        RECT 107.265 208.145 107.595 208.995 ;
        RECT 107.265 208.015 107.485 208.145 ;
        RECT 107.765 208.065 108.015 209.205 ;
        RECT 108.205 208.565 108.455 208.985 ;
        RECT 108.685 208.735 109.015 209.205 ;
        RECT 109.245 208.565 109.495 208.985 ;
        RECT 108.205 208.395 109.495 208.565 ;
        RECT 109.675 208.565 110.005 208.995 ;
        RECT 109.675 208.395 110.130 208.565 ;
        RECT 107.265 207.380 107.455 208.015 ;
        RECT 108.195 207.895 108.410 208.225 ;
        RECT 107.625 207.565 107.935 207.895 ;
        RECT 108.105 207.565 108.410 207.895 ;
        RECT 108.585 207.565 108.870 208.225 ;
        RECT 109.065 207.565 109.330 208.225 ;
        RECT 109.545 207.565 109.790 208.225 ;
        RECT 107.765 207.395 107.935 207.565 ;
        RECT 109.960 207.395 110.130 208.395 ;
        RECT 107.265 206.870 107.595 207.380 ;
        RECT 107.765 207.225 110.130 207.395 ;
        RECT 110.485 208.145 110.815 208.995 ;
        RECT 110.485 207.380 110.675 208.145 ;
        RECT 110.985 208.065 111.235 209.205 ;
        RECT 111.425 208.565 111.675 208.985 ;
        RECT 111.905 208.735 112.235 209.205 ;
        RECT 112.465 208.565 112.715 208.985 ;
        RECT 111.425 208.395 112.715 208.565 ;
        RECT 112.895 208.565 113.225 208.995 ;
        RECT 114.155 208.735 114.495 208.995 ;
        RECT 114.665 208.745 114.915 209.205 ;
        RECT 112.895 208.395 113.350 208.565 ;
        RECT 111.415 207.895 111.630 208.225 ;
        RECT 110.845 207.565 111.155 207.895 ;
        RECT 111.325 207.565 111.630 207.895 ;
        RECT 111.805 207.565 112.090 208.225 ;
        RECT 112.285 207.565 112.550 208.225 ;
        RECT 112.765 207.565 113.010 208.225 ;
        RECT 110.985 207.395 111.155 207.565 ;
        RECT 113.180 207.395 113.350 208.395 ;
        RECT 107.765 206.655 108.095 207.055 ;
        RECT 109.145 206.885 109.475 207.225 ;
        RECT 109.645 206.655 109.975 207.055 ;
        RECT 110.485 206.870 110.815 207.380 ;
        RECT 110.985 207.225 113.350 207.395 ;
        RECT 110.985 206.655 111.315 207.055 ;
        RECT 112.365 206.885 112.695 207.225 ;
        RECT 114.155 207.130 114.415 208.735 ;
        RECT 115.105 208.565 115.435 208.995 ;
        RECT 114.585 208.395 115.435 208.565 ;
        RECT 115.605 208.535 115.775 209.035 ;
        RECT 115.985 208.745 116.235 209.205 ;
        RECT 116.445 208.535 116.615 209.035 ;
        RECT 116.915 208.745 117.165 209.205 ;
        RECT 117.405 208.535 117.575 209.035 ;
        RECT 114.585 207.475 114.755 208.395 ;
        RECT 115.605 208.365 117.575 208.535 ;
        RECT 115.075 207.645 115.405 208.205 ;
        RECT 115.605 208.185 115.905 208.190 ;
        RECT 115.595 208.015 115.905 208.185 ;
        RECT 115.605 207.895 115.905 208.015 ;
        RECT 115.605 207.565 115.985 207.895 ;
        RECT 114.585 207.380 115.405 207.475 ;
        RECT 114.585 207.305 115.600 207.380 ;
        RECT 112.865 206.655 113.195 207.055 ;
        RECT 114.155 206.870 114.495 207.130 ;
        RECT 114.665 206.655 114.995 207.135 ;
        RECT 115.185 206.870 115.600 207.305 ;
        RECT 116.295 207.170 116.515 207.895 ;
        RECT 116.775 207.565 117.155 208.195 ;
        RECT 117.385 207.565 117.640 208.195 ;
        RECT 118.755 208.040 119.045 209.205 ;
        RECT 119.215 208.065 119.475 209.205 ;
        RECT 119.645 208.055 119.975 209.035 ;
        RECT 120.145 208.065 120.425 209.205 ;
        RECT 120.595 208.115 121.805 209.205 ;
        RECT 119.235 207.645 119.570 207.895 ;
        RECT 115.770 206.985 116.720 207.170 ;
        RECT 116.950 206.965 117.155 207.565 ;
        RECT 119.740 207.455 119.910 208.055 ;
        RECT 120.080 207.625 120.415 207.895 ;
        RECT 117.325 206.655 117.665 207.380 ;
        RECT 118.755 206.655 119.045 207.380 ;
        RECT 119.215 206.825 119.910 207.455 ;
        RECT 120.115 206.655 120.425 207.455 ;
        RECT 120.595 207.405 121.115 207.945 ;
        RECT 121.285 207.575 121.805 208.115 ;
        RECT 120.595 206.655 121.805 207.405 ;
        RECT 121.975 206.935 122.255 209.035 ;
        RECT 122.445 208.445 123.230 209.205 ;
        RECT 123.625 208.375 124.010 209.035 ;
        RECT 123.625 208.275 124.035 208.375 ;
        RECT 122.425 208.065 124.035 208.275 ;
        RECT 124.335 208.185 124.535 208.975 ;
        RECT 122.425 207.465 122.700 208.065 ;
        RECT 124.205 208.015 124.535 208.185 ;
        RECT 124.705 208.025 125.025 209.205 ;
        RECT 125.195 208.770 130.540 209.205 ;
        RECT 124.205 207.895 124.385 208.015 ;
        RECT 122.870 207.645 123.225 207.895 ;
        RECT 123.420 207.845 123.885 207.895 ;
        RECT 123.415 207.675 123.885 207.845 ;
        RECT 123.420 207.645 123.885 207.675 ;
        RECT 124.055 207.645 124.385 207.895 ;
        RECT 124.560 207.645 125.025 207.845 ;
        RECT 122.425 207.285 123.675 207.465 ;
        RECT 123.310 207.215 123.675 207.285 ;
        RECT 123.845 207.265 125.025 207.435 ;
        RECT 122.485 206.655 122.655 207.115 ;
        RECT 123.845 207.045 124.175 207.265 ;
        RECT 122.925 206.865 124.175 207.045 ;
        RECT 124.345 206.655 124.515 207.095 ;
        RECT 124.685 206.850 125.025 207.265 ;
        RECT 126.780 207.200 127.120 208.030 ;
        RECT 128.600 207.520 128.950 208.770 ;
        RECT 130.720 208.695 132.375 208.985 ;
        RECT 130.720 208.355 132.310 208.525 ;
        RECT 132.545 208.405 132.825 209.205 ;
        RECT 130.720 208.065 131.040 208.355 ;
        RECT 132.140 208.235 132.310 208.355 ;
        RECT 130.720 207.325 131.070 207.895 ;
        RECT 131.240 207.565 131.950 208.185 ;
        RECT 132.140 208.065 132.865 208.235 ;
        RECT 133.035 208.065 133.305 209.035 ;
        RECT 132.695 207.895 132.865 208.065 ;
        RECT 132.120 207.565 132.525 207.895 ;
        RECT 132.695 207.565 132.965 207.895 ;
        RECT 132.695 207.395 132.865 207.565 ;
        RECT 131.255 207.225 132.865 207.395 ;
        RECT 133.135 207.330 133.305 208.065 ;
        RECT 125.195 206.655 130.540 207.200 ;
        RECT 130.725 206.655 131.055 207.155 ;
        RECT 131.255 206.875 131.425 207.225 ;
        RECT 131.625 206.655 131.955 207.055 ;
        RECT 132.125 206.875 132.295 207.225 ;
        RECT 132.465 206.655 132.845 207.055 ;
        RECT 133.035 206.985 133.305 207.330 ;
        RECT 133.485 206.835 133.745 209.025 ;
        RECT 133.915 208.475 134.255 209.205 ;
        RECT 134.435 208.295 134.705 209.025 ;
        RECT 133.935 208.075 134.705 208.295 ;
        RECT 134.885 208.315 135.115 209.025 ;
        RECT 135.285 208.495 135.615 209.205 ;
        RECT 135.785 208.315 136.045 209.025 ;
        RECT 136.235 208.770 141.580 209.205 ;
        RECT 134.885 208.075 136.045 208.315 ;
        RECT 133.935 207.405 134.225 208.075 ;
        RECT 134.405 207.585 134.870 207.895 ;
        RECT 135.050 207.585 135.575 207.895 ;
        RECT 133.935 207.205 135.165 207.405 ;
        RECT 134.005 206.655 134.675 207.025 ;
        RECT 134.855 206.835 135.165 207.205 ;
        RECT 135.345 206.945 135.575 207.585 ;
        RECT 135.755 207.565 136.055 207.895 ;
        RECT 135.755 206.655 136.045 207.385 ;
        RECT 137.820 207.200 138.160 208.030 ;
        RECT 139.640 207.520 139.990 208.770 ;
        RECT 141.755 208.115 144.345 209.205 ;
        RECT 141.755 207.425 142.965 207.945 ;
        RECT 143.135 207.595 144.345 208.115 ;
        RECT 144.515 208.040 144.805 209.205 ;
        RECT 144.975 208.065 145.360 209.025 ;
        RECT 145.575 208.405 145.865 209.205 ;
        RECT 146.035 208.865 147.400 209.035 ;
        RECT 146.035 208.235 146.205 208.865 ;
        RECT 145.530 208.065 146.205 208.235 ;
        RECT 136.235 206.655 141.580 207.200 ;
        RECT 141.755 206.655 144.345 207.425 ;
        RECT 144.975 207.395 145.150 208.065 ;
        RECT 145.530 207.895 145.700 208.065 ;
        RECT 146.375 207.895 146.700 208.695 ;
        RECT 147.070 208.655 147.400 208.865 ;
        RECT 147.070 208.405 148.025 208.655 ;
        RECT 145.335 207.645 145.700 207.895 ;
        RECT 145.895 207.645 146.145 207.895 ;
        RECT 145.335 207.565 145.525 207.645 ;
        RECT 145.895 207.565 146.065 207.645 ;
        RECT 146.355 207.565 146.700 207.895 ;
        RECT 146.870 207.565 147.145 208.230 ;
        RECT 147.330 207.565 147.685 208.230 ;
        RECT 147.855 207.395 148.025 208.405 ;
        RECT 148.195 208.065 148.485 209.205 ;
        RECT 149.575 208.050 149.915 209.035 ;
        RECT 150.085 208.775 150.495 209.205 ;
        RECT 151.240 208.785 151.570 209.205 ;
        RECT 151.740 208.605 152.065 209.035 ;
        RECT 150.085 208.435 152.065 208.605 ;
        RECT 148.210 207.565 148.485 207.895 ;
        RECT 144.515 206.655 144.805 207.380 ;
        RECT 144.975 206.825 145.485 207.395 ;
        RECT 146.030 207.225 147.430 207.395 ;
        RECT 145.655 206.655 145.825 207.215 ;
        RECT 146.030 206.825 146.360 207.225 ;
        RECT 146.535 206.655 146.865 207.055 ;
        RECT 147.100 207.035 147.430 207.225 ;
        RECT 147.600 207.205 148.025 207.395 ;
        RECT 149.575 207.395 149.830 208.050 ;
        RECT 150.085 207.895 150.350 208.435 ;
        RECT 150.565 208.095 151.190 208.265 ;
        RECT 150.000 207.565 150.350 207.895 ;
        RECT 150.520 207.565 150.850 207.895 ;
        RECT 151.020 207.395 151.190 208.095 ;
        RECT 148.195 207.035 148.485 207.305 ;
        RECT 147.100 206.825 148.485 207.035 ;
        RECT 149.575 207.020 149.935 207.395 ;
        RECT 150.200 206.655 150.370 207.395 ;
        RECT 150.650 207.225 151.190 207.395 ;
        RECT 151.360 208.025 152.065 208.435 ;
        RECT 152.540 208.105 152.870 209.205 ;
        RECT 153.255 208.335 153.530 209.035 ;
        RECT 153.700 208.660 153.955 209.205 ;
        RECT 154.125 208.695 154.605 209.035 ;
        RECT 154.780 208.650 155.385 209.205 ;
        RECT 154.770 208.550 155.385 208.650 ;
        RECT 154.770 208.525 154.955 208.550 ;
        RECT 150.650 207.020 150.820 207.225 ;
        RECT 151.360 206.825 151.530 208.025 ;
        RECT 151.700 207.645 152.270 207.855 ;
        RECT 152.440 207.645 153.085 207.855 ;
        RECT 151.760 207.305 152.930 207.475 ;
        RECT 151.760 206.825 152.090 207.305 ;
        RECT 152.260 206.655 152.430 207.125 ;
        RECT 152.600 206.840 152.930 207.305 ;
        RECT 153.255 207.305 153.425 208.335 ;
        RECT 153.700 208.205 154.455 208.455 ;
        RECT 154.625 208.280 154.955 208.525 ;
        RECT 153.700 208.170 154.470 208.205 ;
        RECT 153.700 208.160 154.485 208.170 ;
        RECT 153.595 208.145 154.490 208.160 ;
        RECT 153.595 208.130 154.510 208.145 ;
        RECT 153.595 208.120 154.530 208.130 ;
        RECT 153.595 208.110 154.555 208.120 ;
        RECT 153.595 208.080 154.625 208.110 ;
        RECT 153.595 208.050 154.645 208.080 ;
        RECT 153.595 208.020 154.665 208.050 ;
        RECT 153.595 207.995 154.695 208.020 ;
        RECT 153.595 207.960 154.730 207.995 ;
        RECT 153.595 207.955 154.760 207.960 ;
        RECT 153.595 207.560 153.825 207.955 ;
        RECT 154.370 207.950 154.760 207.955 ;
        RECT 154.395 207.940 154.760 207.950 ;
        RECT 154.410 207.935 154.760 207.940 ;
        RECT 154.425 207.930 154.760 207.935 ;
        RECT 155.125 207.930 155.385 208.380 ;
        RECT 155.555 208.115 156.765 209.205 ;
        RECT 154.425 207.925 155.385 207.930 ;
        RECT 154.435 207.915 155.385 207.925 ;
        RECT 154.445 207.910 155.385 207.915 ;
        RECT 154.455 207.900 155.385 207.910 ;
        RECT 154.460 207.890 155.385 207.900 ;
        RECT 154.465 207.885 155.385 207.890 ;
        RECT 154.475 207.870 155.385 207.885 ;
        RECT 154.480 207.855 155.385 207.870 ;
        RECT 154.490 207.830 155.385 207.855 ;
        RECT 153.995 207.360 154.325 207.785 ;
        RECT 154.075 207.335 154.325 207.360 ;
        RECT 153.255 206.825 153.515 207.305 ;
        RECT 153.685 206.655 153.935 207.195 ;
        RECT 154.105 206.875 154.325 207.335 ;
        RECT 154.495 207.760 155.385 207.830 ;
        RECT 154.495 207.035 154.665 207.760 ;
        RECT 154.835 207.205 155.385 207.590 ;
        RECT 155.555 207.405 156.075 207.945 ;
        RECT 156.245 207.575 156.765 208.115 ;
        RECT 156.935 208.115 158.145 209.205 ;
        RECT 156.935 207.575 157.455 208.115 ;
        RECT 157.625 207.405 158.145 207.945 ;
        RECT 154.495 206.865 155.385 207.035 ;
        RECT 155.555 206.655 156.765 207.405 ;
        RECT 156.935 206.655 158.145 207.405 ;
        RECT 2.750 206.485 158.230 206.655 ;
        RECT 2.835 205.735 4.045 206.485 ;
        RECT 4.765 205.935 4.935 206.315 ;
        RECT 5.115 206.105 5.445 206.485 ;
        RECT 4.765 205.765 5.430 205.935 ;
        RECT 5.625 205.810 5.885 206.315 ;
        RECT 2.835 205.195 3.355 205.735 ;
        RECT 3.525 205.025 4.045 205.565 ;
        RECT 4.695 205.215 5.025 205.585 ;
        RECT 5.260 205.510 5.430 205.765 ;
        RECT 5.260 205.180 5.545 205.510 ;
        RECT 5.260 205.035 5.430 205.180 ;
        RECT 2.835 203.935 4.045 205.025 ;
        RECT 4.765 204.865 5.430 205.035 ;
        RECT 5.715 205.010 5.885 205.810 ;
        RECT 4.765 204.105 4.935 204.865 ;
        RECT 5.115 203.935 5.445 204.695 ;
        RECT 5.615 204.105 5.885 205.010 ;
        RECT 6.055 205.810 6.315 206.315 ;
        RECT 6.495 206.105 6.825 206.485 ;
        RECT 7.005 205.935 7.175 206.315 ;
        RECT 6.055 205.010 6.225 205.810 ;
        RECT 6.510 205.765 7.175 205.935 ;
        RECT 6.510 205.510 6.680 205.765 ;
        RECT 7.440 205.745 7.695 206.315 ;
        RECT 7.865 206.085 8.195 206.485 ;
        RECT 8.620 205.950 9.150 206.315 ;
        RECT 8.620 205.915 8.795 205.950 ;
        RECT 7.865 205.745 8.795 205.915 ;
        RECT 9.340 205.805 9.615 206.315 ;
        RECT 6.395 205.180 6.680 205.510 ;
        RECT 6.915 205.215 7.245 205.585 ;
        RECT 6.510 205.035 6.680 205.180 ;
        RECT 7.440 205.075 7.610 205.745 ;
        RECT 7.865 205.575 8.035 205.745 ;
        RECT 7.780 205.245 8.035 205.575 ;
        RECT 8.260 205.245 8.455 205.575 ;
        RECT 6.055 204.105 6.325 205.010 ;
        RECT 6.510 204.865 7.175 205.035 ;
        RECT 6.495 203.935 6.825 204.695 ;
        RECT 7.005 204.105 7.175 204.865 ;
        RECT 7.440 204.105 7.775 205.075 ;
        RECT 7.945 203.935 8.115 205.075 ;
        RECT 8.285 204.275 8.455 205.245 ;
        RECT 8.625 204.615 8.795 205.745 ;
        RECT 8.965 204.955 9.135 205.755 ;
        RECT 9.335 205.635 9.615 205.805 ;
        RECT 9.340 205.155 9.615 205.635 ;
        RECT 9.785 204.955 9.975 206.315 ;
        RECT 10.155 205.950 10.665 206.485 ;
        RECT 10.885 205.675 11.130 206.280 ;
        RECT 11.850 205.675 12.095 206.280 ;
        RECT 12.315 205.950 12.825 206.485 ;
        RECT 10.175 205.505 11.405 205.675 ;
        RECT 8.965 204.785 9.975 204.955 ;
        RECT 10.145 204.940 10.895 205.130 ;
        RECT 8.625 204.445 9.750 204.615 ;
        RECT 10.145 204.275 10.315 204.940 ;
        RECT 11.065 204.695 11.405 205.505 ;
        RECT 8.285 204.105 10.315 204.275 ;
        RECT 10.485 203.935 10.655 204.695 ;
        RECT 10.890 204.285 11.405 204.695 ;
        RECT 11.575 205.505 12.805 205.675 ;
        RECT 11.575 204.695 11.915 205.505 ;
        RECT 12.085 204.940 12.835 205.130 ;
        RECT 11.575 204.285 12.090 204.695 ;
        RECT 12.325 203.935 12.495 204.695 ;
        RECT 12.665 204.275 12.835 204.940 ;
        RECT 13.005 204.955 13.195 206.315 ;
        RECT 13.365 205.465 13.640 206.315 ;
        RECT 13.830 205.950 14.360 206.315 ;
        RECT 14.785 206.085 15.115 206.485 ;
        RECT 14.185 205.915 14.360 205.950 ;
        RECT 13.365 205.295 13.645 205.465 ;
        RECT 13.365 205.155 13.640 205.295 ;
        RECT 13.845 204.955 14.015 205.755 ;
        RECT 13.005 204.785 14.015 204.955 ;
        RECT 14.185 205.745 15.115 205.915 ;
        RECT 15.285 205.745 15.540 206.315 ;
        RECT 14.185 204.615 14.355 205.745 ;
        RECT 14.945 205.575 15.115 205.745 ;
        RECT 13.230 204.445 14.355 204.615 ;
        RECT 14.525 205.245 14.720 205.575 ;
        RECT 14.945 205.245 15.200 205.575 ;
        RECT 14.525 204.275 14.695 205.245 ;
        RECT 15.370 205.075 15.540 205.745 ;
        RECT 12.665 204.105 14.695 204.275 ;
        RECT 14.865 203.935 15.035 205.075 ;
        RECT 15.205 204.105 15.540 205.075 ;
        RECT 15.720 205.745 15.975 206.315 ;
        RECT 16.145 206.085 16.475 206.485 ;
        RECT 16.900 205.950 17.430 206.315 ;
        RECT 16.900 205.915 17.075 205.950 ;
        RECT 16.145 205.745 17.075 205.915 ;
        RECT 15.720 205.075 15.890 205.745 ;
        RECT 16.145 205.575 16.315 205.745 ;
        RECT 16.060 205.245 16.315 205.575 ;
        RECT 16.540 205.245 16.735 205.575 ;
        RECT 15.720 204.105 16.055 205.075 ;
        RECT 16.225 203.935 16.395 205.075 ;
        RECT 16.565 204.275 16.735 205.245 ;
        RECT 16.905 204.615 17.075 205.745 ;
        RECT 17.245 204.955 17.415 205.755 ;
        RECT 17.620 205.465 17.895 206.315 ;
        RECT 17.615 205.295 17.895 205.465 ;
        RECT 17.620 205.155 17.895 205.295 ;
        RECT 18.065 204.955 18.255 206.315 ;
        RECT 18.435 205.950 18.945 206.485 ;
        RECT 19.165 205.675 19.410 206.280 ;
        RECT 19.860 205.745 20.115 206.315 ;
        RECT 20.285 206.085 20.615 206.485 ;
        RECT 21.040 205.950 21.570 206.315 ;
        RECT 21.760 206.145 22.035 206.315 ;
        RECT 21.755 205.975 22.035 206.145 ;
        RECT 21.040 205.915 21.215 205.950 ;
        RECT 20.285 205.745 21.215 205.915 ;
        RECT 18.455 205.505 19.685 205.675 ;
        RECT 17.245 204.785 18.255 204.955 ;
        RECT 18.425 204.940 19.175 205.130 ;
        RECT 16.905 204.445 18.030 204.615 ;
        RECT 18.425 204.275 18.595 204.940 ;
        RECT 19.345 204.695 19.685 205.505 ;
        RECT 16.565 204.105 18.595 204.275 ;
        RECT 18.765 203.935 18.935 204.695 ;
        RECT 19.170 204.285 19.685 204.695 ;
        RECT 19.860 205.075 20.030 205.745 ;
        RECT 20.285 205.575 20.455 205.745 ;
        RECT 20.200 205.245 20.455 205.575 ;
        RECT 20.680 205.245 20.875 205.575 ;
        RECT 19.860 204.105 20.195 205.075 ;
        RECT 20.365 203.935 20.535 205.075 ;
        RECT 20.705 204.275 20.875 205.245 ;
        RECT 21.045 204.615 21.215 205.745 ;
        RECT 21.385 204.955 21.555 205.755 ;
        RECT 21.760 205.155 22.035 205.975 ;
        RECT 22.205 204.955 22.395 206.315 ;
        RECT 22.575 205.950 23.085 206.485 ;
        RECT 23.305 205.675 23.550 206.280 ;
        RECT 24.000 205.745 24.255 206.315 ;
        RECT 24.425 206.085 24.755 206.485 ;
        RECT 25.180 205.950 25.710 206.315 ;
        RECT 25.180 205.915 25.355 205.950 ;
        RECT 24.425 205.745 25.355 205.915 ;
        RECT 25.900 205.805 26.175 206.315 ;
        RECT 22.595 205.505 23.825 205.675 ;
        RECT 21.385 204.785 22.395 204.955 ;
        RECT 22.565 204.940 23.315 205.130 ;
        RECT 21.045 204.445 22.170 204.615 ;
        RECT 22.565 204.275 22.735 204.940 ;
        RECT 23.485 204.695 23.825 205.505 ;
        RECT 20.705 204.105 22.735 204.275 ;
        RECT 22.905 203.935 23.075 204.695 ;
        RECT 23.310 204.285 23.825 204.695 ;
        RECT 24.000 205.075 24.170 205.745 ;
        RECT 24.425 205.575 24.595 205.745 ;
        RECT 24.340 205.245 24.595 205.575 ;
        RECT 24.820 205.245 25.015 205.575 ;
        RECT 24.000 204.105 24.335 205.075 ;
        RECT 24.505 203.935 24.675 205.075 ;
        RECT 24.845 204.275 25.015 205.245 ;
        RECT 25.185 204.615 25.355 205.745 ;
        RECT 25.525 204.955 25.695 205.755 ;
        RECT 25.895 205.635 26.175 205.805 ;
        RECT 25.900 205.155 26.175 205.635 ;
        RECT 26.345 204.955 26.535 206.315 ;
        RECT 26.715 205.950 27.225 206.485 ;
        RECT 27.445 205.675 27.690 206.280 ;
        RECT 28.595 205.760 28.885 206.485 ;
        RECT 29.075 205.675 29.315 206.485 ;
        RECT 29.485 205.675 29.815 206.315 ;
        RECT 29.985 205.675 30.255 206.485 ;
        RECT 30.435 205.985 30.735 206.315 ;
        RECT 30.905 206.005 31.180 206.485 ;
        RECT 26.735 205.505 27.965 205.675 ;
        RECT 25.525 204.785 26.535 204.955 ;
        RECT 26.705 204.940 27.455 205.130 ;
        RECT 25.185 204.445 26.310 204.615 ;
        RECT 26.705 204.275 26.875 204.940 ;
        RECT 27.625 204.695 27.965 205.505 ;
        RECT 29.055 205.245 29.405 205.495 ;
        RECT 24.845 204.105 26.875 204.275 ;
        RECT 27.045 203.935 27.215 204.695 ;
        RECT 27.450 204.285 27.965 204.695 ;
        RECT 28.595 203.935 28.885 205.100 ;
        RECT 29.575 205.075 29.745 205.675 ;
        RECT 29.915 205.245 30.265 205.495 ;
        RECT 30.435 205.075 30.605 205.985 ;
        RECT 31.360 205.835 31.655 206.225 ;
        RECT 31.825 206.005 32.080 206.485 ;
        RECT 32.255 205.835 32.515 206.225 ;
        RECT 32.685 206.005 32.965 206.485 ;
        RECT 30.775 205.245 31.125 205.815 ;
        RECT 31.360 205.665 33.010 205.835 ;
        RECT 31.295 205.325 32.435 205.495 ;
        RECT 31.295 205.075 31.465 205.325 ;
        RECT 32.605 205.155 33.010 205.665 ;
        RECT 29.065 204.905 29.745 205.075 ;
        RECT 29.065 204.120 29.395 204.905 ;
        RECT 29.925 203.935 30.255 205.075 ;
        RECT 30.435 204.905 31.465 205.075 ;
        RECT 32.255 204.985 33.010 205.155 ;
        RECT 33.200 205.775 33.455 206.305 ;
        RECT 33.625 206.025 33.930 206.485 ;
        RECT 34.175 206.105 35.245 206.275 ;
        RECT 33.200 205.125 33.410 205.775 ;
        RECT 34.175 205.750 34.495 206.105 ;
        RECT 34.170 205.575 34.495 205.750 ;
        RECT 33.580 205.275 34.495 205.575 ;
        RECT 34.665 205.535 34.905 205.935 ;
        RECT 35.075 205.875 35.245 206.105 ;
        RECT 35.415 206.045 35.605 206.485 ;
        RECT 35.775 206.035 36.725 206.315 ;
        RECT 36.945 206.125 37.295 206.295 ;
        RECT 35.075 205.705 35.605 205.875 ;
        RECT 33.580 205.245 34.320 205.275 ;
        RECT 30.435 204.105 30.745 204.905 ;
        RECT 32.255 204.735 32.515 204.985 ;
        RECT 30.915 203.935 31.225 204.735 ;
        RECT 31.395 204.565 32.515 204.735 ;
        RECT 31.395 204.105 31.655 204.565 ;
        RECT 31.825 203.935 32.080 204.395 ;
        RECT 32.255 204.105 32.515 204.565 ;
        RECT 32.685 203.935 32.970 204.805 ;
        RECT 33.200 204.245 33.455 205.125 ;
        RECT 33.625 203.935 33.930 205.075 ;
        RECT 34.150 204.655 34.320 205.245 ;
        RECT 34.665 205.165 35.205 205.535 ;
        RECT 35.385 205.425 35.605 205.705 ;
        RECT 35.775 205.255 35.945 206.035 ;
        RECT 35.540 205.085 35.945 205.255 ;
        RECT 36.115 205.245 36.465 205.865 ;
        RECT 35.540 204.995 35.710 205.085 ;
        RECT 36.635 205.075 36.845 205.865 ;
        RECT 34.490 204.825 35.710 204.995 ;
        RECT 36.170 204.915 36.845 205.075 ;
        RECT 34.150 204.485 34.950 204.655 ;
        RECT 34.270 203.935 34.600 204.315 ;
        RECT 34.780 204.195 34.950 204.485 ;
        RECT 35.540 204.445 35.710 204.825 ;
        RECT 35.880 204.905 36.845 204.915 ;
        RECT 37.035 205.735 37.295 206.125 ;
        RECT 37.505 206.025 37.835 206.485 ;
        RECT 38.710 206.095 39.565 206.265 ;
        RECT 39.770 206.095 40.265 206.265 ;
        RECT 40.435 206.125 40.765 206.485 ;
        RECT 37.035 205.045 37.205 205.735 ;
        RECT 37.375 205.385 37.545 205.565 ;
        RECT 37.715 205.555 38.505 205.805 ;
        RECT 38.710 205.385 38.880 206.095 ;
        RECT 39.050 205.585 39.405 205.805 ;
        RECT 37.375 205.215 39.065 205.385 ;
        RECT 35.880 204.615 36.340 204.905 ;
        RECT 37.035 204.875 38.535 205.045 ;
        RECT 37.035 204.735 37.205 204.875 ;
        RECT 36.645 204.565 37.205 204.735 ;
        RECT 35.120 203.935 35.370 204.395 ;
        RECT 35.540 204.105 36.410 204.445 ;
        RECT 36.645 204.105 36.815 204.565 ;
        RECT 37.650 204.535 38.725 204.705 ;
        RECT 36.985 203.935 37.355 204.395 ;
        RECT 37.650 204.195 37.820 204.535 ;
        RECT 37.990 203.935 38.320 204.365 ;
        RECT 38.555 204.195 38.725 204.535 ;
        RECT 38.895 204.435 39.065 205.215 ;
        RECT 39.235 204.995 39.405 205.585 ;
        RECT 39.575 205.185 39.925 205.805 ;
        RECT 39.235 204.605 39.700 204.995 ;
        RECT 40.095 204.735 40.265 206.095 ;
        RECT 40.435 204.905 40.895 205.955 ;
        RECT 39.870 204.565 40.265 204.735 ;
        RECT 39.870 204.435 40.040 204.565 ;
        RECT 38.895 204.105 39.575 204.435 ;
        RECT 39.790 204.105 40.040 204.435 ;
        RECT 40.210 203.935 40.460 204.395 ;
        RECT 40.630 204.120 40.955 204.905 ;
        RECT 41.125 204.105 41.295 206.225 ;
        RECT 41.465 206.105 41.795 206.485 ;
        RECT 41.965 205.935 42.220 206.225 ;
        RECT 41.470 205.765 42.220 205.935 ;
        RECT 41.470 204.775 41.700 205.765 ;
        RECT 42.400 205.745 42.655 206.315 ;
        RECT 42.825 206.085 43.155 206.485 ;
        RECT 43.580 205.950 44.110 206.315 ;
        RECT 43.580 205.915 43.755 205.950 ;
        RECT 42.825 205.745 43.755 205.915 ;
        RECT 41.870 204.945 42.220 205.595 ;
        RECT 42.400 205.075 42.570 205.745 ;
        RECT 42.825 205.575 42.995 205.745 ;
        RECT 42.740 205.245 42.995 205.575 ;
        RECT 43.220 205.245 43.415 205.575 ;
        RECT 41.470 204.605 42.220 204.775 ;
        RECT 41.465 203.935 41.795 204.435 ;
        RECT 41.965 204.105 42.220 204.605 ;
        RECT 42.400 204.105 42.735 205.075 ;
        RECT 42.905 203.935 43.075 205.075 ;
        RECT 43.245 204.275 43.415 205.245 ;
        RECT 43.585 204.615 43.755 205.745 ;
        RECT 43.925 204.955 44.095 205.755 ;
        RECT 44.300 205.465 44.575 206.315 ;
        RECT 44.295 205.295 44.575 205.465 ;
        RECT 44.300 205.155 44.575 205.295 ;
        RECT 44.745 204.955 44.935 206.315 ;
        RECT 45.115 205.950 45.625 206.485 ;
        RECT 45.845 205.675 46.090 206.280 ;
        RECT 46.810 205.675 47.055 206.280 ;
        RECT 47.275 205.950 47.785 206.485 ;
        RECT 45.135 205.505 46.365 205.675 ;
        RECT 43.925 204.785 44.935 204.955 ;
        RECT 45.105 204.940 45.855 205.130 ;
        RECT 43.585 204.445 44.710 204.615 ;
        RECT 45.105 204.275 45.275 204.940 ;
        RECT 46.025 204.695 46.365 205.505 ;
        RECT 43.245 204.105 45.275 204.275 ;
        RECT 45.445 203.935 45.615 204.695 ;
        RECT 45.850 204.285 46.365 204.695 ;
        RECT 46.535 205.505 47.765 205.675 ;
        RECT 46.535 204.695 46.875 205.505 ;
        RECT 47.045 204.940 47.795 205.130 ;
        RECT 46.535 204.285 47.050 204.695 ;
        RECT 47.285 203.935 47.455 204.695 ;
        RECT 47.625 204.275 47.795 204.940 ;
        RECT 47.965 204.955 48.155 206.315 ;
        RECT 48.325 205.465 48.600 206.315 ;
        RECT 48.790 205.950 49.320 206.315 ;
        RECT 49.745 206.085 50.075 206.485 ;
        RECT 49.145 205.915 49.320 205.950 ;
        RECT 48.325 205.295 48.605 205.465 ;
        RECT 48.325 205.155 48.600 205.295 ;
        RECT 48.805 204.955 48.975 205.755 ;
        RECT 47.965 204.785 48.975 204.955 ;
        RECT 49.145 205.745 50.075 205.915 ;
        RECT 50.245 205.745 50.500 206.315 ;
        RECT 49.145 204.615 49.315 205.745 ;
        RECT 49.905 205.575 50.075 205.745 ;
        RECT 48.190 204.445 49.315 204.615 ;
        RECT 49.485 205.245 49.680 205.575 ;
        RECT 49.905 205.245 50.160 205.575 ;
        RECT 49.485 204.275 49.655 205.245 ;
        RECT 50.330 205.075 50.500 205.745 ;
        RECT 47.625 204.105 49.655 204.275 ;
        RECT 49.825 203.935 49.995 205.075 ;
        RECT 50.165 204.105 50.500 205.075 ;
        RECT 50.675 205.745 51.060 206.315 ;
        RECT 51.230 206.025 51.555 206.485 ;
        RECT 52.075 205.855 52.355 206.315 ;
        RECT 50.675 205.075 50.955 205.745 ;
        RECT 51.230 205.685 52.355 205.855 ;
        RECT 51.230 205.575 51.680 205.685 ;
        RECT 51.125 205.245 51.680 205.575 ;
        RECT 52.545 205.515 52.945 206.315 ;
        RECT 53.345 206.025 53.615 206.485 ;
        RECT 53.785 205.855 54.070 206.315 ;
        RECT 50.675 204.105 51.060 205.075 ;
        RECT 51.230 204.785 51.680 205.245 ;
        RECT 51.850 204.955 52.945 205.515 ;
        RECT 51.230 204.565 52.355 204.785 ;
        RECT 51.230 203.935 51.555 204.395 ;
        RECT 52.075 204.105 52.355 204.565 ;
        RECT 52.545 204.105 52.945 204.955 ;
        RECT 53.115 205.685 54.070 205.855 ;
        RECT 54.355 205.760 54.645 206.485 ;
        RECT 53.115 204.785 53.325 205.685 ;
        RECT 54.930 205.570 55.100 206.485 ;
        RECT 55.270 205.810 55.545 206.155 ;
        RECT 55.735 206.085 56.115 206.485 ;
        RECT 56.285 205.915 56.455 206.265 ;
        RECT 56.625 206.085 56.955 206.485 ;
        RECT 57.155 205.915 57.325 206.265 ;
        RECT 57.525 205.985 57.860 206.485 ;
        RECT 53.495 204.955 54.185 205.515 ;
        RECT 53.115 204.565 54.070 204.785 ;
        RECT 53.345 203.935 53.615 204.395 ;
        RECT 53.785 204.105 54.070 204.565 ;
        RECT 54.355 203.935 54.645 205.100 ;
        RECT 54.930 203.935 55.100 205.115 ;
        RECT 55.270 205.075 55.440 205.810 ;
        RECT 55.715 205.745 57.325 205.915 ;
        RECT 55.715 205.575 55.885 205.745 ;
        RECT 55.610 205.245 55.885 205.575 ;
        RECT 56.055 205.245 56.460 205.575 ;
        RECT 55.715 205.075 55.885 205.245 ;
        RECT 56.630 205.125 57.340 205.575 ;
        RECT 57.510 205.245 57.865 205.815 ;
        RECT 58.055 205.675 58.295 206.485 ;
        RECT 58.465 205.675 58.795 206.315 ;
        RECT 58.965 205.675 59.235 206.485 ;
        RECT 59.415 205.940 64.760 206.485 ;
        RECT 58.035 205.245 58.385 205.495 ;
        RECT 55.270 204.105 55.545 205.075 ;
        RECT 55.715 204.905 56.440 205.075 ;
        RECT 56.630 204.955 57.345 205.125 ;
        RECT 58.555 205.075 58.725 205.675 ;
        RECT 58.895 205.245 59.245 205.495 ;
        RECT 61.000 205.110 61.340 205.940 ;
        RECT 64.935 205.715 67.525 206.485 ;
        RECT 67.695 205.855 68.035 206.315 ;
        RECT 68.205 206.025 68.375 206.485 ;
        RECT 68.545 206.105 69.715 206.315 ;
        RECT 68.545 205.855 68.795 206.105 ;
        RECT 69.385 206.085 69.715 206.105 ;
        RECT 69.995 205.940 75.340 206.485 ;
        RECT 56.270 204.785 56.440 204.905 ;
        RECT 57.540 204.785 57.865 205.075 ;
        RECT 55.755 203.935 56.035 204.735 ;
        RECT 56.270 204.615 57.865 204.785 ;
        RECT 58.045 204.905 58.725 205.075 ;
        RECT 56.205 204.155 57.865 204.445 ;
        RECT 58.045 204.120 58.375 204.905 ;
        RECT 58.905 203.935 59.235 205.075 ;
        RECT 62.820 204.370 63.170 205.620 ;
        RECT 64.935 205.195 66.145 205.715 ;
        RECT 67.695 205.685 68.795 205.855 ;
        RECT 68.965 205.665 69.825 205.915 ;
        RECT 66.315 205.025 67.525 205.545 ;
        RECT 67.695 205.245 68.455 205.495 ;
        RECT 68.625 205.245 69.375 205.495 ;
        RECT 69.545 205.075 69.825 205.665 ;
        RECT 71.580 205.110 71.920 205.940 ;
        RECT 75.515 205.715 79.025 206.485 ;
        RECT 80.115 205.760 80.405 206.485 ;
        RECT 80.575 205.715 84.085 206.485 ;
        RECT 59.415 203.935 64.760 204.370 ;
        RECT 64.935 203.935 67.525 205.025 ;
        RECT 67.695 203.935 67.955 205.075 ;
        RECT 68.125 204.905 69.825 205.075 ;
        RECT 68.125 204.105 68.455 204.905 ;
        RECT 68.625 203.935 68.795 204.735 ;
        RECT 68.965 204.105 69.295 204.905 ;
        RECT 69.465 203.935 69.720 204.735 ;
        RECT 73.400 204.370 73.750 205.620 ;
        RECT 75.515 205.195 77.165 205.715 ;
        RECT 77.335 205.025 79.025 205.545 ;
        RECT 80.575 205.195 82.225 205.715 ;
        RECT 84.920 205.705 85.420 206.315 ;
        RECT 69.995 203.935 75.340 204.370 ;
        RECT 75.515 203.935 79.025 205.025 ;
        RECT 80.115 203.935 80.405 205.100 ;
        RECT 82.395 205.025 84.085 205.545 ;
        RECT 84.715 205.245 85.065 205.495 ;
        RECT 85.250 205.075 85.420 205.705 ;
        RECT 86.050 205.835 86.380 206.315 ;
        RECT 86.550 206.025 86.775 206.485 ;
        RECT 86.945 205.835 87.275 206.315 ;
        RECT 86.050 205.665 87.275 205.835 ;
        RECT 87.465 205.685 87.715 206.485 ;
        RECT 87.885 205.685 88.225 206.315 ;
        RECT 85.590 205.295 85.920 205.495 ;
        RECT 86.090 205.295 86.420 205.495 ;
        RECT 86.590 205.295 87.010 205.495 ;
        RECT 87.185 205.325 87.880 205.495 ;
        RECT 87.185 205.075 87.355 205.325 ;
        RECT 88.050 205.075 88.225 205.685 ;
        RECT 80.575 203.935 84.085 205.025 ;
        RECT 84.920 204.905 87.355 205.075 ;
        RECT 84.920 204.105 85.250 204.905 ;
        RECT 85.420 203.935 85.750 204.735 ;
        RECT 86.050 204.105 86.380 204.905 ;
        RECT 87.025 203.935 87.275 204.735 ;
        RECT 87.545 203.935 87.715 205.075 ;
        RECT 87.885 204.105 88.225 205.075 ;
        RECT 88.865 205.760 89.195 206.270 ;
        RECT 89.365 206.085 89.695 206.485 ;
        RECT 90.745 205.915 91.075 206.255 ;
        RECT 91.245 206.085 91.575 206.485 ;
        RECT 88.865 204.995 89.055 205.760 ;
        RECT 89.365 205.745 91.730 205.915 ;
        RECT 89.365 205.575 89.535 205.745 ;
        RECT 89.225 205.245 89.535 205.575 ;
        RECT 89.705 205.245 90.010 205.575 ;
        RECT 88.865 204.145 89.195 204.995 ;
        RECT 89.365 203.935 89.615 205.075 ;
        RECT 89.795 204.915 90.010 205.245 ;
        RECT 90.185 204.915 90.470 205.575 ;
        RECT 90.665 204.915 90.930 205.575 ;
        RECT 91.145 204.915 91.390 205.575 ;
        RECT 91.560 204.745 91.730 205.745 ;
        RECT 92.075 205.715 94.665 206.485 ;
        RECT 92.075 205.195 93.285 205.715 ;
        RECT 95.500 205.705 96.000 206.315 ;
        RECT 93.455 205.025 94.665 205.545 ;
        RECT 95.295 205.245 95.645 205.495 ;
        RECT 95.830 205.075 96.000 205.705 ;
        RECT 96.630 205.835 96.960 206.315 ;
        RECT 97.130 206.025 97.355 206.485 ;
        RECT 97.525 205.835 97.855 206.315 ;
        RECT 96.630 205.665 97.855 205.835 ;
        RECT 98.045 205.685 98.295 206.485 ;
        RECT 98.465 205.685 98.805 206.315 ;
        RECT 96.170 205.295 96.500 205.495 ;
        RECT 96.670 205.295 97.000 205.495 ;
        RECT 97.170 205.295 97.590 205.495 ;
        RECT 97.765 205.325 98.460 205.495 ;
        RECT 97.765 205.075 97.935 205.325 ;
        RECT 98.630 205.075 98.805 205.685 ;
        RECT 89.805 204.575 91.095 204.745 ;
        RECT 89.805 204.155 90.055 204.575 ;
        RECT 90.285 203.935 90.615 204.405 ;
        RECT 90.845 204.155 91.095 204.575 ;
        RECT 91.275 204.575 91.730 204.745 ;
        RECT 91.275 204.145 91.605 204.575 ;
        RECT 92.075 203.935 94.665 205.025 ;
        RECT 95.500 204.905 97.935 205.075 ;
        RECT 95.500 204.105 95.830 204.905 ;
        RECT 96.000 203.935 96.330 204.735 ;
        RECT 96.630 204.105 96.960 204.905 ;
        RECT 97.605 203.935 97.855 204.735 ;
        RECT 98.125 203.935 98.295 205.075 ;
        RECT 98.465 204.105 98.805 205.075 ;
        RECT 98.975 205.745 99.485 206.315 ;
        RECT 99.655 205.925 99.825 206.485 ;
        RECT 100.030 205.915 100.360 206.315 ;
        RECT 100.535 206.085 100.865 206.485 ;
        RECT 101.100 206.105 102.485 206.315 ;
        RECT 101.100 205.915 101.430 206.105 ;
        RECT 100.030 205.745 101.430 205.915 ;
        RECT 101.600 205.745 102.025 205.935 ;
        RECT 102.195 205.835 102.485 206.105 ;
        RECT 102.670 205.915 102.925 206.265 ;
        RECT 103.095 206.085 103.425 206.485 ;
        RECT 103.595 205.915 103.765 206.265 ;
        RECT 103.935 206.085 104.315 206.485 ;
        RECT 102.670 205.745 104.335 205.915 ;
        RECT 104.505 205.810 104.780 206.155 ;
        RECT 98.975 205.075 99.150 205.745 ;
        RECT 99.335 205.495 99.525 205.575 ;
        RECT 99.895 205.495 100.065 205.575 ;
        RECT 99.335 205.245 99.700 205.495 ;
        RECT 99.895 205.245 100.145 205.495 ;
        RECT 100.355 205.245 100.700 205.575 ;
        RECT 99.530 205.075 99.700 205.245 ;
        RECT 98.975 204.115 99.360 205.075 ;
        RECT 99.530 204.905 100.205 205.075 ;
        RECT 99.575 203.935 99.865 204.735 ;
        RECT 100.035 204.275 100.205 204.905 ;
        RECT 100.375 204.445 100.700 205.245 ;
        RECT 100.870 204.910 101.145 205.575 ;
        RECT 101.330 204.910 101.685 205.575 ;
        RECT 101.855 204.735 102.025 205.745 ;
        RECT 104.165 205.575 104.335 205.745 ;
        RECT 102.210 205.245 102.485 205.575 ;
        RECT 102.655 205.245 103.000 205.575 ;
        RECT 103.170 205.245 103.995 205.575 ;
        RECT 104.165 205.245 104.440 205.575 ;
        RECT 101.070 204.485 102.025 204.735 ;
        RECT 101.070 204.275 101.400 204.485 ;
        RECT 100.035 204.105 101.400 204.275 ;
        RECT 102.195 203.935 102.485 205.075 ;
        RECT 102.675 204.785 103.000 205.075 ;
        RECT 103.170 204.955 103.365 205.245 ;
        RECT 104.165 205.075 104.335 205.245 ;
        RECT 104.610 205.075 104.780 205.810 ;
        RECT 105.875 205.760 106.165 206.485 ;
        RECT 106.335 205.715 108.005 206.485 ;
        RECT 106.335 205.195 107.085 205.715 ;
        RECT 108.195 205.675 108.435 206.485 ;
        RECT 108.605 205.675 108.935 206.315 ;
        RECT 109.105 205.675 109.375 206.485 ;
        RECT 109.885 206.085 110.215 206.485 ;
        RECT 110.385 205.915 110.715 206.255 ;
        RECT 111.765 206.085 112.095 206.485 ;
        RECT 109.730 205.745 112.095 205.915 ;
        RECT 112.265 205.760 112.595 206.270 ;
        RECT 103.675 204.905 104.335 205.075 ;
        RECT 103.675 204.785 103.845 204.905 ;
        RECT 102.675 204.615 103.845 204.785 ;
        RECT 102.655 204.155 103.845 204.445 ;
        RECT 104.015 203.935 104.295 204.735 ;
        RECT 104.505 204.105 104.780 205.075 ;
        RECT 105.875 203.935 106.165 205.100 ;
        RECT 107.255 205.025 108.005 205.545 ;
        RECT 108.175 205.245 108.525 205.495 ;
        RECT 108.695 205.075 108.865 205.675 ;
        RECT 109.035 205.245 109.385 205.495 ;
        RECT 106.335 203.935 108.005 205.025 ;
        RECT 108.185 204.905 108.865 205.075 ;
        RECT 108.185 204.120 108.515 204.905 ;
        RECT 109.045 203.935 109.375 205.075 ;
        RECT 109.730 204.745 109.900 205.745 ;
        RECT 111.925 205.575 112.095 205.745 ;
        RECT 110.070 204.915 110.315 205.575 ;
        RECT 110.530 204.915 110.795 205.575 ;
        RECT 110.990 204.915 111.275 205.575 ;
        RECT 111.450 205.245 111.755 205.575 ;
        RECT 111.925 205.245 112.235 205.575 ;
        RECT 111.450 204.915 111.665 205.245 ;
        RECT 109.730 204.575 110.185 204.745 ;
        RECT 109.855 204.145 110.185 204.575 ;
        RECT 110.365 204.575 111.655 204.745 ;
        RECT 110.365 204.155 110.615 204.575 ;
        RECT 110.845 203.935 111.175 204.405 ;
        RECT 111.405 204.155 111.655 204.575 ;
        RECT 111.845 203.935 112.095 205.075 ;
        RECT 112.405 204.995 112.595 205.760 ;
        RECT 112.975 205.855 113.305 206.215 ;
        RECT 113.925 206.025 114.175 206.485 ;
        RECT 114.345 206.025 114.905 206.315 ;
        RECT 112.975 205.665 114.365 205.855 ;
        RECT 114.195 205.575 114.365 205.665 ;
        RECT 112.265 204.145 112.595 204.995 ;
        RECT 112.790 205.245 113.465 205.495 ;
        RECT 113.685 205.245 114.025 205.495 ;
        RECT 114.195 205.245 114.485 205.575 ;
        RECT 112.790 204.885 113.055 205.245 ;
        RECT 114.195 204.995 114.365 205.245 ;
        RECT 113.425 204.825 114.365 204.995 ;
        RECT 112.975 203.935 113.255 204.605 ;
        RECT 113.425 204.275 113.725 204.825 ;
        RECT 114.655 204.655 114.905 206.025 ;
        RECT 115.075 205.940 120.420 206.485 ;
        RECT 116.660 205.110 117.000 205.940 ;
        RECT 120.595 205.715 123.185 206.485 ;
        RECT 123.825 205.760 124.155 206.270 ;
        RECT 124.325 206.085 124.655 206.485 ;
        RECT 125.705 205.915 126.035 206.255 ;
        RECT 126.205 206.085 126.535 206.485 ;
        RECT 113.925 203.935 114.255 204.655 ;
        RECT 114.445 204.105 114.905 204.655 ;
        RECT 118.480 204.370 118.830 205.620 ;
        RECT 120.595 205.195 121.805 205.715 ;
        RECT 121.975 205.025 123.185 205.545 ;
        RECT 115.075 203.935 120.420 204.370 ;
        RECT 120.595 203.935 123.185 205.025 ;
        RECT 123.825 204.995 124.015 205.760 ;
        RECT 124.325 205.745 126.690 205.915 ;
        RECT 124.325 205.575 124.495 205.745 ;
        RECT 124.185 205.245 124.495 205.575 ;
        RECT 124.665 205.245 124.970 205.575 ;
        RECT 123.825 204.145 124.155 204.995 ;
        RECT 124.325 203.935 124.575 205.075 ;
        RECT 124.755 204.915 124.970 205.245 ;
        RECT 125.145 204.915 125.430 205.575 ;
        RECT 125.625 204.915 125.890 205.575 ;
        RECT 126.105 204.915 126.350 205.575 ;
        RECT 126.520 204.745 126.690 205.745 ;
        RECT 127.035 205.715 130.545 206.485 ;
        RECT 131.635 205.760 131.925 206.485 ;
        RECT 132.095 205.735 133.305 206.485 ;
        RECT 127.035 205.195 128.685 205.715 ;
        RECT 128.855 205.025 130.545 205.545 ;
        RECT 132.095 205.195 132.615 205.735 ;
        RECT 133.475 205.685 133.785 206.485 ;
        RECT 133.990 205.685 134.685 206.315 ;
        RECT 134.860 205.955 135.150 206.305 ;
        RECT 135.345 206.125 135.675 206.485 ;
        RECT 135.845 205.955 136.075 206.260 ;
        RECT 134.860 205.785 136.075 205.955 ;
        RECT 124.765 204.575 126.055 204.745 ;
        RECT 124.765 204.155 125.015 204.575 ;
        RECT 125.245 203.935 125.575 204.405 ;
        RECT 125.805 204.155 126.055 204.575 ;
        RECT 126.235 204.575 126.690 204.745 ;
        RECT 126.235 204.145 126.565 204.575 ;
        RECT 127.035 203.935 130.545 205.025 ;
        RECT 131.635 203.935 131.925 205.100 ;
        RECT 132.785 205.025 133.305 205.565 ;
        RECT 133.485 205.245 133.820 205.515 ;
        RECT 133.990 205.085 134.160 205.685 ;
        RECT 136.265 205.615 136.435 206.180 ;
        RECT 136.695 205.940 142.040 206.485 ;
        RECT 134.330 205.245 134.665 205.495 ;
        RECT 134.920 205.465 135.180 205.575 ;
        RECT 134.915 205.295 135.180 205.465 ;
        RECT 134.920 205.245 135.180 205.295 ;
        RECT 135.360 205.245 135.745 205.575 ;
        RECT 135.915 205.445 136.435 205.615 ;
        RECT 132.095 203.935 133.305 205.025 ;
        RECT 133.475 203.935 133.755 205.075 ;
        RECT 133.925 204.105 134.255 205.085 ;
        RECT 134.425 203.935 134.685 205.075 ;
        RECT 134.860 203.935 135.180 205.075 ;
        RECT 135.360 204.195 135.555 205.245 ;
        RECT 135.915 205.065 136.085 205.445 ;
        RECT 135.735 204.785 136.085 205.065 ;
        RECT 136.275 204.915 136.520 205.275 ;
        RECT 138.280 205.110 138.620 205.940 ;
        RECT 142.215 205.715 143.885 206.485 ;
        RECT 144.055 205.745 144.545 206.315 ;
        RECT 144.715 205.915 144.945 206.315 ;
        RECT 145.115 206.085 145.535 206.485 ;
        RECT 145.705 205.915 145.875 206.315 ;
        RECT 144.715 205.745 145.875 205.915 ;
        RECT 146.045 205.745 146.495 206.485 ;
        RECT 146.665 205.745 147.105 206.305 ;
        RECT 147.275 205.940 152.620 206.485 ;
        RECT 135.735 204.105 136.065 204.785 ;
        RECT 136.265 203.935 136.520 204.735 ;
        RECT 140.100 204.370 140.450 205.620 ;
        RECT 142.215 205.195 142.965 205.715 ;
        RECT 143.135 205.025 143.885 205.545 ;
        RECT 136.695 203.935 142.040 204.370 ;
        RECT 142.215 203.935 143.885 205.025 ;
        RECT 144.055 205.075 144.225 205.745 ;
        RECT 144.395 205.245 144.800 205.575 ;
        RECT 144.055 204.905 144.825 205.075 ;
        RECT 144.065 203.935 144.395 204.735 ;
        RECT 144.575 204.275 144.825 204.905 ;
        RECT 145.015 204.445 145.265 205.575 ;
        RECT 145.465 205.245 145.710 205.575 ;
        RECT 145.895 205.295 146.285 205.575 ;
        RECT 145.465 204.445 145.665 205.245 ;
        RECT 146.455 205.125 146.625 205.575 ;
        RECT 145.835 204.955 146.625 205.125 ;
        RECT 145.835 204.275 146.005 204.955 ;
        RECT 144.575 204.105 146.005 204.275 ;
        RECT 146.175 203.935 146.490 204.785 ;
        RECT 146.795 204.735 147.105 205.745 ;
        RECT 148.860 205.110 149.200 205.940 ;
        RECT 152.795 205.715 156.305 206.485 ;
        RECT 156.935 205.735 158.145 206.485 ;
        RECT 146.665 204.105 147.105 204.735 ;
        RECT 150.680 204.370 151.030 205.620 ;
        RECT 152.795 205.195 154.445 205.715 ;
        RECT 154.615 205.025 156.305 205.545 ;
        RECT 147.275 203.935 152.620 204.370 ;
        RECT 152.795 203.935 156.305 205.025 ;
        RECT 156.935 205.025 157.455 205.565 ;
        RECT 157.625 205.195 158.145 205.735 ;
        RECT 156.935 203.935 158.145 205.025 ;
        RECT 2.750 203.765 158.230 203.935 ;
        RECT 2.835 202.675 4.045 203.765 ;
        RECT 5.140 203.095 5.395 203.595 ;
        RECT 5.565 203.265 5.895 203.765 ;
        RECT 5.140 202.925 5.890 203.095 ;
        RECT 2.835 201.965 3.355 202.505 ;
        RECT 3.525 202.135 4.045 202.675 ;
        RECT 5.140 202.105 5.490 202.755 ;
        RECT 2.835 201.215 4.045 201.965 ;
        RECT 5.660 201.935 5.890 202.925 ;
        RECT 5.140 201.765 5.890 201.935 ;
        RECT 5.140 201.475 5.395 201.765 ;
        RECT 5.565 201.215 5.895 201.595 ;
        RECT 6.065 201.475 6.235 203.595 ;
        RECT 6.405 202.795 6.730 203.580 ;
        RECT 6.900 203.305 7.150 203.765 ;
        RECT 7.320 203.265 7.570 203.595 ;
        RECT 7.785 203.265 8.465 203.595 ;
        RECT 7.320 203.135 7.490 203.265 ;
        RECT 7.095 202.965 7.490 203.135 ;
        RECT 6.465 201.745 6.925 202.795 ;
        RECT 7.095 201.605 7.265 202.965 ;
        RECT 7.660 202.705 8.125 203.095 ;
        RECT 7.435 201.895 7.785 202.515 ;
        RECT 7.955 202.115 8.125 202.705 ;
        RECT 8.295 202.485 8.465 203.265 ;
        RECT 8.635 203.165 8.805 203.505 ;
        RECT 9.040 203.335 9.370 203.765 ;
        RECT 9.540 203.165 9.710 203.505 ;
        RECT 10.005 203.305 10.375 203.765 ;
        RECT 8.635 202.995 9.710 203.165 ;
        RECT 10.545 203.135 10.715 203.595 ;
        RECT 10.950 203.255 11.820 203.595 ;
        RECT 11.990 203.305 12.240 203.765 ;
        RECT 10.155 202.965 10.715 203.135 ;
        RECT 10.155 202.825 10.325 202.965 ;
        RECT 8.825 202.655 10.325 202.825 ;
        RECT 11.020 202.795 11.480 203.085 ;
        RECT 8.295 202.315 9.985 202.485 ;
        RECT 7.955 201.895 8.310 202.115 ;
        RECT 8.480 201.605 8.650 202.315 ;
        RECT 8.855 201.895 9.645 202.145 ;
        RECT 9.815 202.135 9.985 202.315 ;
        RECT 10.155 201.965 10.325 202.655 ;
        RECT 6.595 201.215 6.925 201.575 ;
        RECT 7.095 201.435 7.590 201.605 ;
        RECT 7.795 201.435 8.650 201.605 ;
        RECT 9.525 201.215 9.855 201.675 ;
        RECT 10.065 201.575 10.325 201.965 ;
        RECT 10.515 202.785 11.480 202.795 ;
        RECT 11.650 202.875 11.820 203.255 ;
        RECT 12.410 203.215 12.580 203.505 ;
        RECT 12.760 203.385 13.090 203.765 ;
        RECT 12.410 203.045 13.210 203.215 ;
        RECT 10.515 202.625 11.190 202.785 ;
        RECT 11.650 202.705 12.870 202.875 ;
        RECT 10.515 201.835 10.725 202.625 ;
        RECT 11.650 202.615 11.820 202.705 ;
        RECT 10.895 201.835 11.245 202.455 ;
        RECT 11.415 202.445 11.820 202.615 ;
        RECT 11.415 201.665 11.585 202.445 ;
        RECT 11.755 201.995 11.975 202.275 ;
        RECT 12.155 202.165 12.695 202.535 ;
        RECT 13.040 202.455 13.210 203.045 ;
        RECT 13.430 202.625 13.735 203.765 ;
        RECT 13.905 202.575 14.160 203.455 ;
        RECT 13.040 202.425 13.780 202.455 ;
        RECT 11.755 201.825 12.285 201.995 ;
        RECT 10.065 201.405 10.415 201.575 ;
        RECT 10.635 201.385 11.585 201.665 ;
        RECT 11.755 201.215 11.945 201.655 ;
        RECT 12.115 201.595 12.285 201.825 ;
        RECT 12.455 201.765 12.695 202.165 ;
        RECT 12.865 202.125 13.780 202.425 ;
        RECT 12.865 201.950 13.190 202.125 ;
        RECT 12.865 201.595 13.185 201.950 ;
        RECT 13.950 201.925 14.160 202.575 ;
        RECT 12.115 201.425 13.185 201.595 ;
        RECT 13.430 201.215 13.735 201.675 ;
        RECT 13.905 201.395 14.160 201.925 ;
        RECT 14.335 202.690 14.605 203.595 ;
        RECT 14.775 203.005 15.105 203.765 ;
        RECT 15.285 202.835 15.455 203.595 ;
        RECT 14.335 201.890 14.505 202.690 ;
        RECT 14.790 202.665 15.455 202.835 ;
        RECT 14.790 202.520 14.960 202.665 ;
        RECT 15.715 202.600 16.005 203.765 ;
        RECT 16.175 202.915 16.555 203.595 ;
        RECT 17.145 202.915 17.315 203.765 ;
        RECT 17.485 203.085 17.815 203.595 ;
        RECT 17.985 203.255 18.155 203.765 ;
        RECT 18.325 203.085 18.725 203.595 ;
        RECT 17.485 202.915 18.725 203.085 ;
        RECT 14.675 202.190 14.960 202.520 ;
        RECT 14.790 201.935 14.960 202.190 ;
        RECT 15.195 202.115 15.525 202.485 ;
        RECT 16.175 201.955 16.345 202.915 ;
        RECT 16.515 202.575 17.820 202.745 ;
        RECT 18.905 202.665 19.225 203.595 ;
        RECT 16.515 202.125 16.760 202.575 ;
        RECT 16.930 202.205 17.480 202.405 ;
        RECT 17.650 202.375 17.820 202.575 ;
        RECT 18.595 202.495 19.225 202.665 ;
        RECT 19.405 203.155 19.735 203.585 ;
        RECT 19.915 203.325 20.110 203.765 ;
        RECT 20.280 203.155 20.610 203.585 ;
        RECT 19.405 202.985 20.610 203.155 ;
        RECT 19.405 202.655 20.300 202.985 ;
        RECT 20.780 202.815 21.055 203.585 ;
        RECT 20.470 202.625 21.055 202.815 ;
        RECT 21.420 202.795 21.810 202.970 ;
        RECT 22.295 202.965 22.625 203.765 ;
        RECT 22.795 202.975 23.330 203.595 ;
        RECT 21.420 202.625 22.845 202.795 ;
        RECT 17.650 202.205 18.025 202.375 ;
        RECT 18.195 201.955 18.425 202.455 ;
        RECT 14.335 201.385 14.595 201.890 ;
        RECT 14.790 201.765 15.455 201.935 ;
        RECT 14.775 201.215 15.105 201.595 ;
        RECT 15.285 201.385 15.455 201.765 ;
        RECT 15.715 201.215 16.005 201.940 ;
        RECT 16.175 201.785 18.425 201.955 ;
        RECT 16.225 201.215 16.555 201.605 ;
        RECT 16.725 201.465 16.895 201.785 ;
        RECT 18.595 201.615 18.765 202.495 ;
        RECT 19.410 202.125 19.705 202.455 ;
        RECT 19.885 202.125 20.300 202.455 ;
        RECT 17.065 201.215 17.395 201.605 ;
        RECT 17.810 201.445 18.765 201.615 ;
        RECT 18.935 201.215 19.225 202.050 ;
        RECT 19.405 201.215 19.705 201.945 ;
        RECT 19.885 201.505 20.115 202.125 ;
        RECT 20.470 201.955 20.645 202.625 ;
        RECT 20.315 201.775 20.645 201.955 ;
        RECT 20.815 201.805 21.055 202.455 ;
        RECT 21.295 201.895 21.650 202.455 ;
        RECT 20.315 201.395 20.540 201.775 ;
        RECT 21.820 201.725 21.990 202.625 ;
        RECT 22.160 201.895 22.425 202.455 ;
        RECT 22.675 202.125 22.845 202.625 ;
        RECT 23.015 201.955 23.330 202.975 ;
        RECT 24.455 203.005 24.970 203.415 ;
        RECT 25.205 203.005 25.375 203.765 ;
        RECT 25.545 203.425 27.575 203.595 ;
        RECT 24.455 202.195 24.795 203.005 ;
        RECT 25.545 202.760 25.715 203.425 ;
        RECT 26.110 203.085 27.235 203.255 ;
        RECT 24.965 202.570 25.715 202.760 ;
        RECT 25.885 202.745 26.895 202.915 ;
        RECT 24.455 202.025 25.685 202.195 ;
        RECT 20.710 201.215 21.040 201.605 ;
        RECT 21.400 201.215 21.640 201.725 ;
        RECT 21.820 201.395 22.100 201.725 ;
        RECT 22.330 201.215 22.545 201.725 ;
        RECT 22.715 201.385 23.330 201.955 ;
        RECT 24.730 201.420 24.975 202.025 ;
        RECT 25.195 201.215 25.705 201.750 ;
        RECT 25.885 201.385 26.075 202.745 ;
        RECT 26.245 201.725 26.520 202.545 ;
        RECT 26.725 201.945 26.895 202.745 ;
        RECT 27.065 201.955 27.235 203.085 ;
        RECT 27.405 202.455 27.575 203.425 ;
        RECT 27.745 202.625 27.915 203.765 ;
        RECT 28.085 202.625 28.420 203.595 ;
        RECT 28.605 202.815 28.880 203.585 ;
        RECT 29.050 203.155 29.380 203.585 ;
        RECT 29.550 203.325 29.745 203.765 ;
        RECT 29.925 203.155 30.255 203.585 ;
        RECT 29.050 202.985 30.255 203.155 ;
        RECT 28.605 202.625 29.190 202.815 ;
        RECT 29.360 202.655 30.255 202.985 ;
        RECT 30.900 203.095 31.155 203.595 ;
        RECT 31.325 203.265 31.655 203.765 ;
        RECT 30.900 202.925 31.650 203.095 ;
        RECT 27.405 202.125 27.600 202.455 ;
        RECT 27.825 202.125 28.080 202.455 ;
        RECT 27.825 201.955 27.995 202.125 ;
        RECT 28.250 201.955 28.420 202.625 ;
        RECT 27.065 201.785 27.995 201.955 ;
        RECT 27.065 201.750 27.240 201.785 ;
        RECT 26.245 201.555 26.525 201.725 ;
        RECT 26.245 201.385 26.520 201.555 ;
        RECT 26.710 201.385 27.240 201.750 ;
        RECT 27.665 201.215 27.995 201.615 ;
        RECT 28.165 201.385 28.420 201.955 ;
        RECT 28.605 201.805 28.845 202.455 ;
        RECT 29.015 201.955 29.190 202.625 ;
        RECT 29.360 202.125 29.775 202.455 ;
        RECT 29.955 202.125 30.250 202.455 ;
        RECT 29.015 201.775 29.345 201.955 ;
        RECT 28.620 201.215 28.950 201.605 ;
        RECT 29.120 201.395 29.345 201.775 ;
        RECT 29.545 201.505 29.775 202.125 ;
        RECT 30.900 202.105 31.250 202.755 ;
        RECT 29.955 201.215 30.255 201.945 ;
        RECT 31.420 201.935 31.650 202.925 ;
        RECT 30.900 201.765 31.650 201.935 ;
        RECT 30.900 201.475 31.155 201.765 ;
        RECT 31.325 201.215 31.655 201.595 ;
        RECT 31.825 201.475 31.995 203.595 ;
        RECT 32.165 202.795 32.490 203.580 ;
        RECT 32.660 203.305 32.910 203.765 ;
        RECT 33.080 203.265 33.330 203.595 ;
        RECT 33.545 203.265 34.225 203.595 ;
        RECT 33.080 203.135 33.250 203.265 ;
        RECT 32.855 202.965 33.250 203.135 ;
        RECT 32.225 201.745 32.685 202.795 ;
        RECT 32.855 201.605 33.025 202.965 ;
        RECT 33.420 202.705 33.885 203.095 ;
        RECT 33.195 201.895 33.545 202.515 ;
        RECT 33.715 202.115 33.885 202.705 ;
        RECT 34.055 202.485 34.225 203.265 ;
        RECT 34.395 203.165 34.565 203.505 ;
        RECT 34.800 203.335 35.130 203.765 ;
        RECT 35.300 203.165 35.470 203.505 ;
        RECT 35.765 203.305 36.135 203.765 ;
        RECT 34.395 202.995 35.470 203.165 ;
        RECT 36.305 203.135 36.475 203.595 ;
        RECT 36.710 203.255 37.580 203.595 ;
        RECT 37.750 203.305 38.000 203.765 ;
        RECT 35.915 202.965 36.475 203.135 ;
        RECT 35.915 202.825 36.085 202.965 ;
        RECT 34.585 202.655 36.085 202.825 ;
        RECT 36.780 202.795 37.240 203.085 ;
        RECT 34.055 202.315 35.745 202.485 ;
        RECT 33.715 201.895 34.070 202.115 ;
        RECT 34.240 201.605 34.410 202.315 ;
        RECT 34.615 201.895 35.405 202.145 ;
        RECT 35.575 202.135 35.745 202.315 ;
        RECT 35.915 201.965 36.085 202.655 ;
        RECT 32.355 201.215 32.685 201.575 ;
        RECT 32.855 201.435 33.350 201.605 ;
        RECT 33.555 201.435 34.410 201.605 ;
        RECT 35.285 201.215 35.615 201.675 ;
        RECT 35.825 201.575 36.085 201.965 ;
        RECT 36.275 202.785 37.240 202.795 ;
        RECT 37.410 202.875 37.580 203.255 ;
        RECT 38.170 203.215 38.340 203.505 ;
        RECT 38.520 203.385 38.850 203.765 ;
        RECT 38.170 203.045 38.970 203.215 ;
        RECT 36.275 202.625 36.950 202.785 ;
        RECT 37.410 202.705 38.630 202.875 ;
        RECT 36.275 201.835 36.485 202.625 ;
        RECT 37.410 202.615 37.580 202.705 ;
        RECT 36.655 201.835 37.005 202.455 ;
        RECT 37.175 202.445 37.580 202.615 ;
        RECT 37.175 201.665 37.345 202.445 ;
        RECT 37.515 201.995 37.735 202.275 ;
        RECT 37.915 202.165 38.455 202.535 ;
        RECT 38.800 202.455 38.970 203.045 ;
        RECT 39.190 202.625 39.495 203.765 ;
        RECT 39.665 202.575 39.920 203.455 ;
        RECT 40.105 202.625 40.435 203.765 ;
        RECT 40.965 202.795 41.295 203.580 ;
        RECT 40.615 202.625 41.295 202.795 ;
        RECT 38.800 202.425 39.540 202.455 ;
        RECT 37.515 201.825 38.045 201.995 ;
        RECT 35.825 201.405 36.175 201.575 ;
        RECT 36.395 201.385 37.345 201.665 ;
        RECT 37.515 201.215 37.705 201.655 ;
        RECT 37.875 201.595 38.045 201.825 ;
        RECT 38.215 201.765 38.455 202.165 ;
        RECT 38.625 202.125 39.540 202.425 ;
        RECT 38.625 201.950 38.950 202.125 ;
        RECT 38.625 201.595 38.945 201.950 ;
        RECT 39.710 201.925 39.920 202.575 ;
        RECT 40.095 202.205 40.445 202.455 ;
        RECT 40.615 202.025 40.785 202.625 ;
        RECT 41.475 202.600 41.765 203.765 ;
        RECT 42.860 203.095 43.115 203.595 ;
        RECT 43.285 203.265 43.615 203.765 ;
        RECT 42.860 202.925 43.610 203.095 ;
        RECT 40.955 202.205 41.305 202.455 ;
        RECT 42.860 202.105 43.210 202.755 ;
        RECT 37.875 201.425 38.945 201.595 ;
        RECT 39.190 201.215 39.495 201.675 ;
        RECT 39.665 201.395 39.920 201.925 ;
        RECT 40.105 201.215 40.375 202.025 ;
        RECT 40.545 201.385 40.875 202.025 ;
        RECT 41.045 201.215 41.285 202.025 ;
        RECT 41.475 201.215 41.765 201.940 ;
        RECT 43.380 201.935 43.610 202.925 ;
        RECT 42.860 201.765 43.610 201.935 ;
        RECT 42.860 201.475 43.115 201.765 ;
        RECT 43.285 201.215 43.615 201.595 ;
        RECT 43.785 201.475 43.955 203.595 ;
        RECT 44.125 202.795 44.450 203.580 ;
        RECT 44.620 203.305 44.870 203.765 ;
        RECT 45.040 203.265 45.290 203.595 ;
        RECT 45.505 203.265 46.185 203.595 ;
        RECT 45.040 203.135 45.210 203.265 ;
        RECT 44.815 202.965 45.210 203.135 ;
        RECT 44.185 201.745 44.645 202.795 ;
        RECT 44.815 201.605 44.985 202.965 ;
        RECT 45.380 202.705 45.845 203.095 ;
        RECT 45.155 201.895 45.505 202.515 ;
        RECT 45.675 202.115 45.845 202.705 ;
        RECT 46.015 202.485 46.185 203.265 ;
        RECT 46.355 203.165 46.525 203.505 ;
        RECT 46.760 203.335 47.090 203.765 ;
        RECT 47.260 203.165 47.430 203.505 ;
        RECT 47.725 203.305 48.095 203.765 ;
        RECT 46.355 202.995 47.430 203.165 ;
        RECT 48.265 203.135 48.435 203.595 ;
        RECT 48.670 203.255 49.540 203.595 ;
        RECT 49.710 203.305 49.960 203.765 ;
        RECT 47.875 202.965 48.435 203.135 ;
        RECT 47.875 202.825 48.045 202.965 ;
        RECT 46.545 202.655 48.045 202.825 ;
        RECT 48.740 202.795 49.200 203.085 ;
        RECT 46.015 202.315 47.705 202.485 ;
        RECT 45.675 201.895 46.030 202.115 ;
        RECT 46.200 201.605 46.370 202.315 ;
        RECT 46.575 201.895 47.365 202.145 ;
        RECT 47.535 202.135 47.705 202.315 ;
        RECT 47.875 201.965 48.045 202.655 ;
        RECT 44.315 201.215 44.645 201.575 ;
        RECT 44.815 201.435 45.310 201.605 ;
        RECT 45.515 201.435 46.370 201.605 ;
        RECT 47.245 201.215 47.575 201.675 ;
        RECT 47.785 201.575 48.045 201.965 ;
        RECT 48.235 202.785 49.200 202.795 ;
        RECT 49.370 202.875 49.540 203.255 ;
        RECT 50.130 203.215 50.300 203.505 ;
        RECT 50.480 203.385 50.810 203.765 ;
        RECT 50.130 203.045 50.930 203.215 ;
        RECT 48.235 202.625 48.910 202.785 ;
        RECT 49.370 202.705 50.590 202.875 ;
        RECT 48.235 201.835 48.445 202.625 ;
        RECT 49.370 202.615 49.540 202.705 ;
        RECT 48.615 201.835 48.965 202.455 ;
        RECT 49.135 202.445 49.540 202.615 ;
        RECT 49.135 201.665 49.305 202.445 ;
        RECT 49.475 201.995 49.695 202.275 ;
        RECT 49.875 202.165 50.415 202.535 ;
        RECT 50.760 202.455 50.930 203.045 ;
        RECT 51.150 202.625 51.455 203.765 ;
        RECT 51.625 202.575 51.880 203.455 ;
        RECT 50.760 202.425 51.500 202.455 ;
        RECT 49.475 201.825 50.005 201.995 ;
        RECT 47.785 201.405 48.135 201.575 ;
        RECT 48.355 201.385 49.305 201.665 ;
        RECT 49.475 201.215 49.665 201.655 ;
        RECT 49.835 201.595 50.005 201.825 ;
        RECT 50.175 201.765 50.415 202.165 ;
        RECT 50.585 202.125 51.500 202.425 ;
        RECT 50.585 201.950 50.910 202.125 ;
        RECT 50.585 201.595 50.905 201.950 ;
        RECT 51.670 201.925 51.880 202.575 ;
        RECT 49.835 201.425 50.905 201.595 ;
        RECT 51.150 201.215 51.455 201.675 ;
        RECT 51.625 201.395 51.880 201.925 ;
        RECT 52.065 201.395 52.325 203.585 ;
        RECT 52.495 203.035 52.835 203.765 ;
        RECT 53.015 202.855 53.285 203.585 ;
        RECT 52.515 202.635 53.285 202.855 ;
        RECT 53.465 202.875 53.695 203.585 ;
        RECT 53.865 203.055 54.195 203.765 ;
        RECT 54.365 202.875 54.625 203.585 ;
        RECT 53.465 202.635 54.625 202.875 ;
        RECT 54.815 202.690 55.085 203.595 ;
        RECT 55.255 203.005 55.585 203.765 ;
        RECT 55.765 202.835 55.935 203.595 ;
        RECT 52.515 201.965 52.805 202.635 ;
        RECT 52.985 202.145 53.450 202.455 ;
        RECT 53.630 202.145 54.155 202.455 ;
        RECT 52.515 201.765 53.745 201.965 ;
        RECT 52.585 201.215 53.255 201.585 ;
        RECT 53.435 201.395 53.745 201.765 ;
        RECT 53.925 201.505 54.155 202.145 ;
        RECT 54.335 202.125 54.635 202.455 ;
        RECT 54.335 201.215 54.625 201.945 ;
        RECT 54.815 201.890 54.985 202.690 ;
        RECT 55.270 202.665 55.935 202.835 ;
        RECT 55.270 202.520 55.440 202.665 ;
        RECT 55.155 202.190 55.440 202.520 ;
        RECT 55.270 201.935 55.440 202.190 ;
        RECT 55.675 202.115 56.005 202.485 ;
        RECT 56.195 202.160 56.475 203.595 ;
        RECT 56.645 202.990 57.355 203.765 ;
        RECT 57.525 202.820 57.855 203.595 ;
        RECT 56.705 202.605 57.855 202.820 ;
        RECT 54.815 201.385 55.075 201.890 ;
        RECT 55.270 201.765 55.935 201.935 ;
        RECT 55.255 201.215 55.585 201.595 ;
        RECT 55.765 201.385 55.935 201.765 ;
        RECT 56.195 201.385 56.535 202.160 ;
        RECT 56.705 202.035 56.990 202.605 ;
        RECT 57.175 202.205 57.645 202.435 ;
        RECT 58.050 202.405 58.265 203.520 ;
        RECT 58.445 203.045 58.775 203.765 ;
        RECT 58.555 202.405 58.785 202.745 ;
        RECT 57.815 202.225 58.265 202.405 ;
        RECT 57.815 202.205 58.145 202.225 ;
        RECT 58.455 202.205 58.785 202.405 ;
        RECT 58.955 202.160 59.235 203.595 ;
        RECT 59.405 202.990 60.115 203.765 ;
        RECT 60.285 202.820 60.615 203.595 ;
        RECT 59.465 202.605 60.615 202.820 ;
        RECT 56.705 201.845 57.415 202.035 ;
        RECT 57.115 201.705 57.415 201.845 ;
        RECT 57.605 201.845 58.785 202.035 ;
        RECT 57.605 201.765 57.935 201.845 ;
        RECT 57.115 201.695 57.430 201.705 ;
        RECT 57.115 201.685 57.440 201.695 ;
        RECT 57.115 201.680 57.450 201.685 ;
        RECT 56.705 201.215 56.875 201.675 ;
        RECT 57.115 201.670 57.455 201.680 ;
        RECT 57.115 201.665 57.460 201.670 ;
        RECT 57.115 201.655 57.465 201.665 ;
        RECT 57.115 201.650 57.470 201.655 ;
        RECT 57.115 201.385 57.475 201.650 ;
        RECT 58.105 201.215 58.275 201.675 ;
        RECT 58.445 201.385 58.785 201.845 ;
        RECT 58.955 201.385 59.295 202.160 ;
        RECT 59.465 202.035 59.750 202.605 ;
        RECT 59.935 202.205 60.405 202.435 ;
        RECT 60.810 202.405 61.025 203.520 ;
        RECT 61.205 203.045 61.535 203.765 ;
        RECT 62.725 203.095 62.895 203.595 ;
        RECT 63.135 203.305 63.385 203.765 ;
        RECT 63.685 203.095 63.855 203.595 ;
        RECT 64.065 203.305 64.315 203.765 ;
        RECT 64.525 203.095 64.695 203.595 ;
        RECT 62.725 202.925 64.695 203.095 ;
        RECT 64.865 203.125 65.195 203.555 ;
        RECT 65.385 203.305 65.635 203.765 ;
        RECT 65.805 203.295 66.145 203.555 ;
        RECT 64.865 202.955 65.715 203.125 ;
        RECT 61.315 202.405 61.545 202.745 ;
        RECT 60.575 202.225 61.025 202.405 ;
        RECT 60.575 202.205 60.905 202.225 ;
        RECT 61.215 202.205 61.545 202.405 ;
        RECT 62.660 202.125 62.915 202.755 ;
        RECT 63.145 202.125 63.525 202.755 ;
        RECT 64.395 202.455 64.695 202.750 ;
        RECT 59.465 201.845 60.175 202.035 ;
        RECT 59.875 201.705 60.175 201.845 ;
        RECT 60.365 201.845 61.545 202.035 ;
        RECT 60.365 201.765 60.695 201.845 ;
        RECT 59.875 201.695 60.190 201.705 ;
        RECT 59.875 201.685 60.200 201.695 ;
        RECT 59.875 201.680 60.210 201.685 ;
        RECT 59.465 201.215 59.635 201.675 ;
        RECT 59.875 201.670 60.215 201.680 ;
        RECT 59.875 201.665 60.220 201.670 ;
        RECT 59.875 201.655 60.225 201.665 ;
        RECT 59.875 201.650 60.230 201.655 ;
        RECT 59.875 201.385 60.235 201.650 ;
        RECT 60.865 201.215 61.035 201.675 ;
        RECT 61.205 201.385 61.545 201.845 ;
        RECT 62.635 201.215 62.975 201.940 ;
        RECT 63.145 201.525 63.350 202.125 ;
        RECT 63.785 201.730 64.005 202.455 ;
        RECT 64.315 202.405 64.695 202.455 ;
        RECT 64.315 202.235 64.705 202.405 ;
        RECT 64.315 202.125 64.695 202.235 ;
        RECT 64.895 202.205 65.225 202.765 ;
        RECT 65.545 202.035 65.715 202.955 ;
        RECT 64.895 201.940 65.715 202.035 ;
        RECT 64.700 201.865 65.715 201.940 ;
        RECT 63.580 201.545 64.530 201.730 ;
        RECT 64.700 201.430 65.115 201.865 ;
        RECT 65.305 201.215 65.635 201.695 ;
        RECT 65.885 201.690 66.145 203.295 ;
        RECT 67.235 202.600 67.525 203.765 ;
        RECT 67.695 202.675 68.905 203.765 ;
        RECT 69.085 202.965 69.415 203.765 ;
        RECT 69.595 203.425 71.025 203.595 ;
        RECT 69.595 202.795 69.845 203.425 ;
        RECT 67.695 201.965 68.215 202.505 ;
        RECT 68.385 202.135 68.905 202.675 ;
        RECT 69.075 202.625 69.845 202.795 ;
        RECT 65.805 201.430 66.145 201.690 ;
        RECT 67.235 201.215 67.525 201.940 ;
        RECT 67.695 201.215 68.905 201.965 ;
        RECT 69.075 201.955 69.245 202.625 ;
        RECT 69.415 202.125 69.820 202.455 ;
        RECT 70.035 202.125 70.285 203.255 ;
        RECT 70.485 202.455 70.685 203.255 ;
        RECT 70.855 202.745 71.025 203.425 ;
        RECT 71.195 202.915 71.510 203.765 ;
        RECT 71.685 202.965 72.125 203.595 ;
        RECT 70.855 202.575 71.645 202.745 ;
        RECT 70.485 202.125 70.730 202.455 ;
        RECT 70.915 202.125 71.305 202.405 ;
        RECT 71.475 202.125 71.645 202.575 ;
        RECT 71.815 201.955 72.125 202.965 ;
        RECT 69.075 201.385 69.565 201.955 ;
        RECT 69.735 201.785 70.895 201.955 ;
        RECT 69.735 201.385 69.965 201.785 ;
        RECT 70.135 201.215 70.555 201.615 ;
        RECT 70.725 201.385 70.895 201.785 ;
        RECT 71.065 201.215 71.515 201.955 ;
        RECT 71.685 201.395 72.125 201.955 ;
        RECT 72.295 202.965 72.735 203.595 ;
        RECT 72.295 201.955 72.605 202.965 ;
        RECT 72.910 202.915 73.225 203.765 ;
        RECT 73.395 203.425 74.825 203.595 ;
        RECT 73.395 202.745 73.565 203.425 ;
        RECT 72.775 202.575 73.565 202.745 ;
        RECT 72.775 202.125 72.945 202.575 ;
        RECT 73.735 202.455 73.935 203.255 ;
        RECT 73.115 202.125 73.505 202.405 ;
        RECT 73.690 202.125 73.935 202.455 ;
        RECT 74.135 202.125 74.385 203.255 ;
        RECT 74.575 202.795 74.825 203.425 ;
        RECT 75.005 202.965 75.335 203.765 ;
        RECT 76.180 202.795 76.510 203.595 ;
        RECT 76.680 202.965 77.010 203.765 ;
        RECT 77.310 202.795 77.640 203.595 ;
        RECT 78.285 202.965 78.535 203.765 ;
        RECT 74.575 202.625 75.345 202.795 ;
        RECT 76.180 202.625 78.615 202.795 ;
        RECT 78.805 202.625 78.975 203.765 ;
        RECT 79.145 202.625 79.485 203.595 ;
        RECT 79.660 203.410 80.740 203.580 ;
        RECT 79.660 202.625 79.995 203.410 ;
        RECT 74.600 202.125 75.005 202.455 ;
        RECT 75.175 201.955 75.345 202.625 ;
        RECT 75.975 202.205 76.325 202.455 ;
        RECT 76.510 201.995 76.680 202.625 ;
        RECT 76.850 202.205 77.180 202.405 ;
        RECT 77.350 202.205 77.680 202.405 ;
        RECT 77.850 202.205 78.270 202.405 ;
        RECT 78.445 202.375 78.615 202.625 ;
        RECT 79.255 202.575 79.485 202.625 ;
        RECT 78.445 202.205 79.140 202.375 ;
        RECT 72.295 201.395 72.735 201.955 ;
        RECT 72.905 201.215 73.355 201.955 ;
        RECT 73.525 201.785 74.685 201.955 ;
        RECT 73.525 201.385 73.695 201.785 ;
        RECT 73.865 201.215 74.285 201.615 ;
        RECT 74.455 201.385 74.685 201.785 ;
        RECT 74.855 201.385 75.345 201.955 ;
        RECT 76.180 201.385 76.680 201.995 ;
        RECT 77.310 201.865 78.535 202.035 ;
        RECT 79.310 202.015 79.485 202.575 ;
        RECT 80.165 202.455 80.400 203.135 ;
        RECT 80.570 202.795 80.740 203.410 ;
        RECT 81.005 202.965 81.320 203.765 ;
        RECT 80.570 202.625 80.885 202.795 ;
        RECT 79.660 202.125 79.995 202.455 ;
        RECT 80.165 202.125 80.545 202.455 ;
        RECT 77.310 201.385 77.640 201.865 ;
        RECT 77.810 201.215 78.035 201.675 ;
        RECT 78.205 201.385 78.535 201.865 ;
        RECT 78.725 201.215 78.975 202.015 ;
        RECT 79.145 201.385 79.485 202.015 ;
        RECT 80.715 201.955 80.885 202.625 ;
        RECT 79.660 201.785 80.885 201.955 ;
        RECT 81.055 201.785 81.325 202.795 ;
        RECT 81.495 202.675 84.085 203.765 ;
        RECT 81.495 201.985 82.705 202.505 ;
        RECT 82.875 202.155 84.085 202.675 ;
        RECT 84.255 202.625 84.515 203.765 ;
        RECT 84.755 203.255 86.370 203.585 ;
        RECT 84.765 202.455 84.935 203.015 ;
        RECT 85.195 202.915 86.370 203.085 ;
        RECT 86.540 202.965 86.820 203.765 ;
        RECT 85.195 202.625 85.525 202.915 ;
        RECT 86.200 202.795 86.370 202.915 ;
        RECT 85.695 202.455 85.940 202.745 ;
        RECT 86.200 202.625 86.860 202.795 ;
        RECT 87.030 202.625 87.305 203.595 ;
        RECT 87.475 203.330 92.820 203.765 ;
        RECT 86.690 202.455 86.860 202.625 ;
        RECT 84.260 202.205 84.595 202.455 ;
        RECT 84.765 202.125 85.480 202.455 ;
        RECT 85.695 202.125 86.520 202.455 ;
        RECT 86.690 202.125 86.965 202.455 ;
        RECT 84.765 202.035 85.015 202.125 ;
        RECT 79.660 201.515 79.915 201.785 ;
        RECT 80.085 201.215 80.415 201.615 ;
        RECT 80.585 201.515 80.755 201.785 ;
        RECT 80.925 201.215 81.255 201.615 ;
        RECT 81.495 201.215 84.085 201.985 ;
        RECT 84.255 201.215 84.515 202.035 ;
        RECT 84.685 201.615 85.015 202.035 ;
        RECT 86.690 201.955 86.860 202.125 ;
        RECT 85.195 201.785 86.860 201.955 ;
        RECT 87.135 201.890 87.305 202.625 ;
        RECT 85.195 201.385 85.455 201.785 ;
        RECT 85.625 201.215 85.955 201.615 ;
        RECT 86.125 201.435 86.295 201.785 ;
        RECT 86.465 201.215 86.840 201.615 ;
        RECT 87.030 201.545 87.305 201.890 ;
        RECT 89.060 201.760 89.400 202.590 ;
        RECT 90.880 202.080 91.230 203.330 ;
        RECT 92.995 202.600 93.285 203.765 ;
        RECT 93.955 202.815 94.245 203.585 ;
        RECT 94.815 203.225 95.075 203.585 ;
        RECT 95.245 203.395 95.575 203.765 ;
        RECT 95.745 203.225 96.005 203.585 ;
        RECT 94.815 202.995 96.005 203.225 ;
        RECT 96.195 203.045 96.525 203.765 ;
        RECT 96.695 202.815 96.960 203.585 ;
        RECT 97.140 202.965 97.395 203.765 ;
        RECT 97.595 202.915 97.925 203.595 ;
        RECT 93.955 202.635 96.450 202.815 ;
        RECT 93.925 202.125 94.195 202.455 ;
        RECT 94.375 202.125 94.810 202.455 ;
        RECT 94.990 202.125 95.565 202.455 ;
        RECT 95.745 202.125 96.025 202.455 ;
        RECT 96.225 201.945 96.450 202.635 ;
        RECT 87.475 201.215 92.820 201.760 ;
        RECT 92.995 201.215 93.285 201.940 ;
        RECT 93.965 201.755 96.450 201.945 ;
        RECT 93.965 201.395 94.190 201.755 ;
        RECT 94.370 201.215 94.700 201.585 ;
        RECT 94.880 201.395 95.135 201.755 ;
        RECT 95.700 201.215 96.445 201.585 ;
        RECT 96.625 201.395 96.960 202.815 ;
        RECT 97.140 202.425 97.385 202.785 ;
        RECT 97.575 202.635 97.925 202.915 ;
        RECT 97.575 202.255 97.745 202.635 ;
        RECT 98.105 202.455 98.300 203.505 ;
        RECT 98.480 202.625 98.800 203.765 ;
        RECT 98.975 202.675 101.565 203.765 ;
        RECT 101.740 203.255 103.395 203.545 ;
        RECT 97.225 202.085 97.745 202.255 ;
        RECT 97.915 202.125 98.300 202.455 ;
        RECT 98.480 202.405 98.740 202.455 ;
        RECT 98.480 202.235 98.745 202.405 ;
        RECT 98.480 202.125 98.740 202.235 ;
        RECT 97.225 201.520 97.395 202.085 ;
        RECT 98.975 201.985 100.185 202.505 ;
        RECT 100.355 202.155 101.565 202.675 ;
        RECT 101.740 202.915 103.330 203.085 ;
        RECT 103.565 202.965 103.845 203.765 ;
        RECT 101.740 202.625 102.060 202.915 ;
        RECT 103.160 202.795 103.330 202.915 ;
        RECT 102.255 202.575 102.970 202.745 ;
        RECT 103.160 202.625 103.885 202.795 ;
        RECT 104.055 202.625 104.325 203.595 ;
        RECT 104.495 203.330 109.840 203.765 ;
        RECT 97.585 201.745 98.800 201.915 ;
        RECT 97.585 201.440 97.815 201.745 ;
        RECT 97.985 201.215 98.315 201.575 ;
        RECT 98.510 201.395 98.800 201.745 ;
        RECT 98.975 201.215 101.565 201.985 ;
        RECT 101.740 201.885 102.090 202.455 ;
        RECT 102.260 202.125 102.970 202.575 ;
        RECT 103.715 202.455 103.885 202.625 ;
        RECT 103.140 202.125 103.545 202.455 ;
        RECT 103.715 202.125 103.985 202.455 ;
        RECT 103.715 201.955 103.885 202.125 ;
        RECT 102.275 201.785 103.885 201.955 ;
        RECT 104.155 201.890 104.325 202.625 ;
        RECT 101.745 201.215 102.075 201.715 ;
        RECT 102.275 201.435 102.445 201.785 ;
        RECT 102.645 201.215 102.975 201.615 ;
        RECT 103.145 201.435 103.315 201.785 ;
        RECT 103.485 201.215 103.865 201.615 ;
        RECT 104.055 201.545 104.325 201.890 ;
        RECT 106.080 201.760 106.420 202.590 ;
        RECT 107.900 202.080 108.250 203.330 ;
        RECT 110.015 202.675 112.605 203.765 ;
        RECT 110.015 201.985 111.225 202.505 ;
        RECT 111.395 202.155 112.605 202.675 ;
        RECT 113.235 202.585 113.555 203.765 ;
        RECT 113.725 202.745 113.925 203.535 ;
        RECT 114.250 202.935 114.635 203.595 ;
        RECT 115.030 203.005 115.815 203.765 ;
        RECT 114.225 202.835 114.635 202.935 ;
        RECT 113.725 202.575 114.055 202.745 ;
        RECT 114.225 202.625 115.835 202.835 ;
        RECT 113.875 202.455 114.055 202.575 ;
        RECT 113.235 202.205 113.700 202.405 ;
        RECT 113.875 202.205 114.205 202.455 ;
        RECT 114.375 202.405 114.840 202.455 ;
        RECT 114.375 202.235 114.845 202.405 ;
        RECT 114.375 202.205 114.840 202.235 ;
        RECT 115.035 202.205 115.390 202.455 ;
        RECT 115.560 202.025 115.835 202.625 ;
        RECT 104.495 201.215 109.840 201.760 ;
        RECT 110.015 201.215 112.605 201.985 ;
        RECT 113.235 201.825 114.415 201.995 ;
        RECT 113.235 201.410 113.575 201.825 ;
        RECT 113.745 201.215 113.915 201.655 ;
        RECT 114.085 201.605 114.415 201.825 ;
        RECT 114.585 201.845 115.835 202.025 ;
        RECT 114.585 201.775 114.950 201.845 ;
        RECT 114.085 201.425 115.335 201.605 ;
        RECT 115.605 201.215 115.775 201.675 ;
        RECT 116.005 201.495 116.285 203.595 ;
        RECT 116.455 202.675 118.125 203.765 ;
        RECT 116.455 201.985 117.205 202.505 ;
        RECT 117.375 202.155 118.125 202.675 ;
        RECT 118.755 202.600 119.045 203.765 ;
        RECT 119.675 202.965 120.000 203.765 ;
        RECT 119.695 202.205 120.025 202.790 ;
        RECT 120.195 202.455 120.380 203.545 ;
        RECT 120.550 202.795 120.800 203.595 ;
        RECT 120.970 202.965 121.710 203.765 ;
        RECT 121.895 202.795 122.225 203.595 ;
        RECT 122.395 202.965 123.205 203.765 ;
        RECT 120.550 202.625 123.035 202.795 ;
        RECT 122.865 202.455 123.035 202.625 ;
        RECT 120.195 202.205 120.680 202.455 ;
        RECT 121.025 202.125 121.285 202.455 ;
        RECT 116.455 201.215 118.125 201.985 ;
        RECT 118.755 201.215 119.045 201.940 ;
        RECT 119.675 201.835 120.860 202.005 ;
        RECT 119.675 201.385 119.940 201.835 ;
        RECT 120.110 201.215 120.400 201.665 ;
        RECT 120.570 201.385 120.860 201.835 ;
        RECT 121.040 201.520 121.285 202.125 ;
        RECT 121.535 201.520 121.805 202.455 ;
        RECT 121.985 202.205 122.465 202.455 ;
        RECT 121.985 201.520 122.195 202.205 ;
        RECT 122.865 202.125 123.205 202.455 ;
        RECT 122.865 202.035 123.035 202.125 ;
        RECT 122.365 201.865 123.035 202.035 ;
        RECT 122.365 201.385 122.705 201.865 ;
        RECT 122.885 201.215 123.195 201.695 ;
        RECT 123.375 201.385 123.635 203.595 ;
        RECT 123.815 202.625 124.085 203.595 ;
        RECT 124.295 202.965 124.575 203.765 ;
        RECT 124.745 203.255 126.400 203.545 ;
        RECT 124.810 202.915 126.400 203.085 ;
        RECT 124.810 202.795 124.980 202.915 ;
        RECT 124.255 202.625 124.980 202.795 ;
        RECT 123.815 201.890 123.985 202.625 ;
        RECT 124.255 202.455 124.425 202.625 ;
        RECT 124.155 202.125 124.425 202.455 ;
        RECT 124.595 202.125 125.000 202.455 ;
        RECT 125.170 202.125 125.880 202.745 ;
        RECT 126.080 202.625 126.400 202.915 ;
        RECT 126.575 202.675 130.085 203.765 ;
        RECT 124.255 201.955 124.425 202.125 ;
        RECT 123.815 201.545 124.085 201.890 ;
        RECT 124.255 201.785 125.865 201.955 ;
        RECT 126.050 201.885 126.400 202.455 ;
        RECT 126.575 201.985 128.225 202.505 ;
        RECT 128.395 202.155 130.085 202.675 ;
        RECT 130.720 202.625 130.975 203.765 ;
        RECT 131.145 202.725 131.455 203.595 ;
        RECT 131.655 203.305 131.945 203.765 ;
        RECT 132.115 203.385 133.425 203.555 ;
        RECT 132.115 203.135 132.285 203.385 ;
        RECT 133.955 203.305 134.175 203.765 ;
        RECT 134.345 203.135 134.680 203.595 ;
        RECT 131.625 202.965 132.285 203.135 ;
        RECT 132.455 202.965 134.680 203.135 ;
        RECT 124.275 201.215 124.655 201.615 ;
        RECT 124.825 201.435 124.995 201.785 ;
        RECT 125.165 201.215 125.495 201.615 ;
        RECT 125.695 201.435 125.865 201.785 ;
        RECT 126.065 201.215 126.395 201.715 ;
        RECT 126.575 201.215 130.085 201.985 ;
        RECT 130.720 201.215 130.975 202.015 ;
        RECT 131.145 201.880 131.315 202.725 ;
        RECT 131.625 202.455 131.795 202.965 ;
        RECT 132.455 202.795 132.625 202.965 ;
        RECT 131.485 202.125 131.795 202.455 ;
        RECT 131.965 202.625 132.625 202.795 ;
        RECT 131.965 202.125 132.135 202.625 ;
        RECT 132.905 202.445 133.720 202.755 ;
        RECT 132.905 202.410 133.075 202.445 ;
        RECT 131.625 201.935 131.795 202.125 ;
        RECT 131.145 201.385 131.395 201.880 ;
        RECT 131.625 201.765 132.235 201.935 ;
        RECT 132.445 201.895 133.075 202.410 ;
        RECT 133.255 201.865 133.720 202.155 ;
        RECT 133.990 201.885 134.180 202.755 ;
        RECT 132.065 201.595 132.235 201.765 ;
        RECT 131.565 201.215 131.895 201.595 ;
        RECT 132.065 201.425 133.360 201.595 ;
        RECT 133.530 201.550 133.720 201.865 ;
        RECT 133.980 201.215 134.180 201.715 ;
        RECT 134.350 201.385 134.680 202.965 ;
        RECT 134.855 202.675 136.525 203.765 ;
        RECT 134.855 201.985 135.605 202.505 ;
        RECT 135.775 202.155 136.525 202.675 ;
        RECT 136.695 202.895 136.970 203.595 ;
        RECT 137.140 203.220 137.395 203.765 ;
        RECT 137.565 203.255 138.045 203.595 ;
        RECT 138.220 203.210 138.825 203.765 ;
        RECT 138.995 203.330 144.340 203.765 ;
        RECT 138.210 203.110 138.825 203.210 ;
        RECT 138.210 203.085 138.395 203.110 ;
        RECT 134.855 201.215 136.525 201.985 ;
        RECT 136.695 201.865 136.865 202.895 ;
        RECT 137.140 202.765 137.895 203.015 ;
        RECT 138.065 202.840 138.395 203.085 ;
        RECT 137.140 202.730 137.910 202.765 ;
        RECT 137.140 202.720 137.925 202.730 ;
        RECT 137.035 202.705 137.930 202.720 ;
        RECT 137.035 202.690 137.950 202.705 ;
        RECT 137.035 202.680 137.970 202.690 ;
        RECT 137.035 202.670 137.995 202.680 ;
        RECT 137.035 202.640 138.065 202.670 ;
        RECT 137.035 202.610 138.085 202.640 ;
        RECT 137.035 202.580 138.105 202.610 ;
        RECT 137.035 202.555 138.135 202.580 ;
        RECT 137.035 202.520 138.170 202.555 ;
        RECT 137.035 202.515 138.200 202.520 ;
        RECT 137.035 202.120 137.265 202.515 ;
        RECT 137.810 202.510 138.200 202.515 ;
        RECT 137.835 202.500 138.200 202.510 ;
        RECT 137.850 202.495 138.200 202.500 ;
        RECT 137.865 202.490 138.200 202.495 ;
        RECT 138.565 202.490 138.825 202.940 ;
        RECT 137.865 202.485 138.825 202.490 ;
        RECT 137.875 202.475 138.825 202.485 ;
        RECT 137.885 202.470 138.825 202.475 ;
        RECT 137.895 202.460 138.825 202.470 ;
        RECT 137.900 202.450 138.825 202.460 ;
        RECT 137.905 202.445 138.825 202.450 ;
        RECT 137.915 202.430 138.825 202.445 ;
        RECT 137.920 202.415 138.825 202.430 ;
        RECT 137.930 202.390 138.825 202.415 ;
        RECT 137.435 201.920 137.765 202.345 ;
        RECT 136.695 201.385 136.955 201.865 ;
        RECT 137.125 201.215 137.375 201.755 ;
        RECT 137.545 201.435 137.765 201.920 ;
        RECT 137.935 202.320 138.825 202.390 ;
        RECT 137.935 201.595 138.105 202.320 ;
        RECT 138.275 201.765 138.825 202.150 ;
        RECT 140.580 201.760 140.920 202.590 ;
        RECT 142.400 202.080 142.750 203.330 ;
        RECT 144.515 202.600 144.805 203.765 ;
        RECT 144.975 202.795 145.285 203.595 ;
        RECT 145.455 202.965 145.765 203.765 ;
        RECT 145.935 203.135 146.195 203.595 ;
        RECT 146.365 203.305 146.620 203.765 ;
        RECT 146.795 203.135 147.055 203.595 ;
        RECT 145.935 202.965 147.055 203.135 ;
        RECT 144.975 202.625 146.005 202.795 ;
        RECT 137.935 201.425 138.825 201.595 ;
        RECT 138.995 201.215 144.340 201.760 ;
        RECT 144.515 201.215 144.805 201.940 ;
        RECT 144.975 201.715 145.145 202.625 ;
        RECT 145.315 201.885 145.665 202.455 ;
        RECT 145.835 202.375 146.005 202.625 ;
        RECT 146.795 202.715 147.055 202.965 ;
        RECT 147.225 202.895 147.510 203.765 ;
        RECT 146.795 202.545 147.550 202.715 ;
        RECT 147.735 202.675 150.325 203.765 ;
        RECT 145.835 202.205 146.975 202.375 ;
        RECT 147.145 202.035 147.550 202.545 ;
        RECT 145.900 201.865 147.550 202.035 ;
        RECT 147.735 201.985 148.945 202.505 ;
        RECT 149.115 202.155 150.325 202.675 ;
        RECT 150.965 202.705 151.295 203.555 ;
        RECT 144.975 201.385 145.275 201.715 ;
        RECT 145.445 201.215 145.720 201.695 ;
        RECT 145.900 201.475 146.195 201.865 ;
        RECT 146.365 201.215 146.620 201.695 ;
        RECT 146.795 201.475 147.055 201.865 ;
        RECT 147.225 201.215 147.505 201.695 ;
        RECT 147.735 201.215 150.325 201.985 ;
        RECT 150.965 201.940 151.155 202.705 ;
        RECT 151.465 202.625 151.715 203.765 ;
        RECT 151.905 203.125 152.155 203.545 ;
        RECT 152.385 203.295 152.715 203.765 ;
        RECT 152.945 203.125 153.195 203.545 ;
        RECT 151.905 202.955 153.195 203.125 ;
        RECT 153.375 203.125 153.705 203.555 ;
        RECT 153.375 202.955 153.830 203.125 ;
        RECT 151.895 202.455 152.110 202.785 ;
        RECT 151.325 202.125 151.635 202.455 ;
        RECT 151.805 202.125 152.110 202.455 ;
        RECT 152.285 202.125 152.570 202.785 ;
        RECT 152.765 202.125 153.030 202.785 ;
        RECT 153.245 202.125 153.490 202.785 ;
        RECT 151.465 201.955 151.635 202.125 ;
        RECT 153.660 201.955 153.830 202.955 ;
        RECT 154.175 202.675 156.765 203.765 ;
        RECT 150.965 201.430 151.295 201.940 ;
        RECT 151.465 201.785 153.830 201.955 ;
        RECT 154.175 201.985 155.385 202.505 ;
        RECT 155.555 202.155 156.765 202.675 ;
        RECT 156.935 202.675 158.145 203.765 ;
        RECT 156.935 202.135 157.455 202.675 ;
        RECT 151.465 201.215 151.795 201.615 ;
        RECT 152.845 201.445 153.175 201.785 ;
        RECT 153.345 201.215 153.675 201.615 ;
        RECT 154.175 201.215 156.765 201.985 ;
        RECT 157.625 201.965 158.145 202.505 ;
        RECT 156.935 201.215 158.145 201.965 ;
        RECT 2.750 201.045 158.230 201.215 ;
        RECT 2.835 200.295 4.045 201.045 ;
        RECT 4.220 200.495 4.475 200.785 ;
        RECT 4.645 200.665 4.975 201.045 ;
        RECT 4.220 200.325 4.970 200.495 ;
        RECT 2.835 199.755 3.355 200.295 ;
        RECT 3.525 199.585 4.045 200.125 ;
        RECT 2.835 198.495 4.045 199.585 ;
        RECT 4.220 199.505 4.570 200.155 ;
        RECT 4.740 199.335 4.970 200.325 ;
        RECT 4.220 199.165 4.970 199.335 ;
        RECT 4.220 198.665 4.475 199.165 ;
        RECT 4.645 198.495 4.975 198.995 ;
        RECT 5.145 198.665 5.315 200.785 ;
        RECT 5.675 200.685 6.005 201.045 ;
        RECT 6.175 200.655 6.670 200.825 ;
        RECT 6.875 200.655 7.730 200.825 ;
        RECT 5.545 199.465 6.005 200.515 ;
        RECT 5.485 198.680 5.810 199.465 ;
        RECT 6.175 199.295 6.345 200.655 ;
        RECT 6.515 199.745 6.865 200.365 ;
        RECT 7.035 200.145 7.390 200.365 ;
        RECT 7.035 199.555 7.205 200.145 ;
        RECT 7.560 199.945 7.730 200.655 ;
        RECT 8.605 200.585 8.935 201.045 ;
        RECT 9.145 200.685 9.495 200.855 ;
        RECT 7.935 200.115 8.725 200.365 ;
        RECT 9.145 200.295 9.405 200.685 ;
        RECT 9.715 200.595 10.665 200.875 ;
        RECT 10.835 200.605 11.025 201.045 ;
        RECT 11.195 200.665 12.265 200.835 ;
        RECT 8.895 199.945 9.065 200.125 ;
        RECT 6.175 199.125 6.570 199.295 ;
        RECT 6.740 199.165 7.205 199.555 ;
        RECT 7.375 199.775 9.065 199.945 ;
        RECT 6.400 198.995 6.570 199.125 ;
        RECT 7.375 198.995 7.545 199.775 ;
        RECT 9.235 199.605 9.405 200.295 ;
        RECT 7.905 199.435 9.405 199.605 ;
        RECT 9.595 199.635 9.805 200.425 ;
        RECT 9.975 199.805 10.325 200.425 ;
        RECT 10.495 199.815 10.665 200.595 ;
        RECT 11.195 200.435 11.365 200.665 ;
        RECT 10.835 200.265 11.365 200.435 ;
        RECT 10.835 199.985 11.055 200.265 ;
        RECT 11.535 200.095 11.775 200.495 ;
        RECT 10.495 199.645 10.900 199.815 ;
        RECT 11.235 199.725 11.775 200.095 ;
        RECT 11.945 200.310 12.265 200.665 ;
        RECT 12.510 200.585 12.815 201.045 ;
        RECT 12.985 200.335 13.240 200.865 ;
        RECT 11.945 200.135 12.270 200.310 ;
        RECT 11.945 199.835 12.860 200.135 ;
        RECT 12.120 199.805 12.860 199.835 ;
        RECT 9.595 199.475 10.270 199.635 ;
        RECT 10.730 199.555 10.900 199.645 ;
        RECT 9.595 199.465 10.560 199.475 ;
        RECT 9.235 199.295 9.405 199.435 ;
        RECT 5.980 198.495 6.230 198.955 ;
        RECT 6.400 198.665 6.650 198.995 ;
        RECT 6.865 198.665 7.545 198.995 ;
        RECT 7.715 199.095 8.790 199.265 ;
        RECT 9.235 199.125 9.795 199.295 ;
        RECT 10.100 199.175 10.560 199.465 ;
        RECT 10.730 199.385 11.950 199.555 ;
        RECT 7.715 198.755 7.885 199.095 ;
        RECT 8.120 198.495 8.450 198.925 ;
        RECT 8.620 198.755 8.790 199.095 ;
        RECT 9.085 198.495 9.455 198.955 ;
        RECT 9.625 198.665 9.795 199.125 ;
        RECT 10.730 199.005 10.900 199.385 ;
        RECT 12.120 199.215 12.290 199.805 ;
        RECT 13.030 199.685 13.240 200.335 ;
        RECT 13.420 200.495 13.675 200.785 ;
        RECT 13.845 200.665 14.175 201.045 ;
        RECT 13.420 200.325 14.170 200.495 ;
        RECT 10.030 198.665 10.900 199.005 ;
        RECT 11.490 199.045 12.290 199.215 ;
        RECT 11.070 198.495 11.320 198.955 ;
        RECT 11.490 198.755 11.660 199.045 ;
        RECT 11.840 198.495 12.170 198.875 ;
        RECT 12.510 198.495 12.815 199.635 ;
        RECT 12.985 198.805 13.240 199.685 ;
        RECT 13.420 199.505 13.770 200.155 ;
        RECT 13.940 199.335 14.170 200.325 ;
        RECT 13.420 199.165 14.170 199.335 ;
        RECT 13.420 198.665 13.675 199.165 ;
        RECT 13.845 198.495 14.175 198.995 ;
        RECT 14.345 198.665 14.515 200.785 ;
        RECT 14.875 200.685 15.205 201.045 ;
        RECT 15.375 200.655 15.870 200.825 ;
        RECT 16.075 200.655 16.930 200.825 ;
        RECT 14.745 199.465 15.205 200.515 ;
        RECT 14.685 198.680 15.010 199.465 ;
        RECT 15.375 199.295 15.545 200.655 ;
        RECT 15.715 199.745 16.065 200.365 ;
        RECT 16.235 200.145 16.590 200.365 ;
        RECT 16.235 199.555 16.405 200.145 ;
        RECT 16.760 199.945 16.930 200.655 ;
        RECT 17.805 200.585 18.135 201.045 ;
        RECT 18.345 200.685 18.695 200.855 ;
        RECT 17.135 200.115 17.925 200.365 ;
        RECT 18.345 200.295 18.605 200.685 ;
        RECT 18.915 200.595 19.865 200.875 ;
        RECT 20.035 200.605 20.225 201.045 ;
        RECT 20.395 200.665 21.465 200.835 ;
        RECT 18.095 199.945 18.265 200.125 ;
        RECT 15.375 199.125 15.770 199.295 ;
        RECT 15.940 199.165 16.405 199.555 ;
        RECT 16.575 199.775 18.265 199.945 ;
        RECT 15.600 198.995 15.770 199.125 ;
        RECT 16.575 198.995 16.745 199.775 ;
        RECT 18.435 199.605 18.605 200.295 ;
        RECT 17.105 199.435 18.605 199.605 ;
        RECT 18.795 199.635 19.005 200.425 ;
        RECT 19.175 199.805 19.525 200.425 ;
        RECT 19.695 199.815 19.865 200.595 ;
        RECT 20.395 200.435 20.565 200.665 ;
        RECT 20.035 200.265 20.565 200.435 ;
        RECT 20.035 199.985 20.255 200.265 ;
        RECT 20.735 200.095 20.975 200.495 ;
        RECT 19.695 199.645 20.100 199.815 ;
        RECT 20.435 199.725 20.975 200.095 ;
        RECT 21.145 200.310 21.465 200.665 ;
        RECT 21.710 200.585 22.015 201.045 ;
        RECT 22.185 200.335 22.440 200.865 ;
        RECT 21.145 200.135 21.470 200.310 ;
        RECT 21.145 199.835 22.060 200.135 ;
        RECT 21.320 199.805 22.060 199.835 ;
        RECT 18.795 199.475 19.470 199.635 ;
        RECT 19.930 199.555 20.100 199.645 ;
        RECT 18.795 199.465 19.760 199.475 ;
        RECT 18.435 199.295 18.605 199.435 ;
        RECT 15.180 198.495 15.430 198.955 ;
        RECT 15.600 198.665 15.850 198.995 ;
        RECT 16.065 198.665 16.745 198.995 ;
        RECT 16.915 199.095 17.990 199.265 ;
        RECT 18.435 199.125 18.995 199.295 ;
        RECT 19.300 199.175 19.760 199.465 ;
        RECT 19.930 199.385 21.150 199.555 ;
        RECT 16.915 198.755 17.085 199.095 ;
        RECT 17.320 198.495 17.650 198.925 ;
        RECT 17.820 198.755 17.990 199.095 ;
        RECT 18.285 198.495 18.655 198.955 ;
        RECT 18.825 198.665 18.995 199.125 ;
        RECT 19.930 199.005 20.100 199.385 ;
        RECT 21.320 199.215 21.490 199.805 ;
        RECT 22.230 199.685 22.440 200.335 ;
        RECT 19.230 198.665 20.100 199.005 ;
        RECT 20.690 199.045 21.490 199.215 ;
        RECT 20.270 198.495 20.520 198.955 ;
        RECT 20.690 198.755 20.860 199.045 ;
        RECT 21.040 198.495 21.370 198.875 ;
        RECT 21.710 198.495 22.015 199.635 ;
        RECT 22.185 198.805 22.440 199.685 ;
        RECT 22.620 200.505 22.875 200.835 ;
        RECT 23.045 200.665 23.375 201.045 ;
        RECT 24.505 200.665 25.760 200.835 ;
        RECT 25.945 200.665 26.275 201.045 ;
        RECT 22.620 199.635 22.790 200.505 ;
        RECT 23.100 200.325 25.380 200.495 ;
        RECT 23.100 200.135 23.270 200.325 ;
        RECT 25.210 200.135 25.380 200.325 ;
        RECT 25.590 200.475 25.760 200.665 ;
        RECT 26.445 200.495 26.615 200.875 ;
        RECT 26.785 200.665 27.115 201.045 ;
        RECT 27.285 200.495 27.455 200.875 ;
        RECT 27.625 200.665 27.955 201.045 ;
        RECT 25.590 200.305 26.265 200.475 ;
        RECT 26.445 200.325 27.960 200.495 ;
        RECT 22.960 199.805 23.270 200.135 ;
        RECT 23.440 199.635 23.610 200.135 ;
        RECT 22.620 199.465 23.610 199.635 ;
        RECT 24.010 199.515 24.280 200.135 ;
        RECT 24.495 199.805 24.965 200.135 ;
        RECT 25.210 199.805 25.925 200.135 ;
        RECT 26.095 200.055 26.265 200.305 ;
        RECT 26.095 199.885 27.560 200.055 ;
        RECT 26.095 199.535 26.265 199.885 ;
        RECT 27.730 199.555 27.960 200.325 ;
        RECT 28.595 200.320 28.885 201.045 ;
        RECT 29.515 200.370 29.775 200.875 ;
        RECT 29.955 200.665 30.285 201.045 ;
        RECT 30.465 200.495 30.635 200.875 ;
        RECT 22.620 198.665 22.875 199.465 ;
        RECT 24.510 199.365 26.265 199.535 ;
        RECT 26.095 199.345 26.265 199.365 ;
        RECT 26.445 199.385 27.960 199.555 ;
        RECT 23.045 198.495 23.350 199.295 ;
        RECT 23.520 198.855 23.870 199.195 ;
        RECT 24.060 199.025 25.775 199.195 ;
        RECT 23.520 198.685 25.300 198.855 ;
        RECT 25.605 198.665 25.775 199.025 ;
        RECT 25.945 198.495 26.275 198.875 ;
        RECT 26.445 198.665 26.615 199.385 ;
        RECT 26.785 198.495 27.115 199.215 ;
        RECT 27.285 198.665 27.455 199.385 ;
        RECT 27.625 198.495 27.955 199.215 ;
        RECT 28.595 198.495 28.885 199.660 ;
        RECT 29.515 199.570 29.685 200.370 ;
        RECT 29.970 200.325 30.635 200.495 ;
        RECT 29.970 200.070 30.140 200.325 ;
        RECT 31.360 200.305 31.615 200.875 ;
        RECT 31.785 200.645 32.115 201.045 ;
        RECT 32.540 200.510 33.070 200.875 ;
        RECT 32.540 200.475 32.715 200.510 ;
        RECT 31.785 200.305 32.715 200.475 ;
        RECT 33.260 200.365 33.535 200.875 ;
        RECT 29.855 199.740 30.140 200.070 ;
        RECT 30.375 199.775 30.705 200.145 ;
        RECT 29.970 199.595 30.140 199.740 ;
        RECT 31.360 199.635 31.530 200.305 ;
        RECT 31.785 200.135 31.955 200.305 ;
        RECT 31.700 199.805 31.955 200.135 ;
        RECT 32.180 199.805 32.375 200.135 ;
        RECT 29.515 198.665 29.785 199.570 ;
        RECT 29.970 199.425 30.635 199.595 ;
        RECT 29.955 198.495 30.285 199.255 ;
        RECT 30.465 198.665 30.635 199.425 ;
        RECT 31.360 198.665 31.695 199.635 ;
        RECT 31.865 198.495 32.035 199.635 ;
        RECT 32.205 198.835 32.375 199.805 ;
        RECT 32.545 199.175 32.715 200.305 ;
        RECT 32.885 199.515 33.055 200.315 ;
        RECT 33.255 200.195 33.535 200.365 ;
        RECT 33.260 199.715 33.535 200.195 ;
        RECT 33.705 199.515 33.895 200.875 ;
        RECT 34.075 200.510 34.585 201.045 ;
        RECT 34.805 200.235 35.050 200.840 ;
        RECT 35.770 200.235 36.015 200.840 ;
        RECT 36.235 200.510 36.745 201.045 ;
        RECT 34.095 200.065 35.325 200.235 ;
        RECT 32.885 199.345 33.895 199.515 ;
        RECT 34.065 199.500 34.815 199.690 ;
        RECT 32.545 199.005 33.670 199.175 ;
        RECT 34.065 198.835 34.235 199.500 ;
        RECT 34.985 199.255 35.325 200.065 ;
        RECT 32.205 198.665 34.235 198.835 ;
        RECT 34.405 198.495 34.575 199.255 ;
        RECT 34.810 198.845 35.325 199.255 ;
        RECT 35.495 200.065 36.725 200.235 ;
        RECT 35.495 199.255 35.835 200.065 ;
        RECT 36.005 199.500 36.755 199.690 ;
        RECT 35.495 198.845 36.010 199.255 ;
        RECT 36.245 198.495 36.415 199.255 ;
        RECT 36.585 198.835 36.755 199.500 ;
        RECT 36.925 199.515 37.115 200.875 ;
        RECT 37.285 200.025 37.560 200.875 ;
        RECT 37.750 200.510 38.280 200.875 ;
        RECT 38.705 200.645 39.035 201.045 ;
        RECT 38.105 200.475 38.280 200.510 ;
        RECT 37.285 199.855 37.565 200.025 ;
        RECT 37.285 199.715 37.560 199.855 ;
        RECT 37.765 199.515 37.935 200.315 ;
        RECT 36.925 199.345 37.935 199.515 ;
        RECT 38.105 200.305 39.035 200.475 ;
        RECT 39.205 200.305 39.460 200.875 ;
        RECT 38.105 199.175 38.275 200.305 ;
        RECT 38.865 200.135 39.035 200.305 ;
        RECT 37.150 199.005 38.275 199.175 ;
        RECT 38.445 199.805 38.640 200.135 ;
        RECT 38.865 199.805 39.120 200.135 ;
        RECT 38.445 198.835 38.615 199.805 ;
        RECT 39.290 199.635 39.460 200.305 ;
        RECT 36.585 198.665 38.615 198.835 ;
        RECT 38.785 198.495 38.955 199.635 ;
        RECT 39.125 198.665 39.460 199.635 ;
        RECT 40.095 200.395 40.355 200.875 ;
        RECT 40.525 200.505 40.775 201.045 ;
        RECT 40.095 199.365 40.265 200.395 ;
        RECT 40.945 200.340 41.165 200.825 ;
        RECT 40.435 199.745 40.665 200.140 ;
        RECT 40.835 199.915 41.165 200.340 ;
        RECT 41.335 200.665 42.225 200.835 ;
        RECT 41.335 199.940 41.505 200.665 ;
        RECT 41.675 200.110 42.225 200.495 ;
        RECT 42.485 200.395 42.655 200.875 ;
        RECT 42.825 200.565 43.155 201.045 ;
        RECT 43.380 200.625 44.915 200.875 ;
        RECT 43.380 200.395 43.550 200.625 ;
        RECT 42.485 200.225 43.550 200.395 ;
        RECT 43.730 200.055 44.010 200.455 ;
        RECT 41.335 199.870 42.225 199.940 ;
        RECT 41.330 199.845 42.225 199.870 ;
        RECT 42.400 199.845 42.750 200.055 ;
        RECT 42.920 199.855 43.365 200.055 ;
        RECT 43.535 199.855 44.010 200.055 ;
        RECT 44.280 200.055 44.565 200.455 ;
        RECT 44.745 200.395 44.915 200.625 ;
        RECT 45.085 200.565 45.415 201.045 ;
        RECT 45.630 200.545 45.885 200.875 ;
        RECT 45.700 200.465 45.885 200.545 ;
        RECT 44.745 200.225 45.545 200.395 ;
        RECT 44.280 199.855 44.610 200.055 ;
        RECT 44.780 200.025 45.145 200.055 ;
        RECT 44.780 199.855 45.155 200.025 ;
        RECT 41.320 199.830 42.225 199.845 ;
        RECT 41.315 199.815 42.225 199.830 ;
        RECT 41.305 199.810 42.225 199.815 ;
        RECT 41.300 199.800 42.225 199.810 ;
        RECT 41.295 199.790 42.225 199.800 ;
        RECT 41.285 199.785 42.225 199.790 ;
        RECT 41.275 199.775 42.225 199.785 ;
        RECT 41.265 199.770 42.225 199.775 ;
        RECT 41.265 199.765 41.600 199.770 ;
        RECT 41.250 199.760 41.600 199.765 ;
        RECT 41.235 199.750 41.600 199.760 ;
        RECT 41.210 199.745 41.600 199.750 ;
        RECT 40.435 199.740 41.600 199.745 ;
        RECT 40.435 199.705 41.570 199.740 ;
        RECT 40.435 199.680 41.535 199.705 ;
        RECT 40.435 199.650 41.505 199.680 ;
        RECT 40.435 199.620 41.485 199.650 ;
        RECT 40.435 199.590 41.465 199.620 ;
        RECT 40.435 199.580 41.395 199.590 ;
        RECT 40.435 199.570 41.370 199.580 ;
        RECT 40.435 199.555 41.350 199.570 ;
        RECT 40.435 199.540 41.330 199.555 ;
        RECT 40.540 199.530 41.325 199.540 ;
        RECT 40.540 199.495 41.310 199.530 ;
        RECT 40.095 198.665 40.370 199.365 ;
        RECT 40.540 199.245 41.295 199.495 ;
        RECT 41.465 199.175 41.795 199.420 ;
        RECT 41.965 199.320 42.225 199.770 ;
        RECT 45.375 199.675 45.545 200.225 ;
        RECT 42.485 199.505 45.545 199.675 ;
        RECT 41.610 199.150 41.795 199.175 ;
        RECT 41.610 199.050 42.225 199.150 ;
        RECT 40.540 198.495 40.795 199.040 ;
        RECT 40.965 198.665 41.445 199.005 ;
        RECT 41.620 198.495 42.225 199.050 ;
        RECT 42.485 198.665 42.655 199.505 ;
        RECT 45.715 199.345 45.885 200.465 ;
        RECT 46.165 200.395 46.335 200.875 ;
        RECT 46.505 200.565 46.835 201.045 ;
        RECT 47.060 200.625 48.595 200.875 ;
        RECT 47.060 200.395 47.230 200.625 ;
        RECT 46.165 200.225 47.230 200.395 ;
        RECT 47.410 200.055 47.690 200.455 ;
        RECT 46.080 199.845 46.430 200.055 ;
        RECT 46.600 199.855 47.045 200.055 ;
        RECT 47.215 199.855 47.690 200.055 ;
        RECT 47.960 200.055 48.245 200.455 ;
        RECT 48.425 200.395 48.595 200.625 ;
        RECT 48.765 200.565 49.095 201.045 ;
        RECT 49.310 200.545 49.565 200.875 ;
        RECT 49.380 200.465 49.565 200.545 ;
        RECT 48.425 200.225 49.225 200.395 ;
        RECT 47.960 199.855 48.290 200.055 ;
        RECT 48.460 199.855 48.825 200.055 ;
        RECT 49.055 199.675 49.225 200.225 ;
        RECT 45.675 199.335 45.885 199.345 ;
        RECT 42.825 198.835 43.155 199.335 ;
        RECT 43.325 199.095 44.960 199.335 ;
        RECT 43.325 199.005 43.555 199.095 ;
        RECT 43.665 198.835 43.995 198.875 ;
        RECT 42.825 198.665 43.995 198.835 ;
        RECT 44.185 198.495 44.540 198.915 ;
        RECT 44.710 198.665 44.960 199.095 ;
        RECT 45.130 198.495 45.460 199.255 ;
        RECT 45.630 198.665 45.885 199.335 ;
        RECT 46.165 199.505 49.225 199.675 ;
        RECT 46.165 198.665 46.335 199.505 ;
        RECT 49.395 199.335 49.565 200.465 ;
        RECT 46.505 198.835 46.835 199.335 ;
        RECT 47.005 199.095 48.640 199.335 ;
        RECT 47.005 199.005 47.235 199.095 ;
        RECT 47.345 198.835 47.675 198.875 ;
        RECT 46.505 198.665 47.675 198.835 ;
        RECT 47.865 198.495 48.220 198.915 ;
        RECT 48.390 198.665 48.640 199.095 ;
        RECT 48.810 198.495 49.140 199.255 ;
        RECT 49.310 198.665 49.565 199.335 ;
        RECT 49.775 200.545 50.030 200.875 ;
        RECT 50.245 200.565 50.575 201.045 ;
        RECT 50.745 200.625 52.280 200.875 ;
        RECT 49.775 200.535 49.985 200.545 ;
        RECT 49.775 200.465 49.960 200.535 ;
        RECT 49.775 199.335 49.945 200.465 ;
        RECT 50.745 200.395 50.915 200.625 ;
        RECT 50.115 200.225 50.915 200.395 ;
        RECT 50.115 199.675 50.285 200.225 ;
        RECT 51.095 200.055 51.380 200.455 ;
        RECT 50.515 199.855 50.880 200.055 ;
        RECT 51.050 199.855 51.380 200.055 ;
        RECT 51.650 200.055 51.930 200.455 ;
        RECT 52.110 200.395 52.280 200.625 ;
        RECT 52.505 200.565 52.835 201.045 ;
        RECT 53.005 200.395 53.175 200.875 ;
        RECT 52.110 200.225 53.175 200.395 ;
        RECT 54.355 200.320 54.645 201.045 ;
        RECT 54.815 200.395 55.075 200.875 ;
        RECT 55.245 200.505 55.495 201.045 ;
        RECT 51.650 199.855 52.125 200.055 ;
        RECT 52.295 199.855 52.740 200.055 ;
        RECT 52.910 199.845 53.260 200.055 ;
        RECT 50.115 199.505 53.175 199.675 ;
        RECT 49.775 198.665 50.030 199.335 ;
        RECT 50.200 198.495 50.530 199.255 ;
        RECT 50.700 199.095 52.335 199.335 ;
        RECT 50.700 198.665 50.950 199.095 ;
        RECT 52.105 199.005 52.335 199.095 ;
        RECT 51.120 198.495 51.475 198.915 ;
        RECT 51.665 198.835 51.995 198.875 ;
        RECT 52.505 198.835 52.835 199.335 ;
        RECT 51.665 198.665 52.835 198.835 ;
        RECT 53.005 198.665 53.175 199.505 ;
        RECT 54.355 198.495 54.645 199.660 ;
        RECT 54.815 199.365 54.985 200.395 ;
        RECT 55.665 200.365 55.885 200.825 ;
        RECT 55.635 200.340 55.885 200.365 ;
        RECT 55.155 199.745 55.385 200.140 ;
        RECT 55.555 199.915 55.885 200.340 ;
        RECT 56.055 200.665 56.945 200.835 ;
        RECT 56.055 199.940 56.225 200.665 ;
        RECT 56.395 200.110 56.945 200.495 ;
        RECT 57.120 200.205 57.380 201.045 ;
        RECT 57.555 200.300 57.810 200.875 ;
        RECT 57.980 200.665 58.310 201.045 ;
        RECT 58.525 200.495 58.695 200.875 ;
        RECT 57.980 200.325 58.695 200.495 ;
        RECT 56.055 199.870 56.945 199.940 ;
        RECT 56.050 199.845 56.945 199.870 ;
        RECT 56.040 199.830 56.945 199.845 ;
        RECT 56.035 199.815 56.945 199.830 ;
        RECT 56.025 199.810 56.945 199.815 ;
        RECT 56.020 199.800 56.945 199.810 ;
        RECT 56.015 199.790 56.945 199.800 ;
        RECT 56.005 199.785 56.945 199.790 ;
        RECT 55.995 199.775 56.945 199.785 ;
        RECT 55.985 199.770 56.945 199.775 ;
        RECT 55.985 199.765 56.320 199.770 ;
        RECT 55.970 199.760 56.320 199.765 ;
        RECT 55.955 199.750 56.320 199.760 ;
        RECT 55.930 199.745 56.320 199.750 ;
        RECT 55.155 199.740 56.320 199.745 ;
        RECT 55.155 199.705 56.290 199.740 ;
        RECT 55.155 199.680 56.255 199.705 ;
        RECT 55.155 199.650 56.225 199.680 ;
        RECT 55.155 199.620 56.205 199.650 ;
        RECT 55.155 199.590 56.185 199.620 ;
        RECT 55.155 199.580 56.115 199.590 ;
        RECT 55.155 199.570 56.090 199.580 ;
        RECT 55.155 199.555 56.070 199.570 ;
        RECT 55.155 199.540 56.050 199.555 ;
        RECT 55.260 199.530 56.045 199.540 ;
        RECT 55.260 199.495 56.030 199.530 ;
        RECT 54.815 198.665 55.090 199.365 ;
        RECT 55.260 199.245 56.015 199.495 ;
        RECT 56.185 199.175 56.515 199.420 ;
        RECT 56.685 199.320 56.945 199.770 ;
        RECT 56.330 199.150 56.515 199.175 ;
        RECT 56.330 199.050 56.945 199.150 ;
        RECT 55.260 198.495 55.515 199.040 ;
        RECT 55.685 198.665 56.165 199.005 ;
        RECT 56.340 198.495 56.945 199.050 ;
        RECT 57.120 198.495 57.380 199.645 ;
        RECT 57.555 199.570 57.725 200.300 ;
        RECT 57.980 200.135 58.150 200.325 ;
        RECT 58.965 200.315 59.265 201.045 ;
        RECT 57.895 199.805 58.150 200.135 ;
        RECT 57.980 199.595 58.150 199.805 ;
        RECT 58.430 199.775 58.785 200.145 ;
        RECT 59.445 200.135 59.675 200.755 ;
        RECT 59.875 200.485 60.100 200.865 ;
        RECT 60.270 200.655 60.600 201.045 ;
        RECT 59.875 200.305 60.205 200.485 ;
        RECT 58.970 199.805 59.265 200.135 ;
        RECT 59.445 199.805 59.860 200.135 ;
        RECT 60.030 199.635 60.205 200.305 ;
        RECT 60.375 199.805 60.615 200.455 ;
        RECT 60.805 200.315 61.105 201.045 ;
        RECT 61.285 200.135 61.515 200.755 ;
        RECT 61.715 200.485 61.940 200.865 ;
        RECT 62.110 200.655 62.440 201.045 ;
        RECT 62.635 200.500 67.980 201.045 ;
        RECT 68.155 200.500 73.500 201.045 ;
        RECT 73.675 200.500 79.020 201.045 ;
        RECT 61.715 200.305 62.045 200.485 ;
        RECT 60.810 199.805 61.105 200.135 ;
        RECT 61.285 199.805 61.700 200.135 ;
        RECT 61.870 199.635 62.045 200.305 ;
        RECT 62.215 199.805 62.455 200.455 ;
        RECT 64.220 199.670 64.560 200.500 ;
        RECT 57.555 198.665 57.810 199.570 ;
        RECT 57.980 199.425 58.695 199.595 ;
        RECT 57.980 198.495 58.310 199.255 ;
        RECT 58.525 198.665 58.695 199.425 ;
        RECT 58.965 199.275 59.860 199.605 ;
        RECT 60.030 199.445 60.615 199.635 ;
        RECT 58.965 199.105 60.170 199.275 ;
        RECT 58.965 198.675 59.295 199.105 ;
        RECT 59.475 198.495 59.670 198.935 ;
        RECT 59.840 198.675 60.170 199.105 ;
        RECT 60.340 198.675 60.615 199.445 ;
        RECT 60.805 199.275 61.700 199.605 ;
        RECT 61.870 199.445 62.455 199.635 ;
        RECT 60.805 199.105 62.010 199.275 ;
        RECT 60.805 198.675 61.135 199.105 ;
        RECT 61.315 198.495 61.510 198.935 ;
        RECT 61.680 198.675 62.010 199.105 ;
        RECT 62.180 198.675 62.455 199.445 ;
        RECT 66.040 198.930 66.390 200.180 ;
        RECT 69.740 199.670 70.080 200.500 ;
        RECT 71.560 198.930 71.910 200.180 ;
        RECT 75.260 199.670 75.600 200.500 ;
        RECT 80.115 200.320 80.405 201.045 ;
        RECT 80.575 200.275 84.085 201.045 ;
        RECT 77.080 198.930 77.430 200.180 ;
        RECT 80.575 199.755 82.225 200.275 ;
        RECT 62.635 198.495 67.980 198.930 ;
        RECT 68.155 198.495 73.500 198.930 ;
        RECT 73.675 198.495 79.020 198.930 ;
        RECT 80.115 198.495 80.405 199.660 ;
        RECT 82.395 199.585 84.085 200.105 ;
        RECT 80.575 198.495 84.085 199.585 ;
        RECT 84.725 198.665 84.985 200.875 ;
        RECT 85.165 200.565 85.475 201.045 ;
        RECT 85.655 200.395 85.995 200.875 ;
        RECT 85.325 200.225 85.995 200.395 ;
        RECT 85.325 200.135 85.495 200.225 ;
        RECT 85.155 199.805 85.495 200.135 ;
        RECT 86.165 200.055 86.375 200.740 ;
        RECT 85.895 199.805 86.375 200.055 ;
        RECT 86.555 199.805 86.825 200.740 ;
        RECT 87.075 200.135 87.320 200.740 ;
        RECT 87.500 200.425 87.790 200.875 ;
        RECT 87.960 200.595 88.250 201.045 ;
        RECT 88.420 200.425 88.685 200.875 ;
        RECT 88.905 200.575 89.195 201.045 ;
        RECT 87.500 200.255 88.685 200.425 ;
        RECT 89.365 200.405 89.695 200.875 ;
        RECT 89.865 200.575 90.035 201.045 ;
        RECT 90.205 200.405 90.535 200.875 ;
        RECT 89.365 200.395 90.535 200.405 ;
        RECT 88.935 200.225 90.535 200.395 ;
        RECT 90.705 200.225 90.980 201.045 ;
        RECT 91.155 200.275 94.665 201.045 ;
        RECT 95.845 200.475 96.015 200.875 ;
        RECT 96.255 200.645 96.585 201.045 ;
        RECT 96.855 200.705 98.260 200.875 ;
        RECT 96.855 200.475 97.025 200.705 ;
        RECT 95.845 200.305 97.025 200.475 ;
        RECT 98.090 200.475 98.260 200.705 ;
        RECT 98.430 200.665 98.760 201.045 ;
        RECT 87.075 199.805 87.335 200.135 ;
        RECT 87.680 199.805 88.165 200.055 ;
        RECT 85.325 199.635 85.495 199.805 ;
        RECT 85.325 199.465 87.810 199.635 ;
        RECT 85.155 198.495 85.965 199.295 ;
        RECT 86.135 198.665 86.465 199.465 ;
        RECT 86.650 198.495 87.390 199.295 ;
        RECT 87.560 198.665 87.810 199.465 ;
        RECT 87.980 198.715 88.165 199.805 ;
        RECT 88.335 199.470 88.665 200.055 ;
        RECT 88.935 199.685 89.150 200.225 ;
        RECT 89.320 199.855 90.090 200.055 ;
        RECT 90.260 199.855 90.980 200.055 ;
        RECT 91.155 199.755 92.805 200.275 ;
        RECT 97.195 200.135 97.385 200.365 ;
        RECT 88.935 199.465 89.695 199.685 ;
        RECT 88.360 198.495 88.685 199.295 ;
        RECT 88.895 198.835 89.195 199.295 ;
        RECT 89.365 199.005 89.695 199.465 ;
        RECT 89.865 199.465 90.980 199.675 ;
        RECT 92.975 199.585 94.665 200.105 ;
        RECT 95.815 199.805 96.000 200.135 ;
        RECT 96.255 199.805 96.730 200.135 ;
        RECT 97.040 199.805 97.385 200.135 ;
        RECT 97.645 199.805 97.840 200.380 ;
        RECT 98.090 200.305 98.785 200.475 ;
        RECT 98.955 200.460 99.265 200.875 ;
        RECT 98.615 200.135 98.785 200.305 ;
        RECT 98.110 199.805 98.445 200.135 ;
        RECT 98.615 199.805 98.925 200.135 ;
        RECT 98.615 199.635 98.785 199.805 ;
        RECT 89.865 198.835 90.035 199.465 ;
        RECT 88.895 198.665 90.035 198.835 ;
        RECT 90.205 198.495 90.535 199.295 ;
        RECT 90.705 198.665 90.980 199.465 ;
        RECT 91.155 198.495 94.665 199.585 ;
        RECT 95.845 199.465 98.785 199.635 ;
        RECT 95.845 198.665 96.015 199.465 ;
        RECT 99.095 199.345 99.265 200.460 ;
        RECT 99.445 200.315 99.745 201.045 ;
        RECT 99.925 200.135 100.155 200.755 ;
        RECT 100.355 200.485 100.580 200.865 ;
        RECT 100.750 200.655 101.080 201.045 ;
        RECT 100.355 200.305 100.685 200.485 ;
        RECT 99.450 199.805 99.745 200.135 ;
        RECT 99.925 199.805 100.340 200.135 ;
        RECT 100.510 199.635 100.685 200.305 ;
        RECT 100.855 199.805 101.095 200.455 ;
        RECT 101.275 200.275 104.785 201.045 ;
        RECT 105.875 200.320 106.165 201.045 ;
        RECT 106.335 200.460 106.645 200.875 ;
        RECT 106.840 200.665 107.170 201.045 ;
        RECT 107.340 200.705 108.745 200.875 ;
        RECT 107.340 200.475 107.510 200.705 ;
        RECT 101.275 199.755 102.925 200.275 ;
        RECT 96.775 199.125 98.335 199.295 ;
        RECT 96.775 198.665 97.025 199.125 ;
        RECT 97.225 198.495 97.895 198.875 ;
        RECT 98.085 198.665 98.335 199.125 ;
        RECT 98.510 198.495 98.755 198.955 ;
        RECT 98.925 198.705 99.265 199.345 ;
        RECT 99.445 199.275 100.340 199.605 ;
        RECT 100.510 199.445 101.095 199.635 ;
        RECT 103.095 199.585 104.785 200.105 ;
        RECT 99.445 199.105 100.650 199.275 ;
        RECT 99.445 198.675 99.775 199.105 ;
        RECT 99.955 198.495 100.150 198.935 ;
        RECT 100.320 198.675 100.650 199.105 ;
        RECT 100.820 198.675 101.095 199.445 ;
        RECT 101.275 198.495 104.785 199.585 ;
        RECT 105.875 198.495 106.165 199.660 ;
        RECT 106.335 199.345 106.505 200.460 ;
        RECT 106.815 200.305 107.510 200.475 ;
        RECT 108.575 200.475 108.745 200.705 ;
        RECT 109.015 200.645 109.345 201.045 ;
        RECT 109.585 200.475 109.755 200.875 ;
        RECT 110.015 200.500 115.360 201.045 ;
        RECT 106.815 200.135 106.985 200.305 ;
        RECT 106.675 199.805 106.985 200.135 ;
        RECT 107.155 199.805 107.490 200.135 ;
        RECT 107.760 199.805 107.955 200.380 ;
        RECT 108.215 200.135 108.405 200.365 ;
        RECT 108.575 200.305 109.755 200.475 ;
        RECT 108.215 199.805 108.560 200.135 ;
        RECT 108.870 199.805 109.345 200.135 ;
        RECT 109.600 199.805 109.785 200.135 ;
        RECT 106.815 199.635 106.985 199.805 ;
        RECT 111.600 199.670 111.940 200.500 ;
        RECT 115.535 200.275 118.125 201.045 ;
        RECT 118.755 200.665 119.645 200.835 ;
        RECT 106.815 199.465 109.755 199.635 ;
        RECT 106.335 198.705 106.675 199.345 ;
        RECT 107.265 199.125 108.825 199.295 ;
        RECT 106.845 198.495 107.090 198.955 ;
        RECT 107.265 198.665 107.515 199.125 ;
        RECT 107.705 198.495 108.375 198.875 ;
        RECT 108.575 198.665 108.825 199.125 ;
        RECT 109.585 198.665 109.755 199.465 ;
        RECT 113.420 198.930 113.770 200.180 ;
        RECT 115.535 199.755 116.745 200.275 ;
        RECT 118.755 200.110 119.305 200.495 ;
        RECT 116.915 199.585 118.125 200.105 ;
        RECT 119.475 199.940 119.645 200.665 ;
        RECT 110.015 198.495 115.360 198.930 ;
        RECT 115.535 198.495 118.125 199.585 ;
        RECT 118.755 199.870 119.645 199.940 ;
        RECT 119.815 200.340 120.035 200.825 ;
        RECT 120.205 200.505 120.455 201.045 ;
        RECT 120.625 200.395 120.885 200.875 ;
        RECT 121.080 200.655 121.410 201.045 ;
        RECT 121.580 200.485 121.805 200.865 ;
        RECT 119.815 199.915 120.145 200.340 ;
        RECT 118.755 199.845 119.650 199.870 ;
        RECT 118.755 199.830 119.660 199.845 ;
        RECT 118.755 199.815 119.665 199.830 ;
        RECT 118.755 199.810 119.675 199.815 ;
        RECT 118.755 199.800 119.680 199.810 ;
        RECT 118.755 199.790 119.685 199.800 ;
        RECT 118.755 199.785 119.695 199.790 ;
        RECT 118.755 199.775 119.705 199.785 ;
        RECT 118.755 199.770 119.715 199.775 ;
        RECT 118.755 199.320 119.015 199.770 ;
        RECT 119.380 199.765 119.715 199.770 ;
        RECT 119.380 199.760 119.730 199.765 ;
        RECT 119.380 199.750 119.745 199.760 ;
        RECT 119.380 199.745 119.770 199.750 ;
        RECT 120.315 199.745 120.545 200.140 ;
        RECT 119.380 199.740 120.545 199.745 ;
        RECT 119.410 199.705 120.545 199.740 ;
        RECT 119.445 199.680 120.545 199.705 ;
        RECT 119.475 199.650 120.545 199.680 ;
        RECT 119.495 199.620 120.545 199.650 ;
        RECT 119.515 199.590 120.545 199.620 ;
        RECT 119.585 199.580 120.545 199.590 ;
        RECT 119.610 199.570 120.545 199.580 ;
        RECT 119.630 199.555 120.545 199.570 ;
        RECT 119.650 199.540 120.545 199.555 ;
        RECT 119.655 199.530 120.440 199.540 ;
        RECT 119.670 199.495 120.440 199.530 ;
        RECT 119.185 199.175 119.515 199.420 ;
        RECT 119.685 199.245 120.440 199.495 ;
        RECT 120.715 199.365 120.885 200.395 ;
        RECT 121.065 199.805 121.305 200.455 ;
        RECT 121.475 200.305 121.805 200.485 ;
        RECT 121.475 199.635 121.650 200.305 ;
        RECT 122.005 200.135 122.235 200.755 ;
        RECT 122.415 200.315 122.715 201.045 ;
        RECT 122.935 200.225 123.165 201.045 ;
        RECT 123.335 200.245 123.665 200.875 ;
        RECT 121.820 199.805 122.235 200.135 ;
        RECT 122.415 199.805 122.710 200.135 ;
        RECT 122.915 199.805 123.245 200.055 ;
        RECT 123.415 199.645 123.665 200.245 ;
        RECT 123.835 200.225 124.045 201.045 ;
        RECT 124.280 200.515 124.570 200.865 ;
        RECT 124.765 200.685 125.095 201.045 ;
        RECT 125.265 200.515 125.495 200.820 ;
        RECT 124.280 200.345 125.495 200.515 ;
        RECT 125.685 200.705 125.855 200.740 ;
        RECT 125.685 200.535 125.885 200.705 ;
        RECT 125.685 200.175 125.855 200.535 ;
        RECT 124.340 200.025 124.600 200.135 ;
        RECT 124.335 199.855 124.600 200.025 ;
        RECT 124.340 199.805 124.600 199.855 ;
        RECT 124.780 199.805 125.165 200.135 ;
        RECT 125.335 200.005 125.855 200.175 ;
        RECT 126.115 200.295 127.325 201.045 ;
        RECT 127.495 200.305 127.935 200.865 ;
        RECT 128.105 200.305 128.555 201.045 ;
        RECT 128.725 200.475 128.895 200.875 ;
        RECT 129.065 200.645 129.485 201.045 ;
        RECT 129.655 200.475 129.885 200.875 ;
        RECT 128.725 200.305 129.885 200.475 ;
        RECT 130.055 200.305 130.545 200.875 ;
        RECT 131.635 200.320 131.925 201.045 ;
        RECT 119.185 199.150 119.370 199.175 ;
        RECT 118.755 199.050 119.370 199.150 ;
        RECT 118.755 198.495 119.360 199.050 ;
        RECT 119.535 198.665 120.015 199.005 ;
        RECT 120.185 198.495 120.440 199.040 ;
        RECT 120.610 198.665 120.885 199.365 ;
        RECT 121.065 199.445 121.650 199.635 ;
        RECT 121.065 198.675 121.340 199.445 ;
        RECT 121.820 199.275 122.715 199.605 ;
        RECT 121.510 199.105 122.715 199.275 ;
        RECT 121.510 198.675 121.840 199.105 ;
        RECT 122.010 198.495 122.205 198.935 ;
        RECT 122.385 198.675 122.715 199.105 ;
        RECT 122.935 198.495 123.165 199.635 ;
        RECT 123.335 198.665 123.665 199.645 ;
        RECT 123.835 198.495 124.045 199.635 ;
        RECT 124.280 198.495 124.600 199.635 ;
        RECT 124.780 198.755 124.975 199.805 ;
        RECT 125.335 199.625 125.505 200.005 ;
        RECT 125.155 199.345 125.505 199.625 ;
        RECT 125.695 199.475 125.940 199.835 ;
        RECT 126.115 199.755 126.635 200.295 ;
        RECT 126.805 199.585 127.325 200.125 ;
        RECT 125.155 198.665 125.485 199.345 ;
        RECT 125.685 198.495 125.940 199.295 ;
        RECT 126.115 198.495 127.325 199.585 ;
        RECT 127.495 199.295 127.805 200.305 ;
        RECT 127.975 199.685 128.145 200.135 ;
        RECT 128.315 199.855 128.705 200.135 ;
        RECT 128.890 199.805 129.135 200.135 ;
        RECT 127.975 199.515 128.765 199.685 ;
        RECT 127.495 198.665 127.935 199.295 ;
        RECT 128.110 198.495 128.425 199.345 ;
        RECT 128.595 198.835 128.765 199.515 ;
        RECT 128.935 199.005 129.135 199.805 ;
        RECT 129.335 199.005 129.585 200.135 ;
        RECT 129.800 199.805 130.205 200.135 ;
        RECT 130.375 199.635 130.545 200.305 ;
        RECT 132.095 200.100 132.435 200.875 ;
        RECT 132.605 200.585 132.775 201.045 ;
        RECT 133.015 200.610 133.375 200.875 ;
        RECT 133.015 200.605 133.370 200.610 ;
        RECT 133.015 200.595 133.365 200.605 ;
        RECT 133.015 200.590 133.360 200.595 ;
        RECT 133.015 200.580 133.355 200.590 ;
        RECT 134.005 200.585 134.175 201.045 ;
        RECT 133.015 200.575 133.350 200.580 ;
        RECT 133.015 200.565 133.340 200.575 ;
        RECT 133.015 200.555 133.330 200.565 ;
        RECT 133.015 200.415 133.315 200.555 ;
        RECT 132.605 200.225 133.315 200.415 ;
        RECT 133.505 200.415 133.835 200.495 ;
        RECT 134.345 200.415 134.685 200.875 ;
        RECT 134.855 200.500 140.200 201.045 ;
        RECT 133.505 200.225 134.685 200.415 ;
        RECT 129.775 199.465 130.545 199.635 ;
        RECT 129.775 198.835 130.025 199.465 ;
        RECT 128.595 198.665 130.025 198.835 ;
        RECT 130.205 198.495 130.535 199.295 ;
        RECT 131.635 198.495 131.925 199.660 ;
        RECT 132.095 198.665 132.375 200.100 ;
        RECT 132.605 199.655 132.890 200.225 ;
        RECT 133.075 199.825 133.545 200.055 ;
        RECT 133.715 200.035 134.045 200.055 ;
        RECT 133.715 199.855 134.165 200.035 ;
        RECT 134.355 199.855 134.685 200.055 ;
        RECT 132.605 199.440 133.755 199.655 ;
        RECT 132.545 198.495 133.255 199.270 ;
        RECT 133.425 198.665 133.755 199.440 ;
        RECT 133.950 198.740 134.165 199.855 ;
        RECT 134.455 199.515 134.685 199.855 ;
        RECT 136.440 199.670 136.780 200.500 ;
        RECT 140.375 200.295 141.585 201.045 ;
        RECT 141.840 200.545 142.335 200.875 ;
        RECT 134.345 198.495 134.675 199.215 ;
        RECT 138.260 198.930 138.610 200.180 ;
        RECT 140.375 199.755 140.895 200.295 ;
        RECT 141.065 199.585 141.585 200.125 ;
        RECT 134.855 198.495 140.200 198.930 ;
        RECT 140.375 198.495 141.585 199.585 ;
        RECT 141.755 199.055 141.995 200.365 ;
        RECT 142.165 199.635 142.335 200.545 ;
        RECT 142.555 199.805 142.905 200.770 ;
        RECT 143.085 199.805 143.385 200.775 ;
        RECT 143.565 199.805 143.845 200.775 ;
        RECT 144.025 200.245 144.295 201.045 ;
        RECT 144.465 200.325 144.805 200.835 ;
        RECT 144.040 199.805 144.370 200.055 ;
        RECT 144.040 199.635 144.355 199.805 ;
        RECT 142.165 199.465 144.355 199.635 ;
        RECT 141.760 198.495 142.095 198.875 ;
        RECT 142.265 198.665 142.515 199.465 ;
        RECT 142.735 198.495 143.065 199.215 ;
        RECT 143.250 198.665 143.500 199.465 ;
        RECT 143.965 198.495 144.295 199.295 ;
        RECT 144.545 198.925 144.805 200.325 ;
        RECT 144.985 200.315 145.285 201.045 ;
        RECT 145.465 200.135 145.695 200.755 ;
        RECT 145.895 200.485 146.120 200.865 ;
        RECT 146.290 200.655 146.620 201.045 ;
        RECT 145.895 200.305 146.225 200.485 ;
        RECT 144.990 199.805 145.285 200.135 ;
        RECT 145.465 199.805 145.880 200.135 ;
        RECT 146.050 199.635 146.225 200.305 ;
        RECT 146.395 199.805 146.635 200.455 ;
        RECT 146.815 200.275 149.405 201.045 ;
        RECT 146.815 199.755 148.025 200.275 ;
        RECT 149.575 200.245 149.915 200.875 ;
        RECT 150.085 200.245 150.335 201.045 ;
        RECT 150.525 200.395 150.855 200.875 ;
        RECT 151.025 200.585 151.250 201.045 ;
        RECT 151.420 200.395 151.750 200.875 ;
        RECT 144.465 198.665 144.805 198.925 ;
        RECT 144.985 199.275 145.880 199.605 ;
        RECT 146.050 199.445 146.635 199.635 ;
        RECT 148.195 199.585 149.405 200.105 ;
        RECT 144.985 199.105 146.190 199.275 ;
        RECT 144.985 198.675 145.315 199.105 ;
        RECT 145.495 198.495 145.690 198.935 ;
        RECT 145.860 198.675 146.190 199.105 ;
        RECT 146.360 198.675 146.635 199.445 ;
        RECT 146.815 198.495 149.405 199.585 ;
        RECT 149.575 199.635 149.750 200.245 ;
        RECT 150.525 200.225 151.750 200.395 ;
        RECT 152.380 200.265 152.880 200.875 ;
        RECT 153.255 200.275 156.765 201.045 ;
        RECT 156.935 200.295 158.145 201.045 ;
        RECT 149.920 199.885 150.615 200.055 ;
        RECT 150.445 199.635 150.615 199.885 ;
        RECT 150.790 199.855 151.210 200.055 ;
        RECT 151.380 199.855 151.710 200.055 ;
        RECT 151.880 199.855 152.210 200.055 ;
        RECT 152.380 199.635 152.550 200.265 ;
        RECT 152.735 199.805 153.085 200.055 ;
        RECT 153.255 199.755 154.905 200.275 ;
        RECT 149.575 198.665 149.915 199.635 ;
        RECT 150.085 198.495 150.255 199.635 ;
        RECT 150.445 199.465 152.880 199.635 ;
        RECT 155.075 199.585 156.765 200.105 ;
        RECT 150.525 198.495 150.775 199.295 ;
        RECT 151.420 198.665 151.750 199.465 ;
        RECT 152.050 198.495 152.380 199.295 ;
        RECT 152.550 198.665 152.880 199.465 ;
        RECT 153.255 198.495 156.765 199.585 ;
        RECT 156.935 199.585 157.455 200.125 ;
        RECT 157.625 199.755 158.145 200.295 ;
        RECT 156.935 198.495 158.145 199.585 ;
        RECT 2.750 198.325 158.230 198.495 ;
        RECT 2.835 197.235 4.045 198.325 ;
        RECT 4.215 197.235 5.885 198.325 ;
        RECT 2.835 196.525 3.355 197.065 ;
        RECT 3.525 196.695 4.045 197.235 ;
        RECT 4.215 196.545 4.965 197.065 ;
        RECT 5.135 196.715 5.885 197.235 ;
        RECT 6.055 197.250 6.325 198.155 ;
        RECT 6.495 197.565 6.825 198.325 ;
        RECT 7.005 197.395 7.175 198.155 ;
        RECT 2.835 195.775 4.045 196.525 ;
        RECT 4.215 195.775 5.885 196.545 ;
        RECT 6.055 196.450 6.225 197.250 ;
        RECT 6.510 197.225 7.175 197.395 ;
        RECT 6.510 197.080 6.680 197.225 ;
        RECT 6.395 196.750 6.680 197.080 ;
        RECT 7.440 197.185 7.775 198.155 ;
        RECT 7.945 197.185 8.115 198.325 ;
        RECT 8.285 197.985 10.315 198.155 ;
        RECT 6.510 196.495 6.680 196.750 ;
        RECT 6.915 196.675 7.245 197.045 ;
        RECT 7.440 196.515 7.610 197.185 ;
        RECT 8.285 197.015 8.455 197.985 ;
        RECT 7.780 196.685 8.035 197.015 ;
        RECT 8.260 196.685 8.455 197.015 ;
        RECT 8.625 197.645 9.750 197.815 ;
        RECT 7.865 196.515 8.035 196.685 ;
        RECT 8.625 196.515 8.795 197.645 ;
        RECT 6.055 195.945 6.315 196.450 ;
        RECT 6.510 196.325 7.175 196.495 ;
        RECT 6.495 195.775 6.825 196.155 ;
        RECT 7.005 195.945 7.175 196.325 ;
        RECT 7.440 195.945 7.695 196.515 ;
        RECT 7.865 196.345 8.795 196.515 ;
        RECT 8.965 197.305 9.975 197.475 ;
        RECT 8.965 196.505 9.135 197.305 ;
        RECT 9.340 196.625 9.615 197.105 ;
        RECT 9.335 196.455 9.615 196.625 ;
        RECT 8.620 196.310 8.795 196.345 ;
        RECT 7.865 195.775 8.195 196.175 ;
        RECT 8.620 195.945 9.150 196.310 ;
        RECT 9.340 195.945 9.615 196.455 ;
        RECT 9.785 195.945 9.975 197.305 ;
        RECT 10.145 197.320 10.315 197.985 ;
        RECT 10.485 197.565 10.655 198.325 ;
        RECT 10.890 197.565 11.405 197.975 ;
        RECT 10.145 197.130 10.895 197.320 ;
        RECT 11.065 196.755 11.405 197.565 ;
        RECT 10.175 196.585 11.405 196.755 ;
        RECT 11.575 197.565 12.090 197.975 ;
        RECT 12.325 197.565 12.495 198.325 ;
        RECT 12.665 197.985 14.695 198.155 ;
        RECT 11.575 196.755 11.915 197.565 ;
        RECT 12.665 197.320 12.835 197.985 ;
        RECT 13.230 197.645 14.355 197.815 ;
        RECT 12.085 197.130 12.835 197.320 ;
        RECT 13.005 197.305 14.015 197.475 ;
        RECT 11.575 196.585 12.805 196.755 ;
        RECT 10.155 195.775 10.665 196.310 ;
        RECT 10.885 195.980 11.130 196.585 ;
        RECT 11.850 195.980 12.095 196.585 ;
        RECT 12.315 195.775 12.825 196.310 ;
        RECT 13.005 195.945 13.195 197.305 ;
        RECT 13.365 196.965 13.640 197.105 ;
        RECT 13.365 196.795 13.645 196.965 ;
        RECT 13.365 195.945 13.640 196.795 ;
        RECT 13.845 196.505 14.015 197.305 ;
        RECT 14.185 196.515 14.355 197.645 ;
        RECT 14.525 197.015 14.695 197.985 ;
        RECT 14.865 197.185 15.035 198.325 ;
        RECT 15.205 197.185 15.540 198.155 ;
        RECT 14.525 196.685 14.720 197.015 ;
        RECT 14.945 196.685 15.200 197.015 ;
        RECT 14.945 196.515 15.115 196.685 ;
        RECT 15.370 196.515 15.540 197.185 ;
        RECT 15.715 197.160 16.005 198.325 ;
        RECT 16.175 197.250 16.445 198.155 ;
        RECT 16.615 197.565 16.945 198.325 ;
        RECT 17.125 197.395 17.295 198.155 ;
        RECT 14.185 196.345 15.115 196.515 ;
        RECT 14.185 196.310 14.360 196.345 ;
        RECT 13.830 195.945 14.360 196.310 ;
        RECT 14.785 195.775 15.115 196.175 ;
        RECT 15.285 195.945 15.540 196.515 ;
        RECT 15.715 195.775 16.005 196.500 ;
        RECT 16.175 196.450 16.345 197.250 ;
        RECT 16.630 197.225 17.295 197.395 ;
        RECT 16.630 197.080 16.800 197.225 ;
        RECT 16.515 196.750 16.800 197.080 ;
        RECT 17.560 197.185 17.895 198.155 ;
        RECT 18.065 197.185 18.235 198.325 ;
        RECT 18.405 197.985 20.435 198.155 ;
        RECT 16.630 196.495 16.800 196.750 ;
        RECT 17.035 196.675 17.365 197.045 ;
        RECT 17.560 196.515 17.730 197.185 ;
        RECT 18.405 197.015 18.575 197.985 ;
        RECT 17.900 196.685 18.155 197.015 ;
        RECT 18.380 196.685 18.575 197.015 ;
        RECT 18.745 197.645 19.870 197.815 ;
        RECT 17.985 196.515 18.155 196.685 ;
        RECT 18.745 196.515 18.915 197.645 ;
        RECT 16.175 195.945 16.435 196.450 ;
        RECT 16.630 196.325 17.295 196.495 ;
        RECT 16.615 195.775 16.945 196.155 ;
        RECT 17.125 195.945 17.295 196.325 ;
        RECT 17.560 195.945 17.815 196.515 ;
        RECT 17.985 196.345 18.915 196.515 ;
        RECT 19.085 197.305 20.095 197.475 ;
        RECT 19.085 196.505 19.255 197.305 ;
        RECT 18.740 196.310 18.915 196.345 ;
        RECT 17.985 195.775 18.315 196.175 ;
        RECT 18.740 195.945 19.270 196.310 ;
        RECT 19.460 196.285 19.735 197.105 ;
        RECT 19.455 196.115 19.735 196.285 ;
        RECT 19.460 195.945 19.735 196.115 ;
        RECT 19.905 195.945 20.095 197.305 ;
        RECT 20.265 197.320 20.435 197.985 ;
        RECT 20.605 197.565 20.775 198.325 ;
        RECT 21.010 197.565 21.525 197.975 ;
        RECT 20.265 197.130 21.015 197.320 ;
        RECT 21.185 196.755 21.525 197.565 ;
        RECT 21.700 197.935 22.035 198.155 ;
        RECT 23.040 197.945 23.395 198.325 ;
        RECT 21.700 197.315 21.955 197.935 ;
        RECT 22.205 197.775 22.435 197.815 ;
        RECT 23.565 197.775 23.815 198.155 ;
        RECT 22.205 197.575 23.815 197.775 ;
        RECT 22.205 197.485 22.390 197.575 ;
        RECT 22.980 197.565 23.815 197.575 ;
        RECT 24.065 197.545 24.315 198.325 ;
        RECT 24.485 197.475 24.745 198.155 ;
        RECT 22.545 197.375 22.875 197.405 ;
        RECT 22.545 197.315 24.345 197.375 ;
        RECT 21.700 197.205 24.405 197.315 ;
        RECT 21.700 197.145 22.875 197.205 ;
        RECT 24.205 197.170 24.405 197.205 ;
        RECT 21.695 196.765 22.185 196.965 ;
        RECT 22.375 196.765 22.850 196.975 ;
        RECT 20.295 196.585 21.525 196.755 ;
        RECT 20.275 195.775 20.785 196.310 ;
        RECT 21.005 195.980 21.250 196.585 ;
        RECT 21.700 195.775 22.155 196.540 ;
        RECT 22.630 196.365 22.850 196.765 ;
        RECT 23.095 196.765 23.425 196.975 ;
        RECT 23.095 196.365 23.305 196.765 ;
        RECT 23.595 196.730 24.005 197.035 ;
        RECT 24.235 196.595 24.405 197.170 ;
        RECT 24.135 196.475 24.405 196.595 ;
        RECT 23.560 196.430 24.405 196.475 ;
        RECT 23.560 196.305 24.315 196.430 ;
        RECT 23.560 196.155 23.730 196.305 ;
        RECT 24.575 196.275 24.745 197.475 ;
        RECT 22.430 195.945 23.730 196.155 ;
        RECT 23.985 195.775 24.315 196.135 ;
        RECT 24.485 195.945 24.745 196.275 ;
        RECT 24.915 197.355 25.225 198.155 ;
        RECT 25.395 197.525 25.705 198.325 ;
        RECT 25.875 197.695 26.135 198.155 ;
        RECT 26.305 197.865 26.560 198.325 ;
        RECT 26.735 197.695 26.995 198.155 ;
        RECT 25.875 197.525 26.995 197.695 ;
        RECT 24.915 197.185 25.945 197.355 ;
        RECT 24.915 196.275 25.085 197.185 ;
        RECT 25.255 196.445 25.605 197.015 ;
        RECT 25.775 196.935 25.945 197.185 ;
        RECT 26.735 197.275 26.995 197.525 ;
        RECT 27.165 197.455 27.450 198.325 ;
        RECT 27.680 197.655 27.935 198.155 ;
        RECT 28.105 197.825 28.435 198.325 ;
        RECT 27.680 197.485 28.430 197.655 ;
        RECT 26.735 197.105 27.490 197.275 ;
        RECT 25.775 196.765 26.915 196.935 ;
        RECT 27.085 196.595 27.490 197.105 ;
        RECT 27.680 196.665 28.030 197.315 ;
        RECT 25.840 196.425 27.490 196.595 ;
        RECT 28.200 196.495 28.430 197.485 ;
        RECT 24.915 195.945 25.215 196.275 ;
        RECT 25.385 195.775 25.660 196.255 ;
        RECT 25.840 196.035 26.135 196.425 ;
        RECT 26.305 195.775 26.560 196.255 ;
        RECT 26.735 196.035 26.995 196.425 ;
        RECT 27.680 196.325 28.430 196.495 ;
        RECT 27.165 195.775 27.445 196.255 ;
        RECT 27.680 196.035 27.935 196.325 ;
        RECT 28.105 195.775 28.435 196.155 ;
        RECT 28.605 196.035 28.775 198.155 ;
        RECT 28.945 197.355 29.270 198.140 ;
        RECT 29.440 197.865 29.690 198.325 ;
        RECT 29.860 197.825 30.110 198.155 ;
        RECT 30.325 197.825 31.005 198.155 ;
        RECT 29.860 197.695 30.030 197.825 ;
        RECT 29.635 197.525 30.030 197.695 ;
        RECT 29.005 196.305 29.465 197.355 ;
        RECT 29.635 196.165 29.805 197.525 ;
        RECT 30.200 197.265 30.665 197.655 ;
        RECT 29.975 196.455 30.325 197.075 ;
        RECT 30.495 196.675 30.665 197.265 ;
        RECT 30.835 197.045 31.005 197.825 ;
        RECT 31.175 197.725 31.345 198.065 ;
        RECT 31.580 197.895 31.910 198.325 ;
        RECT 32.080 197.725 32.250 198.065 ;
        RECT 32.545 197.865 32.915 198.325 ;
        RECT 31.175 197.555 32.250 197.725 ;
        RECT 33.085 197.695 33.255 198.155 ;
        RECT 33.490 197.815 34.360 198.155 ;
        RECT 34.530 197.865 34.780 198.325 ;
        RECT 32.695 197.525 33.255 197.695 ;
        RECT 32.695 197.385 32.865 197.525 ;
        RECT 31.365 197.215 32.865 197.385 ;
        RECT 33.560 197.355 34.020 197.645 ;
        RECT 30.835 196.875 32.525 197.045 ;
        RECT 30.495 196.455 30.850 196.675 ;
        RECT 31.020 196.165 31.190 196.875 ;
        RECT 31.395 196.455 32.185 196.705 ;
        RECT 32.355 196.695 32.525 196.875 ;
        RECT 32.695 196.525 32.865 197.215 ;
        RECT 29.135 195.775 29.465 196.135 ;
        RECT 29.635 195.995 30.130 196.165 ;
        RECT 30.335 195.995 31.190 196.165 ;
        RECT 32.065 195.775 32.395 196.235 ;
        RECT 32.605 196.135 32.865 196.525 ;
        RECT 33.055 197.345 34.020 197.355 ;
        RECT 34.190 197.435 34.360 197.815 ;
        RECT 34.950 197.775 35.120 198.065 ;
        RECT 35.300 197.945 35.630 198.325 ;
        RECT 34.950 197.605 35.750 197.775 ;
        RECT 33.055 197.185 33.730 197.345 ;
        RECT 34.190 197.265 35.410 197.435 ;
        RECT 33.055 196.395 33.265 197.185 ;
        RECT 34.190 197.175 34.360 197.265 ;
        RECT 33.435 196.395 33.785 197.015 ;
        RECT 33.955 197.005 34.360 197.175 ;
        RECT 33.955 196.225 34.125 197.005 ;
        RECT 34.295 196.555 34.515 196.835 ;
        RECT 34.695 196.725 35.235 197.095 ;
        RECT 35.580 197.015 35.750 197.605 ;
        RECT 35.970 197.185 36.275 198.325 ;
        RECT 36.445 197.135 36.700 198.015 ;
        RECT 35.580 196.985 36.320 197.015 ;
        RECT 34.295 196.385 34.825 196.555 ;
        RECT 32.605 195.965 32.955 196.135 ;
        RECT 33.175 195.945 34.125 196.225 ;
        RECT 34.295 195.775 34.485 196.215 ;
        RECT 34.655 196.155 34.825 196.385 ;
        RECT 34.995 196.325 35.235 196.725 ;
        RECT 35.405 196.685 36.320 196.985 ;
        RECT 35.405 196.510 35.730 196.685 ;
        RECT 35.405 196.155 35.725 196.510 ;
        RECT 36.490 196.485 36.700 197.135 ;
        RECT 36.875 197.565 37.390 197.975 ;
        RECT 37.625 197.565 37.795 198.325 ;
        RECT 37.965 197.985 39.995 198.155 ;
        RECT 36.875 196.755 37.215 197.565 ;
        RECT 37.965 197.320 38.135 197.985 ;
        RECT 38.530 197.645 39.655 197.815 ;
        RECT 37.385 197.130 38.135 197.320 ;
        RECT 38.305 197.305 39.315 197.475 ;
        RECT 36.875 196.585 38.105 196.755 ;
        RECT 34.655 195.985 35.725 196.155 ;
        RECT 35.970 195.775 36.275 196.235 ;
        RECT 36.445 195.955 36.700 196.485 ;
        RECT 37.150 195.980 37.395 196.585 ;
        RECT 37.615 195.775 38.125 196.310 ;
        RECT 38.305 195.945 38.495 197.305 ;
        RECT 38.665 196.285 38.940 197.105 ;
        RECT 39.145 196.505 39.315 197.305 ;
        RECT 39.485 196.515 39.655 197.645 ;
        RECT 39.825 197.015 39.995 197.985 ;
        RECT 40.165 197.185 40.335 198.325 ;
        RECT 40.505 197.185 40.840 198.155 ;
        RECT 39.825 196.685 40.020 197.015 ;
        RECT 40.245 196.685 40.500 197.015 ;
        RECT 40.245 196.515 40.415 196.685 ;
        RECT 40.670 196.515 40.840 197.185 ;
        RECT 41.475 197.160 41.765 198.325 ;
        RECT 42.120 197.355 42.510 197.530 ;
        RECT 42.995 197.525 43.325 198.325 ;
        RECT 43.495 197.535 44.030 198.155 ;
        RECT 42.120 197.185 43.545 197.355 ;
        RECT 39.485 196.345 40.415 196.515 ;
        RECT 39.485 196.310 39.660 196.345 ;
        RECT 38.665 196.115 38.945 196.285 ;
        RECT 38.665 195.945 38.940 196.115 ;
        RECT 39.130 195.945 39.660 196.310 ;
        RECT 40.085 195.775 40.415 196.175 ;
        RECT 40.585 195.945 40.840 196.515 ;
        RECT 41.475 195.775 41.765 196.500 ;
        RECT 41.995 196.455 42.350 197.015 ;
        RECT 42.520 196.285 42.690 197.185 ;
        RECT 42.860 196.455 43.125 197.015 ;
        RECT 43.375 196.685 43.545 197.185 ;
        RECT 43.715 196.515 44.030 197.535 ;
        RECT 42.100 195.775 42.340 196.285 ;
        RECT 42.520 195.955 42.800 196.285 ;
        RECT 43.030 195.775 43.245 196.285 ;
        RECT 43.415 195.945 44.030 196.515 ;
        RECT 44.235 197.565 44.900 198.155 ;
        RECT 44.235 196.595 44.485 197.565 ;
        RECT 45.070 197.485 45.400 198.325 ;
        RECT 45.910 197.735 46.715 198.155 ;
        RECT 45.570 197.565 47.135 197.735 ;
        RECT 45.570 197.315 45.740 197.565 ;
        RECT 44.820 197.145 45.740 197.315 ;
        RECT 45.910 197.305 46.285 197.395 ;
        RECT 44.820 196.975 44.990 197.145 ;
        RECT 45.910 197.135 46.305 197.305 ;
        RECT 45.910 196.975 46.285 197.135 ;
        RECT 44.655 196.765 44.990 196.975 ;
        RECT 45.160 196.765 45.610 196.975 ;
        RECT 45.800 196.765 46.285 196.975 ;
        RECT 46.475 197.015 46.795 197.395 ;
        RECT 46.965 197.315 47.135 197.565 ;
        RECT 47.305 197.485 47.555 198.325 ;
        RECT 47.750 197.315 48.050 198.155 ;
        RECT 46.965 197.145 48.050 197.315 ;
        RECT 48.375 197.565 49.040 198.155 ;
        RECT 46.475 196.765 46.855 197.015 ;
        RECT 47.035 196.765 47.365 196.975 ;
        RECT 44.235 195.955 44.920 196.595 ;
        RECT 45.090 195.775 45.260 196.595 ;
        RECT 45.430 196.425 47.130 196.595 ;
        RECT 45.430 195.960 45.760 196.425 ;
        RECT 46.745 196.335 47.130 196.425 ;
        RECT 47.535 196.515 47.705 197.145 ;
        RECT 47.875 196.685 48.205 196.975 ;
        RECT 48.375 196.595 48.625 197.565 ;
        RECT 49.210 197.485 49.540 198.325 ;
        RECT 50.050 197.735 50.855 198.155 ;
        RECT 49.710 197.565 51.275 197.735 ;
        RECT 49.710 197.315 49.880 197.565 ;
        RECT 48.960 197.145 49.880 197.315 ;
        RECT 48.960 196.975 49.130 197.145 ;
        RECT 50.050 196.975 50.425 197.395 ;
        RECT 48.795 196.765 49.130 196.975 ;
        RECT 49.300 196.765 49.750 196.975 ;
        RECT 49.940 196.965 50.425 196.975 ;
        RECT 50.615 197.015 50.935 197.395 ;
        RECT 51.105 197.315 51.275 197.565 ;
        RECT 51.445 197.485 51.695 198.325 ;
        RECT 51.890 197.315 52.190 198.155 ;
        RECT 51.105 197.145 52.190 197.315 ;
        RECT 52.550 197.535 53.085 198.155 ;
        RECT 49.940 196.795 50.445 196.965 ;
        RECT 49.940 196.765 50.425 196.795 ;
        RECT 50.615 196.765 50.995 197.015 ;
        RECT 51.175 196.765 51.505 196.975 ;
        RECT 47.535 196.335 48.045 196.515 ;
        RECT 45.930 195.775 46.100 196.245 ;
        RECT 46.360 195.995 47.545 196.165 ;
        RECT 47.715 195.945 48.045 196.335 ;
        RECT 48.375 195.955 49.060 196.595 ;
        RECT 49.230 195.775 49.400 196.595 ;
        RECT 49.570 196.425 51.270 196.595 ;
        RECT 49.570 195.960 49.900 196.425 ;
        RECT 50.885 196.335 51.270 196.425 ;
        RECT 51.675 196.515 51.845 197.145 ;
        RECT 52.015 196.685 52.345 196.975 ;
        RECT 52.550 196.515 52.865 197.535 ;
        RECT 53.255 197.525 53.585 198.325 ;
        RECT 54.850 197.535 55.385 198.155 ;
        RECT 54.070 197.355 54.460 197.530 ;
        RECT 53.035 197.185 54.460 197.355 ;
        RECT 53.035 196.685 53.205 197.185 ;
        RECT 51.675 196.335 52.185 196.515 ;
        RECT 50.070 195.775 50.240 196.245 ;
        RECT 50.500 195.995 51.685 196.165 ;
        RECT 51.855 195.945 52.185 196.335 ;
        RECT 52.550 195.945 53.165 196.515 ;
        RECT 53.455 196.455 53.720 197.015 ;
        RECT 53.890 196.285 54.060 197.185 ;
        RECT 54.230 196.455 54.585 197.015 ;
        RECT 54.850 196.515 55.165 197.535 ;
        RECT 55.555 197.525 55.885 198.325 ;
        RECT 56.370 197.355 56.760 197.530 ;
        RECT 55.335 197.185 56.760 197.355 ;
        RECT 55.335 196.685 55.505 197.185 ;
        RECT 53.335 195.775 53.550 196.285 ;
        RECT 53.780 195.955 54.060 196.285 ;
        RECT 54.240 195.775 54.480 196.285 ;
        RECT 54.850 195.945 55.465 196.515 ;
        RECT 55.755 196.455 56.020 197.015 ;
        RECT 56.190 196.285 56.360 197.185 ;
        RECT 57.120 197.175 57.380 198.325 ;
        RECT 57.555 197.250 57.810 198.155 ;
        RECT 57.980 197.565 58.310 198.325 ;
        RECT 58.525 197.395 58.695 198.155 ;
        RECT 56.530 196.455 56.885 197.015 ;
        RECT 55.635 195.775 55.850 196.285 ;
        RECT 56.080 195.955 56.360 196.285 ;
        RECT 56.540 195.775 56.780 196.285 ;
        RECT 57.120 195.775 57.380 196.615 ;
        RECT 57.555 196.520 57.725 197.250 ;
        RECT 57.980 197.225 58.695 197.395 ;
        RECT 57.980 197.015 58.150 197.225 ;
        RECT 57.895 196.685 58.150 197.015 ;
        RECT 57.555 195.945 57.810 196.520 ;
        RECT 57.980 196.495 58.150 196.685 ;
        RECT 58.430 196.675 58.785 197.045 ;
        RECT 57.980 196.325 58.695 196.495 ;
        RECT 57.980 195.775 58.310 196.155 ;
        RECT 58.525 195.945 58.695 196.325 ;
        RECT 59.885 195.955 60.145 198.145 ;
        RECT 60.315 197.595 60.655 198.325 ;
        RECT 60.835 197.415 61.105 198.145 ;
        RECT 60.335 197.195 61.105 197.415 ;
        RECT 61.285 197.435 61.515 198.145 ;
        RECT 61.685 197.615 62.015 198.325 ;
        RECT 62.185 197.435 62.445 198.145 ;
        RECT 61.285 197.195 62.445 197.435 ;
        RECT 62.635 197.475 62.975 198.115 ;
        RECT 63.145 197.865 63.390 198.325 ;
        RECT 63.565 197.695 63.815 198.155 ;
        RECT 64.005 197.945 64.675 198.325 ;
        RECT 64.875 197.695 65.125 198.155 ;
        RECT 63.565 197.525 65.125 197.695 ;
        RECT 60.335 196.525 60.625 197.195 ;
        RECT 60.805 196.705 61.270 197.015 ;
        RECT 61.450 196.705 61.975 197.015 ;
        RECT 60.335 196.325 61.565 196.525 ;
        RECT 60.405 195.775 61.075 196.145 ;
        RECT 61.255 195.955 61.565 196.325 ;
        RECT 61.745 196.065 61.975 196.705 ;
        RECT 62.155 196.685 62.455 197.015 ;
        RECT 62.155 195.775 62.445 196.505 ;
        RECT 62.635 196.360 62.805 197.475 ;
        RECT 65.885 197.355 66.055 198.155 ;
        RECT 63.115 197.185 66.055 197.355 ;
        RECT 63.115 197.015 63.285 197.185 ;
        RECT 67.235 197.160 67.525 198.325 ;
        RECT 68.705 197.315 68.875 198.155 ;
        RECT 69.045 197.985 70.215 198.155 ;
        RECT 69.045 197.485 69.375 197.985 ;
        RECT 69.885 197.945 70.215 197.985 ;
        RECT 70.405 197.905 70.760 198.325 ;
        RECT 69.545 197.725 69.775 197.815 ;
        RECT 70.930 197.725 71.180 198.155 ;
        RECT 69.545 197.485 71.180 197.725 ;
        RECT 71.350 197.565 71.680 198.325 ;
        RECT 71.850 197.485 72.105 198.155 ;
        RECT 68.705 197.145 71.765 197.315 ;
        RECT 62.975 196.685 63.285 197.015 ;
        RECT 63.455 196.685 63.790 197.015 ;
        RECT 63.115 196.515 63.285 196.685 ;
        RECT 62.635 195.945 62.945 196.360 ;
        RECT 63.115 196.345 63.810 196.515 ;
        RECT 64.060 196.440 64.255 197.015 ;
        RECT 64.515 196.685 64.860 197.015 ;
        RECT 65.170 196.685 65.645 197.015 ;
        RECT 65.900 196.685 66.085 197.015 ;
        RECT 68.620 196.765 68.970 196.975 ;
        RECT 69.140 196.765 69.585 196.965 ;
        RECT 69.755 196.765 70.230 196.965 ;
        RECT 64.515 196.455 64.705 196.685 ;
        RECT 63.140 195.775 63.470 196.155 ;
        RECT 63.640 196.115 63.810 196.345 ;
        RECT 64.875 196.345 66.055 196.515 ;
        RECT 64.875 196.115 65.045 196.345 ;
        RECT 63.640 195.945 65.045 196.115 ;
        RECT 65.315 195.775 65.645 196.175 ;
        RECT 65.885 195.945 66.055 196.345 ;
        RECT 67.235 195.775 67.525 196.500 ;
        RECT 68.705 196.425 69.770 196.595 ;
        RECT 68.705 195.945 68.875 196.425 ;
        RECT 69.045 195.775 69.375 196.255 ;
        RECT 69.600 196.195 69.770 196.425 ;
        RECT 69.950 196.365 70.230 196.765 ;
        RECT 70.500 196.765 70.830 196.965 ;
        RECT 71.000 196.795 71.375 196.965 ;
        RECT 71.000 196.765 71.365 196.795 ;
        RECT 70.500 196.365 70.785 196.765 ;
        RECT 71.595 196.595 71.765 197.145 ;
        RECT 70.965 196.425 71.765 196.595 ;
        RECT 70.965 196.195 71.135 196.425 ;
        RECT 71.935 196.355 72.105 197.485 ;
        RECT 71.920 196.275 72.105 196.355 ;
        RECT 69.600 195.945 71.135 196.195 ;
        RECT 71.305 195.775 71.635 196.255 ;
        RECT 71.850 195.945 72.105 196.275 ;
        RECT 72.305 195.955 72.565 198.145 ;
        RECT 72.735 197.595 73.075 198.325 ;
        RECT 73.255 197.415 73.525 198.145 ;
        RECT 72.755 197.195 73.525 197.415 ;
        RECT 73.705 197.435 73.935 198.145 ;
        RECT 74.105 197.615 74.435 198.325 ;
        RECT 74.605 197.435 74.865 198.145 ;
        RECT 73.705 197.195 74.865 197.435 ;
        RECT 75.055 197.235 76.725 198.325 ;
        RECT 72.755 196.525 73.045 197.195 ;
        RECT 73.225 196.705 73.690 197.015 ;
        RECT 73.870 196.705 74.395 197.015 ;
        RECT 72.755 196.325 73.985 196.525 ;
        RECT 72.825 195.775 73.495 196.145 ;
        RECT 73.675 195.955 73.985 196.325 ;
        RECT 74.165 196.065 74.395 196.705 ;
        RECT 74.575 196.685 74.875 197.015 ;
        RECT 75.055 196.545 75.805 197.065 ;
        RECT 75.975 196.715 76.725 197.235 ;
        RECT 77.560 197.355 77.890 198.155 ;
        RECT 78.060 197.525 78.390 198.325 ;
        RECT 78.690 197.355 79.020 198.155 ;
        RECT 79.665 197.525 79.915 198.325 ;
        RECT 77.560 197.185 79.995 197.355 ;
        RECT 80.185 197.185 80.355 198.325 ;
        RECT 80.525 197.185 80.865 198.155 ;
        RECT 81.035 197.235 84.545 198.325 ;
        RECT 77.355 196.765 77.705 197.015 ;
        RECT 77.890 196.555 78.060 197.185 ;
        RECT 78.230 196.765 78.560 196.965 ;
        RECT 78.730 196.765 79.060 196.965 ;
        RECT 79.230 196.795 79.655 196.965 ;
        RECT 79.825 196.935 79.995 197.185 ;
        RECT 79.230 196.765 79.650 196.795 ;
        RECT 79.825 196.765 80.520 196.935 ;
        RECT 74.575 195.775 74.865 196.505 ;
        RECT 75.055 195.775 76.725 196.545 ;
        RECT 77.560 195.945 78.060 196.555 ;
        RECT 78.690 196.425 79.915 196.595 ;
        RECT 80.690 196.575 80.865 197.185 ;
        RECT 78.690 195.945 79.020 196.425 ;
        RECT 79.190 195.775 79.415 196.235 ;
        RECT 79.585 195.945 79.915 196.425 ;
        RECT 80.105 195.775 80.355 196.575 ;
        RECT 80.525 195.945 80.865 196.575 ;
        RECT 81.035 196.545 82.685 197.065 ;
        RECT 82.855 196.715 84.545 197.235 ;
        RECT 85.185 197.265 85.515 198.115 ;
        RECT 81.035 195.775 84.545 196.545 ;
        RECT 85.185 196.500 85.375 197.265 ;
        RECT 85.685 197.185 85.935 198.325 ;
        RECT 86.125 197.685 86.375 198.105 ;
        RECT 86.605 197.855 86.935 198.325 ;
        RECT 87.165 197.685 87.415 198.105 ;
        RECT 86.125 197.515 87.415 197.685 ;
        RECT 87.595 197.685 87.925 198.115 ;
        RECT 87.595 197.515 88.050 197.685 ;
        RECT 86.115 197.015 86.330 197.345 ;
        RECT 85.545 196.685 85.855 197.015 ;
        RECT 86.025 196.685 86.330 197.015 ;
        RECT 86.505 196.685 86.790 197.345 ;
        RECT 86.985 196.685 87.250 197.345 ;
        RECT 87.465 196.685 87.710 197.345 ;
        RECT 85.685 196.515 85.855 196.685 ;
        RECT 87.880 196.515 88.050 197.515 ;
        RECT 88.395 197.235 89.605 198.325 ;
        RECT 85.185 195.990 85.515 196.500 ;
        RECT 85.685 196.345 88.050 196.515 ;
        RECT 88.395 196.525 88.915 197.065 ;
        RECT 89.085 196.695 89.605 197.235 ;
        RECT 89.780 197.355 90.055 198.155 ;
        RECT 90.225 197.525 90.555 198.325 ;
        RECT 90.725 197.985 91.865 198.155 ;
        RECT 90.725 197.355 90.895 197.985 ;
        RECT 89.780 197.145 90.895 197.355 ;
        RECT 91.065 197.355 91.395 197.815 ;
        RECT 91.565 197.525 91.865 197.985 ;
        RECT 91.065 197.135 91.825 197.355 ;
        RECT 92.995 197.160 93.285 198.325 ;
        RECT 93.455 197.185 93.735 198.325 ;
        RECT 93.905 197.175 94.235 198.155 ;
        RECT 94.405 197.185 94.665 198.325 ;
        RECT 95.295 197.455 95.570 198.155 ;
        RECT 95.740 197.780 95.995 198.325 ;
        RECT 96.165 197.815 96.645 198.155 ;
        RECT 96.820 197.770 97.425 198.325 ;
        RECT 97.595 197.890 102.940 198.325 ;
        RECT 96.810 197.670 97.425 197.770 ;
        RECT 96.810 197.645 96.995 197.670 ;
        RECT 89.780 196.765 90.500 196.965 ;
        RECT 90.670 196.765 91.440 196.965 ;
        RECT 91.610 196.595 91.825 197.135 ;
        RECT 93.970 197.135 94.145 197.175 ;
        RECT 93.465 196.745 93.800 197.015 ;
        RECT 85.685 195.775 86.015 196.175 ;
        RECT 87.065 196.005 87.395 196.345 ;
        RECT 87.565 195.775 87.895 196.175 ;
        RECT 88.395 195.775 89.605 196.525 ;
        RECT 89.780 195.775 90.055 196.595 ;
        RECT 90.225 196.425 91.825 196.595 ;
        RECT 93.970 196.575 94.140 197.135 ;
        RECT 94.310 196.765 94.645 197.015 ;
        RECT 90.225 196.415 91.395 196.425 ;
        RECT 90.225 195.945 90.555 196.415 ;
        RECT 90.725 195.775 90.895 196.245 ;
        RECT 91.065 195.945 91.395 196.415 ;
        RECT 91.565 195.775 91.855 196.245 ;
        RECT 92.995 195.775 93.285 196.500 ;
        RECT 93.455 195.775 93.765 196.575 ;
        RECT 93.970 195.945 94.665 196.575 ;
        RECT 95.295 196.425 95.465 197.455 ;
        RECT 95.740 197.325 96.495 197.575 ;
        RECT 96.665 197.400 96.995 197.645 ;
        RECT 95.740 197.290 96.510 197.325 ;
        RECT 95.740 197.280 96.525 197.290 ;
        RECT 95.635 197.265 96.530 197.280 ;
        RECT 95.635 197.250 96.550 197.265 ;
        RECT 95.635 197.240 96.570 197.250 ;
        RECT 95.635 197.230 96.595 197.240 ;
        RECT 95.635 197.200 96.665 197.230 ;
        RECT 95.635 197.170 96.685 197.200 ;
        RECT 95.635 197.140 96.705 197.170 ;
        RECT 95.635 197.115 96.735 197.140 ;
        RECT 95.635 197.080 96.770 197.115 ;
        RECT 95.635 197.075 96.800 197.080 ;
        RECT 95.635 196.680 95.865 197.075 ;
        RECT 96.410 197.070 96.800 197.075 ;
        RECT 96.435 197.060 96.800 197.070 ;
        RECT 96.450 197.055 96.800 197.060 ;
        RECT 96.465 197.050 96.800 197.055 ;
        RECT 97.165 197.050 97.425 197.500 ;
        RECT 96.465 197.045 97.425 197.050 ;
        RECT 96.475 197.035 97.425 197.045 ;
        RECT 96.485 197.030 97.425 197.035 ;
        RECT 96.495 197.020 97.425 197.030 ;
        RECT 96.500 197.010 97.425 197.020 ;
        RECT 96.505 197.005 97.425 197.010 ;
        RECT 96.515 196.990 97.425 197.005 ;
        RECT 96.520 196.975 97.425 196.990 ;
        RECT 96.530 196.950 97.425 196.975 ;
        RECT 96.035 196.480 96.365 196.905 ;
        RECT 95.295 195.945 95.555 196.425 ;
        RECT 95.725 195.775 95.975 196.315 ;
        RECT 96.145 195.995 96.365 196.480 ;
        RECT 96.535 196.880 97.425 196.950 ;
        RECT 96.535 196.155 96.705 196.880 ;
        RECT 96.875 196.325 97.425 196.710 ;
        RECT 99.180 196.320 99.520 197.150 ;
        RECT 101.000 196.640 101.350 197.890 ;
        RECT 103.580 197.185 103.900 198.325 ;
        RECT 104.080 197.015 104.275 198.065 ;
        RECT 104.455 197.475 104.785 198.155 ;
        RECT 104.985 197.525 105.240 198.325 ;
        RECT 105.465 197.865 105.715 198.325 ;
        RECT 105.925 197.695 106.095 198.155 ;
        RECT 105.420 197.525 106.095 197.695 ;
        RECT 106.265 197.525 106.515 198.325 ;
        RECT 106.685 197.695 106.935 198.115 ;
        RECT 107.145 197.865 107.475 198.325 ;
        RECT 107.665 197.695 107.915 198.115 ;
        RECT 106.685 197.525 107.975 197.695 ;
        RECT 104.455 197.195 104.805 197.475 ;
        RECT 103.640 196.965 103.900 197.015 ;
        RECT 103.635 196.795 103.900 196.965 ;
        RECT 103.640 196.685 103.900 196.795 ;
        RECT 104.080 196.685 104.465 197.015 ;
        RECT 104.635 196.815 104.805 197.195 ;
        RECT 104.995 196.985 105.240 197.345 ;
        RECT 104.635 196.645 105.155 196.815 ;
        RECT 96.535 195.985 97.425 196.155 ;
        RECT 97.595 195.775 102.940 196.320 ;
        RECT 103.580 196.305 104.795 196.475 ;
        RECT 103.580 195.955 103.870 196.305 ;
        RECT 104.065 195.775 104.395 196.135 ;
        RECT 104.565 196.000 104.795 196.305 ;
        RECT 104.985 196.080 105.155 196.645 ;
        RECT 105.420 196.575 105.675 197.525 ;
        RECT 108.205 197.355 108.375 198.155 ;
        RECT 105.885 197.185 108.375 197.355 ;
        RECT 109.555 197.525 109.995 198.155 ;
        RECT 105.885 196.935 106.055 197.185 ;
        RECT 105.885 196.765 106.215 196.935 ;
        RECT 106.395 196.685 106.725 197.015 ;
        RECT 106.955 196.935 107.125 196.950 ;
        RECT 106.955 196.765 107.285 196.935 ;
        RECT 105.420 196.405 106.095 196.575 ;
        RECT 106.395 196.450 106.600 196.685 ;
        RECT 106.955 196.555 107.125 196.765 ;
        RECT 107.515 196.560 107.685 197.015 ;
        RECT 105.420 195.775 105.675 196.235 ;
        RECT 105.925 195.945 106.095 196.405 ;
        RECT 106.860 196.385 107.125 196.555 ;
        RECT 107.295 196.390 107.685 196.560 ;
        RECT 106.860 196.285 107.030 196.385 ;
        RECT 106.345 196.155 106.515 196.235 ;
        RECT 106.285 195.775 106.615 196.155 ;
        RECT 106.855 196.115 107.030 196.285 ;
        RECT 106.860 196.090 107.030 196.115 ;
        RECT 107.295 196.105 107.505 196.390 ;
        RECT 107.865 196.195 108.035 197.185 ;
        RECT 108.225 196.445 108.420 197.015 ;
        RECT 109.555 196.515 109.865 197.525 ;
        RECT 110.170 197.475 110.485 198.325 ;
        RECT 110.655 197.985 112.085 198.155 ;
        RECT 110.655 197.305 110.825 197.985 ;
        RECT 110.035 197.135 110.825 197.305 ;
        RECT 110.035 196.685 110.205 197.135 ;
        RECT 110.995 197.015 111.195 197.815 ;
        RECT 110.375 196.685 110.765 196.965 ;
        RECT 110.950 196.685 111.195 197.015 ;
        RECT 111.395 196.685 111.645 197.815 ;
        RECT 111.835 197.355 112.085 197.985 ;
        RECT 112.265 197.525 112.595 198.325 ;
        RECT 112.775 197.890 118.120 198.325 ;
        RECT 111.835 197.185 112.605 197.355 ;
        RECT 111.860 196.685 112.265 197.015 ;
        RECT 112.435 196.515 112.605 197.185 ;
        RECT 107.705 196.025 108.035 196.195 ;
        RECT 107.790 195.945 108.035 196.025 ;
        RECT 108.205 195.775 108.465 196.255 ;
        RECT 109.555 195.955 109.995 196.515 ;
        RECT 110.165 195.775 110.615 196.515 ;
        RECT 110.785 196.345 111.945 196.515 ;
        RECT 110.785 195.945 110.955 196.345 ;
        RECT 111.125 195.775 111.545 196.175 ;
        RECT 111.715 195.945 111.945 196.345 ;
        RECT 112.115 195.945 112.605 196.515 ;
        RECT 114.360 196.320 114.700 197.150 ;
        RECT 116.180 196.640 116.530 197.890 ;
        RECT 118.755 197.160 119.045 198.325 ;
        RECT 119.215 197.890 124.560 198.325 ;
        RECT 112.775 195.775 118.120 196.320 ;
        RECT 118.755 195.775 119.045 196.500 ;
        RECT 120.800 196.320 121.140 197.150 ;
        RECT 122.620 196.640 122.970 197.890 ;
        RECT 125.195 197.355 125.505 198.155 ;
        RECT 125.675 197.525 125.985 198.325 ;
        RECT 126.155 197.695 126.415 198.155 ;
        RECT 126.585 197.865 126.840 198.325 ;
        RECT 127.015 197.695 127.275 198.155 ;
        RECT 126.155 197.525 127.275 197.695 ;
        RECT 126.635 197.475 126.805 197.525 ;
        RECT 125.195 197.185 126.225 197.355 ;
        RECT 119.215 195.775 124.560 196.320 ;
        RECT 125.195 196.275 125.365 197.185 ;
        RECT 125.535 196.445 125.885 197.015 ;
        RECT 126.055 196.935 126.225 197.185 ;
        RECT 127.015 197.275 127.275 197.525 ;
        RECT 127.445 197.455 127.730 198.325 ;
        RECT 127.015 197.105 127.770 197.275 ;
        RECT 127.955 197.235 131.465 198.325 ;
        RECT 126.055 196.765 127.195 196.935 ;
        RECT 127.365 196.595 127.770 197.105 ;
        RECT 126.120 196.425 127.770 196.595 ;
        RECT 127.955 196.545 129.605 197.065 ;
        RECT 129.775 196.715 131.465 197.235 ;
        RECT 132.185 197.355 132.355 198.155 ;
        RECT 133.115 197.695 133.365 198.155 ;
        RECT 133.565 197.945 134.235 198.325 ;
        RECT 134.425 197.695 134.675 198.155 ;
        RECT 134.850 197.865 135.095 198.325 ;
        RECT 133.115 197.525 134.675 197.695 ;
        RECT 135.265 197.475 135.605 198.115 ;
        RECT 132.185 197.185 135.125 197.355 ;
        RECT 134.955 197.015 135.125 197.185 ;
        RECT 132.155 196.685 132.340 197.015 ;
        RECT 132.595 196.685 133.070 197.015 ;
        RECT 133.380 196.685 133.725 197.015 ;
        RECT 125.195 195.945 125.495 196.275 ;
        RECT 125.665 195.775 125.940 196.255 ;
        RECT 126.120 196.035 126.415 196.425 ;
        RECT 126.585 195.775 126.840 196.255 ;
        RECT 127.015 196.035 127.275 196.425 ;
        RECT 127.445 195.775 127.725 196.255 ;
        RECT 127.955 195.775 131.465 196.545 ;
        RECT 132.185 196.345 133.365 196.515 ;
        RECT 133.535 196.455 133.725 196.685 ;
        RECT 133.985 196.440 134.180 197.015 ;
        RECT 134.450 196.685 134.785 197.015 ;
        RECT 134.955 196.685 135.265 197.015 ;
        RECT 134.955 196.515 135.125 196.685 ;
        RECT 132.185 195.945 132.355 196.345 ;
        RECT 132.595 195.775 132.925 196.175 ;
        RECT 133.195 196.115 133.365 196.345 ;
        RECT 134.430 196.345 135.125 196.515 ;
        RECT 135.435 196.360 135.605 197.475 ;
        RECT 136.275 197.375 136.565 198.145 ;
        RECT 137.135 197.785 137.395 198.145 ;
        RECT 137.565 197.955 137.895 198.325 ;
        RECT 138.065 197.785 138.325 198.145 ;
        RECT 137.135 197.555 138.325 197.785 ;
        RECT 138.515 197.605 138.845 198.325 ;
        RECT 139.015 197.375 139.280 198.145 ;
        RECT 136.275 197.195 138.770 197.375 ;
        RECT 136.245 196.685 136.515 197.015 ;
        RECT 136.695 196.685 137.130 197.015 ;
        RECT 137.310 196.685 137.885 197.015 ;
        RECT 138.065 196.685 138.345 197.015 ;
        RECT 138.545 196.505 138.770 197.195 ;
        RECT 134.430 196.115 134.600 196.345 ;
        RECT 133.195 195.945 134.600 196.115 ;
        RECT 134.770 195.775 135.100 196.155 ;
        RECT 135.295 195.945 135.605 196.360 ;
        RECT 136.285 196.315 138.770 196.505 ;
        RECT 136.285 195.955 136.510 196.315 ;
        RECT 136.690 195.775 137.020 196.145 ;
        RECT 137.200 195.955 137.455 196.315 ;
        RECT 138.020 195.775 138.765 196.145 ;
        RECT 138.945 195.955 139.280 197.375 ;
        RECT 139.455 197.185 139.735 198.325 ;
        RECT 139.905 197.175 140.235 198.155 ;
        RECT 140.405 197.185 140.665 198.325 ;
        RECT 140.835 197.235 144.345 198.325 ;
        RECT 139.465 196.745 139.800 197.015 ;
        RECT 139.970 196.625 140.140 197.175 ;
        RECT 140.310 196.765 140.645 197.015 ;
        RECT 139.970 196.575 140.145 196.625 ;
        RECT 139.455 195.775 139.765 196.575 ;
        RECT 139.970 195.945 140.665 196.575 ;
        RECT 140.835 196.545 142.485 197.065 ;
        RECT 142.655 196.715 144.345 197.235 ;
        RECT 144.515 197.160 144.805 198.325 ;
        RECT 144.975 197.890 150.320 198.325 ;
        RECT 140.835 195.775 144.345 196.545 ;
        RECT 144.515 195.775 144.805 196.500 ;
        RECT 146.560 196.320 146.900 197.150 ;
        RECT 148.380 196.640 148.730 197.890 ;
        RECT 150.585 197.315 150.755 198.155 ;
        RECT 150.925 197.985 152.095 198.155 ;
        RECT 150.925 197.485 151.255 197.985 ;
        RECT 151.765 197.945 152.095 197.985 ;
        RECT 152.285 197.905 152.640 198.325 ;
        RECT 151.425 197.725 151.655 197.815 ;
        RECT 152.810 197.725 153.060 198.155 ;
        RECT 151.425 197.485 153.060 197.725 ;
        RECT 153.230 197.565 153.560 198.325 ;
        RECT 153.730 197.485 153.985 198.155 ;
        RECT 150.585 197.145 153.645 197.315 ;
        RECT 150.500 196.765 150.850 196.975 ;
        RECT 151.020 196.765 151.465 196.965 ;
        RECT 151.635 196.765 152.110 196.965 ;
        RECT 150.585 196.425 151.650 196.595 ;
        RECT 144.975 195.775 150.320 196.320 ;
        RECT 150.585 195.945 150.755 196.425 ;
        RECT 150.925 195.775 151.255 196.255 ;
        RECT 151.480 196.195 151.650 196.425 ;
        RECT 151.830 196.365 152.110 196.765 ;
        RECT 152.380 196.765 152.710 196.965 ;
        RECT 152.880 196.765 153.245 196.965 ;
        RECT 152.380 196.365 152.665 196.765 ;
        RECT 153.475 196.595 153.645 197.145 ;
        RECT 152.845 196.425 153.645 196.595 ;
        RECT 152.845 196.195 153.015 196.425 ;
        RECT 153.815 196.355 153.985 197.485 ;
        RECT 154.175 197.235 156.765 198.325 ;
        RECT 153.800 196.275 153.985 196.355 ;
        RECT 151.480 195.945 153.015 196.195 ;
        RECT 153.185 195.775 153.515 196.255 ;
        RECT 153.730 195.945 153.985 196.275 ;
        RECT 154.175 196.545 155.385 197.065 ;
        RECT 155.555 196.715 156.765 197.235 ;
        RECT 156.935 197.235 158.145 198.325 ;
        RECT 156.935 196.695 157.455 197.235 ;
        RECT 154.175 195.775 156.765 196.545 ;
        RECT 157.625 196.525 158.145 197.065 ;
        RECT 156.935 195.775 158.145 196.525 ;
        RECT 2.750 195.605 158.230 195.775 ;
        RECT 2.835 194.855 4.045 195.605 ;
        RECT 4.220 195.055 4.475 195.345 ;
        RECT 4.645 195.225 4.975 195.605 ;
        RECT 4.220 194.885 4.970 195.055 ;
        RECT 2.835 194.315 3.355 194.855 ;
        RECT 3.525 194.145 4.045 194.685 ;
        RECT 2.835 193.055 4.045 194.145 ;
        RECT 4.220 194.065 4.570 194.715 ;
        RECT 4.740 193.895 4.970 194.885 ;
        RECT 4.220 193.725 4.970 193.895 ;
        RECT 4.220 193.225 4.475 193.725 ;
        RECT 4.645 193.055 4.975 193.555 ;
        RECT 5.145 193.225 5.315 195.345 ;
        RECT 5.675 195.245 6.005 195.605 ;
        RECT 6.175 195.215 6.670 195.385 ;
        RECT 6.875 195.215 7.730 195.385 ;
        RECT 5.545 194.025 6.005 195.075 ;
        RECT 5.485 193.240 5.810 194.025 ;
        RECT 6.175 193.855 6.345 195.215 ;
        RECT 6.515 194.305 6.865 194.925 ;
        RECT 7.035 194.705 7.390 194.925 ;
        RECT 7.035 194.115 7.205 194.705 ;
        RECT 7.560 194.505 7.730 195.215 ;
        RECT 8.605 195.145 8.935 195.605 ;
        RECT 9.145 195.245 9.495 195.415 ;
        RECT 7.935 194.675 8.725 194.925 ;
        RECT 9.145 194.855 9.405 195.245 ;
        RECT 9.715 195.155 10.665 195.435 ;
        RECT 10.835 195.165 11.025 195.605 ;
        RECT 11.195 195.225 12.265 195.395 ;
        RECT 8.895 194.505 9.065 194.685 ;
        RECT 6.175 193.685 6.570 193.855 ;
        RECT 6.740 193.725 7.205 194.115 ;
        RECT 7.375 194.335 9.065 194.505 ;
        RECT 6.400 193.555 6.570 193.685 ;
        RECT 7.375 193.555 7.545 194.335 ;
        RECT 9.235 194.165 9.405 194.855 ;
        RECT 7.905 193.995 9.405 194.165 ;
        RECT 9.595 194.195 9.805 194.985 ;
        RECT 9.975 194.365 10.325 194.985 ;
        RECT 10.495 194.375 10.665 195.155 ;
        RECT 11.195 194.995 11.365 195.225 ;
        RECT 10.835 194.825 11.365 194.995 ;
        RECT 10.835 194.545 11.055 194.825 ;
        RECT 11.535 194.655 11.775 195.055 ;
        RECT 10.495 194.205 10.900 194.375 ;
        RECT 11.235 194.285 11.775 194.655 ;
        RECT 11.945 194.870 12.265 195.225 ;
        RECT 12.510 195.145 12.815 195.605 ;
        RECT 12.985 194.895 13.240 195.425 ;
        RECT 11.945 194.695 12.270 194.870 ;
        RECT 11.945 194.395 12.860 194.695 ;
        RECT 12.120 194.365 12.860 194.395 ;
        RECT 9.595 194.035 10.270 194.195 ;
        RECT 10.730 194.115 10.900 194.205 ;
        RECT 9.595 194.025 10.560 194.035 ;
        RECT 9.235 193.855 9.405 193.995 ;
        RECT 5.980 193.055 6.230 193.515 ;
        RECT 6.400 193.225 6.650 193.555 ;
        RECT 6.865 193.225 7.545 193.555 ;
        RECT 7.715 193.655 8.790 193.825 ;
        RECT 9.235 193.685 9.795 193.855 ;
        RECT 10.100 193.735 10.560 194.025 ;
        RECT 10.730 193.945 11.950 194.115 ;
        RECT 7.715 193.315 7.885 193.655 ;
        RECT 8.120 193.055 8.450 193.485 ;
        RECT 8.620 193.315 8.790 193.655 ;
        RECT 9.085 193.055 9.455 193.515 ;
        RECT 9.625 193.225 9.795 193.685 ;
        RECT 10.730 193.565 10.900 193.945 ;
        RECT 12.120 193.775 12.290 194.365 ;
        RECT 13.030 194.245 13.240 194.895 ;
        RECT 13.415 194.835 15.085 195.605 ;
        RECT 15.260 195.055 15.515 195.345 ;
        RECT 15.685 195.225 16.015 195.605 ;
        RECT 15.260 194.885 16.010 195.055 ;
        RECT 13.415 194.315 14.165 194.835 ;
        RECT 10.030 193.225 10.900 193.565 ;
        RECT 11.490 193.605 12.290 193.775 ;
        RECT 11.070 193.055 11.320 193.515 ;
        RECT 11.490 193.315 11.660 193.605 ;
        RECT 11.840 193.055 12.170 193.435 ;
        RECT 12.510 193.055 12.815 194.195 ;
        RECT 12.985 193.365 13.240 194.245 ;
        RECT 14.335 194.145 15.085 194.665 ;
        RECT 13.415 193.055 15.085 194.145 ;
        RECT 15.260 194.065 15.610 194.715 ;
        RECT 15.780 193.895 16.010 194.885 ;
        RECT 15.260 193.725 16.010 193.895 ;
        RECT 15.260 193.225 15.515 193.725 ;
        RECT 15.685 193.055 16.015 193.555 ;
        RECT 16.185 193.225 16.355 195.345 ;
        RECT 16.715 195.245 17.045 195.605 ;
        RECT 17.215 195.215 17.710 195.385 ;
        RECT 17.915 195.215 18.770 195.385 ;
        RECT 16.585 194.025 17.045 195.075 ;
        RECT 16.525 193.240 16.850 194.025 ;
        RECT 17.215 193.855 17.385 195.215 ;
        RECT 17.555 194.305 17.905 194.925 ;
        RECT 18.075 194.705 18.430 194.925 ;
        RECT 18.075 194.115 18.245 194.705 ;
        RECT 18.600 194.505 18.770 195.215 ;
        RECT 19.645 195.145 19.975 195.605 ;
        RECT 20.185 195.245 20.535 195.415 ;
        RECT 18.975 194.675 19.765 194.925 ;
        RECT 20.185 194.855 20.445 195.245 ;
        RECT 20.755 195.155 21.705 195.435 ;
        RECT 21.875 195.165 22.065 195.605 ;
        RECT 22.235 195.225 23.305 195.395 ;
        RECT 19.935 194.505 20.105 194.685 ;
        RECT 17.215 193.685 17.610 193.855 ;
        RECT 17.780 193.725 18.245 194.115 ;
        RECT 18.415 194.335 20.105 194.505 ;
        RECT 17.440 193.555 17.610 193.685 ;
        RECT 18.415 193.555 18.585 194.335 ;
        RECT 20.275 194.165 20.445 194.855 ;
        RECT 18.945 193.995 20.445 194.165 ;
        RECT 20.635 194.195 20.845 194.985 ;
        RECT 21.015 194.365 21.365 194.985 ;
        RECT 21.535 194.375 21.705 195.155 ;
        RECT 22.235 194.995 22.405 195.225 ;
        RECT 21.875 194.825 22.405 194.995 ;
        RECT 21.875 194.545 22.095 194.825 ;
        RECT 22.575 194.655 22.815 195.055 ;
        RECT 21.535 194.205 21.940 194.375 ;
        RECT 22.275 194.285 22.815 194.655 ;
        RECT 22.985 194.870 23.305 195.225 ;
        RECT 23.550 195.145 23.855 195.605 ;
        RECT 24.025 194.895 24.280 195.425 ;
        RECT 24.515 195.125 24.795 195.605 ;
        RECT 24.965 194.955 25.225 195.345 ;
        RECT 25.400 195.125 25.655 195.605 ;
        RECT 25.825 194.955 26.120 195.345 ;
        RECT 26.300 195.125 26.575 195.605 ;
        RECT 26.745 195.105 27.045 195.435 ;
        RECT 22.985 194.695 23.310 194.870 ;
        RECT 22.985 194.395 23.900 194.695 ;
        RECT 23.160 194.365 23.900 194.395 ;
        RECT 20.635 194.035 21.310 194.195 ;
        RECT 21.770 194.115 21.940 194.205 ;
        RECT 20.635 194.025 21.600 194.035 ;
        RECT 20.275 193.855 20.445 193.995 ;
        RECT 17.020 193.055 17.270 193.515 ;
        RECT 17.440 193.225 17.690 193.555 ;
        RECT 17.905 193.225 18.585 193.555 ;
        RECT 18.755 193.655 19.830 193.825 ;
        RECT 20.275 193.685 20.835 193.855 ;
        RECT 21.140 193.735 21.600 194.025 ;
        RECT 21.770 193.945 22.990 194.115 ;
        RECT 18.755 193.315 18.925 193.655 ;
        RECT 19.160 193.055 19.490 193.485 ;
        RECT 19.660 193.315 19.830 193.655 ;
        RECT 20.125 193.055 20.495 193.515 ;
        RECT 20.665 193.225 20.835 193.685 ;
        RECT 21.770 193.565 21.940 193.945 ;
        RECT 23.160 193.775 23.330 194.365 ;
        RECT 24.070 194.245 24.280 194.895 ;
        RECT 21.070 193.225 21.940 193.565 ;
        RECT 22.530 193.605 23.330 193.775 ;
        RECT 22.110 193.055 22.360 193.515 ;
        RECT 22.530 193.315 22.700 193.605 ;
        RECT 22.880 193.055 23.210 193.435 ;
        RECT 23.550 193.055 23.855 194.195 ;
        RECT 24.025 193.365 24.280 194.245 ;
        RECT 24.470 194.785 26.120 194.955 ;
        RECT 24.470 194.275 24.875 194.785 ;
        RECT 25.045 194.445 26.185 194.615 ;
        RECT 24.470 194.105 25.225 194.275 ;
        RECT 24.510 193.055 24.795 193.925 ;
        RECT 24.965 193.855 25.225 194.105 ;
        RECT 26.015 194.195 26.185 194.445 ;
        RECT 26.355 194.365 26.705 194.935 ;
        RECT 26.875 194.195 27.045 195.105 ;
        RECT 27.305 195.055 27.475 195.435 ;
        RECT 27.655 195.225 27.985 195.605 ;
        RECT 27.305 194.885 27.970 195.055 ;
        RECT 28.165 194.930 28.425 195.435 ;
        RECT 27.235 194.335 27.565 194.705 ;
        RECT 27.800 194.630 27.970 194.885 ;
        RECT 26.015 194.025 27.045 194.195 ;
        RECT 27.800 194.300 28.085 194.630 ;
        RECT 27.800 194.155 27.970 194.300 ;
        RECT 24.965 193.685 26.085 193.855 ;
        RECT 24.965 193.225 25.225 193.685 ;
        RECT 25.400 193.055 25.655 193.515 ;
        RECT 25.825 193.225 26.085 193.685 ;
        RECT 26.255 193.055 26.565 193.855 ;
        RECT 26.735 193.225 27.045 194.025 ;
        RECT 27.305 193.985 27.970 194.155 ;
        RECT 28.255 194.130 28.425 194.930 ;
        RECT 28.595 194.880 28.885 195.605 ;
        RECT 29.060 195.055 29.315 195.345 ;
        RECT 29.485 195.225 29.815 195.605 ;
        RECT 29.060 194.885 29.810 195.055 ;
        RECT 27.305 193.225 27.475 193.985 ;
        RECT 27.655 193.055 27.985 193.815 ;
        RECT 28.155 193.225 28.425 194.130 ;
        RECT 28.595 193.055 28.885 194.220 ;
        RECT 29.060 194.065 29.410 194.715 ;
        RECT 29.580 193.895 29.810 194.885 ;
        RECT 29.060 193.725 29.810 193.895 ;
        RECT 29.060 193.225 29.315 193.725 ;
        RECT 29.485 193.055 29.815 193.555 ;
        RECT 29.985 193.225 30.155 195.345 ;
        RECT 30.515 195.245 30.845 195.605 ;
        RECT 31.015 195.215 31.510 195.385 ;
        RECT 31.715 195.215 32.570 195.385 ;
        RECT 30.385 194.025 30.845 195.075 ;
        RECT 30.325 193.240 30.650 194.025 ;
        RECT 31.015 193.855 31.185 195.215 ;
        RECT 31.355 194.305 31.705 194.925 ;
        RECT 31.875 194.705 32.230 194.925 ;
        RECT 31.875 194.115 32.045 194.705 ;
        RECT 32.400 194.505 32.570 195.215 ;
        RECT 33.445 195.145 33.775 195.605 ;
        RECT 33.985 195.245 34.335 195.415 ;
        RECT 32.775 194.675 33.565 194.925 ;
        RECT 33.985 194.855 34.245 195.245 ;
        RECT 34.555 195.155 35.505 195.435 ;
        RECT 35.675 195.165 35.865 195.605 ;
        RECT 36.035 195.225 37.105 195.395 ;
        RECT 33.735 194.505 33.905 194.685 ;
        RECT 31.015 193.685 31.410 193.855 ;
        RECT 31.580 193.725 32.045 194.115 ;
        RECT 32.215 194.335 33.905 194.505 ;
        RECT 31.240 193.555 31.410 193.685 ;
        RECT 32.215 193.555 32.385 194.335 ;
        RECT 34.075 194.165 34.245 194.855 ;
        RECT 32.745 193.995 34.245 194.165 ;
        RECT 34.435 194.195 34.645 194.985 ;
        RECT 34.815 194.365 35.165 194.985 ;
        RECT 35.335 194.375 35.505 195.155 ;
        RECT 36.035 194.995 36.205 195.225 ;
        RECT 35.675 194.825 36.205 194.995 ;
        RECT 35.675 194.545 35.895 194.825 ;
        RECT 36.375 194.655 36.615 195.055 ;
        RECT 35.335 194.205 35.740 194.375 ;
        RECT 36.075 194.285 36.615 194.655 ;
        RECT 36.785 194.870 37.105 195.225 ;
        RECT 37.350 195.145 37.655 195.605 ;
        RECT 37.825 194.895 38.080 195.425 ;
        RECT 36.785 194.695 37.110 194.870 ;
        RECT 36.785 194.395 37.700 194.695 ;
        RECT 36.960 194.365 37.700 194.395 ;
        RECT 34.435 194.035 35.110 194.195 ;
        RECT 35.570 194.115 35.740 194.205 ;
        RECT 34.435 194.025 35.400 194.035 ;
        RECT 34.075 193.855 34.245 193.995 ;
        RECT 30.820 193.055 31.070 193.515 ;
        RECT 31.240 193.225 31.490 193.555 ;
        RECT 31.705 193.225 32.385 193.555 ;
        RECT 32.555 193.655 33.630 193.825 ;
        RECT 34.075 193.685 34.635 193.855 ;
        RECT 34.940 193.735 35.400 194.025 ;
        RECT 35.570 193.945 36.790 194.115 ;
        RECT 32.555 193.315 32.725 193.655 ;
        RECT 32.960 193.055 33.290 193.485 ;
        RECT 33.460 193.315 33.630 193.655 ;
        RECT 33.925 193.055 34.295 193.515 ;
        RECT 34.465 193.225 34.635 193.685 ;
        RECT 35.570 193.565 35.740 193.945 ;
        RECT 36.960 193.775 37.130 194.365 ;
        RECT 37.870 194.245 38.080 194.895 ;
        RECT 34.870 193.225 35.740 193.565 ;
        RECT 36.330 193.605 37.130 193.775 ;
        RECT 35.910 193.055 36.160 193.515 ;
        RECT 36.330 193.315 36.500 193.605 ;
        RECT 36.680 193.055 37.010 193.435 ;
        RECT 37.350 193.055 37.655 194.195 ;
        RECT 37.825 193.365 38.080 194.245 ;
        RECT 38.260 194.865 38.515 195.435 ;
        RECT 38.685 195.205 39.015 195.605 ;
        RECT 39.440 195.070 39.970 195.435 ;
        RECT 39.440 195.035 39.615 195.070 ;
        RECT 38.685 194.865 39.615 195.035 ;
        RECT 38.260 194.195 38.430 194.865 ;
        RECT 38.685 194.695 38.855 194.865 ;
        RECT 38.600 194.365 38.855 194.695 ;
        RECT 39.080 194.365 39.275 194.695 ;
        RECT 38.260 193.225 38.595 194.195 ;
        RECT 38.765 193.055 38.935 194.195 ;
        RECT 39.105 193.395 39.275 194.365 ;
        RECT 39.445 193.735 39.615 194.865 ;
        RECT 39.785 194.075 39.955 194.875 ;
        RECT 40.160 194.585 40.435 195.435 ;
        RECT 40.155 194.415 40.435 194.585 ;
        RECT 40.160 194.275 40.435 194.415 ;
        RECT 40.605 194.075 40.795 195.435 ;
        RECT 40.975 195.070 41.485 195.605 ;
        RECT 41.705 194.795 41.950 195.400 ;
        RECT 42.510 194.975 42.795 195.435 ;
        RECT 42.965 195.145 43.235 195.605 ;
        RECT 42.510 194.805 43.465 194.975 ;
        RECT 40.995 194.625 42.225 194.795 ;
        RECT 39.785 193.905 40.795 194.075 ;
        RECT 40.965 194.060 41.715 194.250 ;
        RECT 39.445 193.565 40.570 193.735 ;
        RECT 40.965 193.395 41.135 194.060 ;
        RECT 41.885 193.815 42.225 194.625 ;
        RECT 42.395 194.075 43.085 194.635 ;
        RECT 43.255 193.905 43.465 194.805 ;
        RECT 39.105 193.225 41.135 193.395 ;
        RECT 41.305 193.055 41.475 193.815 ;
        RECT 41.710 193.405 42.225 193.815 ;
        RECT 42.510 193.685 43.465 193.905 ;
        RECT 43.635 194.635 44.035 195.435 ;
        RECT 44.225 194.975 44.505 195.435 ;
        RECT 45.025 195.145 45.350 195.605 ;
        RECT 44.225 194.805 45.350 194.975 ;
        RECT 45.520 194.865 45.905 195.435 ;
        RECT 44.900 194.695 45.350 194.805 ;
        RECT 43.635 194.075 44.730 194.635 ;
        RECT 44.900 194.365 45.455 194.695 ;
        RECT 42.510 193.225 42.795 193.685 ;
        RECT 42.965 193.055 43.235 193.515 ;
        RECT 43.635 193.225 44.035 194.075 ;
        RECT 44.900 193.905 45.350 194.365 ;
        RECT 45.625 194.195 45.905 194.865 ;
        RECT 44.225 193.685 45.350 193.905 ;
        RECT 44.225 193.225 44.505 193.685 ;
        RECT 45.025 193.055 45.350 193.515 ;
        RECT 45.520 193.225 45.905 194.195 ;
        RECT 46.535 194.785 47.220 195.425 ;
        RECT 47.390 194.785 47.560 195.605 ;
        RECT 47.730 194.955 48.060 195.420 ;
        RECT 48.230 195.135 48.400 195.605 ;
        RECT 48.660 195.215 49.845 195.385 ;
        RECT 50.015 195.045 50.345 195.435 ;
        RECT 49.045 194.955 49.430 195.045 ;
        RECT 47.730 194.785 49.430 194.955 ;
        RECT 49.835 194.865 50.345 195.045 ;
        RECT 50.695 195.105 50.950 195.435 ;
        RECT 51.165 195.125 51.495 195.605 ;
        RECT 51.665 195.185 53.200 195.435 ;
        RECT 50.695 195.095 50.905 195.105 ;
        RECT 50.695 195.025 50.880 195.095 ;
        RECT 46.535 193.815 46.785 194.785 ;
        RECT 46.955 194.405 47.290 194.615 ;
        RECT 47.460 194.405 47.910 194.615 ;
        RECT 48.100 194.405 48.585 194.615 ;
        RECT 47.120 194.235 47.290 194.405 ;
        RECT 48.210 194.245 48.585 194.405 ;
        RECT 48.775 194.365 49.155 194.615 ;
        RECT 49.335 194.405 49.665 194.615 ;
        RECT 47.120 194.065 48.040 194.235 ;
        RECT 46.535 193.225 47.200 193.815 ;
        RECT 47.370 193.055 47.700 193.895 ;
        RECT 47.870 193.815 48.040 194.065 ;
        RECT 48.210 194.075 48.605 194.245 ;
        RECT 48.210 193.985 48.585 194.075 ;
        RECT 48.775 193.985 49.095 194.365 ;
        RECT 49.835 194.235 50.005 194.865 ;
        RECT 50.175 194.405 50.505 194.695 ;
        RECT 49.265 194.065 50.350 194.235 ;
        RECT 49.265 193.815 49.435 194.065 ;
        RECT 47.870 193.645 49.435 193.815 ;
        RECT 48.210 193.225 49.015 193.645 ;
        RECT 49.605 193.055 49.855 193.895 ;
        RECT 50.050 193.225 50.350 194.065 ;
        RECT 50.695 193.895 50.865 195.025 ;
        RECT 51.665 194.955 51.835 195.185 ;
        RECT 51.035 194.785 51.835 194.955 ;
        RECT 51.035 194.235 51.205 194.785 ;
        RECT 52.015 194.615 52.300 195.015 ;
        RECT 51.435 194.415 51.800 194.615 ;
        RECT 51.970 194.415 52.300 194.615 ;
        RECT 52.570 194.615 52.850 195.015 ;
        RECT 53.030 194.955 53.200 195.185 ;
        RECT 53.425 195.125 53.755 195.605 ;
        RECT 53.925 194.955 54.095 195.435 ;
        RECT 53.030 194.785 54.095 194.955 ;
        RECT 54.355 194.880 54.645 195.605 ;
        RECT 54.815 194.865 55.200 195.435 ;
        RECT 55.370 195.145 55.695 195.605 ;
        RECT 56.215 194.975 56.495 195.435 ;
        RECT 52.570 194.415 53.045 194.615 ;
        RECT 53.215 194.415 53.660 194.615 ;
        RECT 53.830 194.405 54.180 194.615 ;
        RECT 51.035 194.065 54.095 194.235 ;
        RECT 50.695 193.225 50.950 193.895 ;
        RECT 51.120 193.055 51.450 193.815 ;
        RECT 51.620 193.655 53.255 193.895 ;
        RECT 51.620 193.225 51.870 193.655 ;
        RECT 53.025 193.565 53.255 193.655 ;
        RECT 52.040 193.055 52.395 193.475 ;
        RECT 52.585 193.395 52.915 193.435 ;
        RECT 53.425 193.395 53.755 193.895 ;
        RECT 52.585 193.225 53.755 193.395 ;
        RECT 53.925 193.225 54.095 194.065 ;
        RECT 54.355 193.055 54.645 194.220 ;
        RECT 54.815 194.195 55.095 194.865 ;
        RECT 55.370 194.805 56.495 194.975 ;
        RECT 55.370 194.695 55.820 194.805 ;
        RECT 55.265 194.365 55.820 194.695 ;
        RECT 56.685 194.635 57.085 195.435 ;
        RECT 57.485 195.145 57.755 195.605 ;
        RECT 57.925 194.975 58.210 195.435 ;
        RECT 54.815 193.225 55.200 194.195 ;
        RECT 55.370 193.905 55.820 194.365 ;
        RECT 55.990 194.075 57.085 194.635 ;
        RECT 55.370 193.685 56.495 193.905 ;
        RECT 55.370 193.055 55.695 193.515 ;
        RECT 56.215 193.225 56.495 193.685 ;
        RECT 56.685 193.225 57.085 194.075 ;
        RECT 57.255 194.805 58.210 194.975 ;
        RECT 58.545 195.065 58.770 195.425 ;
        RECT 58.950 195.235 59.280 195.605 ;
        RECT 59.460 195.065 59.715 195.425 ;
        RECT 60.280 195.235 61.025 195.605 ;
        RECT 58.545 194.875 61.030 195.065 ;
        RECT 57.255 193.905 57.465 194.805 ;
        RECT 57.635 194.075 58.325 194.635 ;
        RECT 58.505 194.365 58.775 194.695 ;
        RECT 58.955 194.365 59.390 194.695 ;
        RECT 59.570 194.365 60.145 194.695 ;
        RECT 60.325 194.365 60.605 194.695 ;
        RECT 60.805 194.185 61.030 194.875 ;
        RECT 58.535 194.005 61.030 194.185 ;
        RECT 61.205 194.005 61.540 195.425 ;
        RECT 61.715 194.805 62.025 195.605 ;
        RECT 62.230 194.805 62.925 195.435 ;
        RECT 63.565 194.880 63.895 195.390 ;
        RECT 64.065 195.205 64.395 195.605 ;
        RECT 65.445 195.035 65.775 195.375 ;
        RECT 65.945 195.205 66.275 195.605 ;
        RECT 61.725 194.365 62.060 194.635 ;
        RECT 62.230 194.205 62.400 194.805 ;
        RECT 62.570 194.365 62.905 194.615 ;
        RECT 63.565 194.245 63.755 194.880 ;
        RECT 64.065 194.865 66.430 195.035 ;
        RECT 64.065 194.695 64.235 194.865 ;
        RECT 63.925 194.365 64.235 194.695 ;
        RECT 64.405 194.365 64.710 194.695 ;
        RECT 57.255 193.685 58.210 193.905 ;
        RECT 57.485 193.055 57.755 193.515 ;
        RECT 57.925 193.225 58.210 193.685 ;
        RECT 58.535 193.235 58.825 194.005 ;
        RECT 59.395 193.595 60.585 193.825 ;
        RECT 59.395 193.235 59.655 193.595 ;
        RECT 59.825 193.055 60.155 193.425 ;
        RECT 60.325 193.235 60.585 193.595 ;
        RECT 60.775 193.055 61.105 193.775 ;
        RECT 61.275 193.235 61.540 194.005 ;
        RECT 61.715 193.055 61.995 194.195 ;
        RECT 62.165 193.225 62.495 194.205 ;
        RECT 62.665 193.055 62.925 194.195 ;
        RECT 63.565 194.115 63.785 194.245 ;
        RECT 63.565 193.265 63.895 194.115 ;
        RECT 64.065 193.055 64.315 194.195 ;
        RECT 64.495 194.035 64.710 194.365 ;
        RECT 64.885 194.035 65.170 194.695 ;
        RECT 65.365 194.035 65.630 194.695 ;
        RECT 65.845 194.035 66.090 194.695 ;
        RECT 66.260 193.865 66.430 194.865 ;
        RECT 66.775 194.835 70.285 195.605 ;
        RECT 66.775 194.315 68.425 194.835 ;
        RECT 70.465 194.795 70.735 195.605 ;
        RECT 70.905 194.795 71.235 195.435 ;
        RECT 71.405 194.795 71.645 195.605 ;
        RECT 71.835 194.865 72.275 195.425 ;
        RECT 72.445 194.865 72.895 195.605 ;
        RECT 73.065 195.035 73.235 195.435 ;
        RECT 73.405 195.205 73.825 195.605 ;
        RECT 73.995 195.035 74.225 195.435 ;
        RECT 73.065 194.865 74.225 195.035 ;
        RECT 74.395 194.865 74.885 195.435 ;
        RECT 68.595 194.145 70.285 194.665 ;
        RECT 70.455 194.365 70.805 194.615 ;
        RECT 70.975 194.195 71.145 194.795 ;
        RECT 71.315 194.365 71.665 194.615 ;
        RECT 64.505 193.695 65.795 193.865 ;
        RECT 64.505 193.275 64.755 193.695 ;
        RECT 64.985 193.055 65.315 193.525 ;
        RECT 65.545 193.275 65.795 193.695 ;
        RECT 65.975 193.695 66.430 193.865 ;
        RECT 65.975 193.265 66.305 193.695 ;
        RECT 66.775 193.055 70.285 194.145 ;
        RECT 70.465 193.055 70.795 194.195 ;
        RECT 70.975 194.025 71.655 194.195 ;
        RECT 71.325 193.240 71.655 194.025 ;
        RECT 71.835 193.855 72.145 194.865 ;
        RECT 72.315 194.245 72.485 194.695 ;
        RECT 72.655 194.415 73.045 194.695 ;
        RECT 73.230 194.365 73.475 194.695 ;
        RECT 72.315 194.075 73.105 194.245 ;
        RECT 71.835 193.225 72.275 193.855 ;
        RECT 72.450 193.055 72.765 193.905 ;
        RECT 72.935 193.395 73.105 194.075 ;
        RECT 73.275 193.565 73.475 194.365 ;
        RECT 73.675 193.565 73.925 194.695 ;
        RECT 74.140 194.365 74.545 194.695 ;
        RECT 74.715 194.195 74.885 194.865 ;
        RECT 75.055 194.835 78.565 195.605 ;
        RECT 78.735 194.855 79.945 195.605 ;
        RECT 80.115 194.880 80.405 195.605 ;
        RECT 75.055 194.315 76.705 194.835 ;
        RECT 74.115 194.025 74.885 194.195 ;
        RECT 76.875 194.145 78.565 194.665 ;
        RECT 78.735 194.315 79.255 194.855 ;
        RECT 80.590 194.825 80.885 195.605 ;
        RECT 81.445 195.075 81.790 195.435 ;
        RECT 82.250 195.245 82.580 195.605 ;
        RECT 82.785 195.075 83.105 195.435 ;
        RECT 81.445 194.905 83.105 195.075 ;
        RECT 79.425 194.145 79.945 194.685 ;
        RECT 74.115 193.395 74.365 194.025 ;
        RECT 72.935 193.225 74.365 193.395 ;
        RECT 74.545 193.055 74.875 193.855 ;
        RECT 75.055 193.055 78.565 194.145 ;
        RECT 78.735 193.055 79.945 194.145 ;
        RECT 80.115 193.055 80.405 194.220 ;
        RECT 80.635 194.195 81.135 194.655 ;
        RECT 81.305 194.365 81.915 194.695 ;
        RECT 82.095 194.445 82.425 194.615 ;
        RECT 82.095 194.195 82.420 194.445 ;
        RECT 80.635 194.015 82.420 194.195 ;
        RECT 80.600 193.665 82.635 193.835 ;
        RECT 80.600 193.585 81.710 193.665 ;
        RECT 80.600 193.225 80.860 193.585 ;
        RECT 81.030 193.055 81.360 193.415 ;
        RECT 81.540 193.225 81.710 193.585 ;
        RECT 81.965 193.055 82.135 193.495 ;
        RECT 82.305 193.405 82.635 193.665 ;
        RECT 82.805 193.575 83.105 194.905 ;
        RECT 83.285 194.865 83.615 195.605 ;
        RECT 83.795 194.805 84.490 195.435 ;
        RECT 84.695 194.805 85.005 195.605 ;
        RECT 83.290 194.065 83.565 194.695 ;
        RECT 83.815 194.365 84.150 194.615 ;
        RECT 84.320 194.205 84.490 194.805 ;
        RECT 86.105 194.795 86.375 195.605 ;
        RECT 86.545 194.795 86.875 195.435 ;
        RECT 87.045 194.795 87.285 195.605 ;
        RECT 87.475 195.060 92.820 195.605 ;
        RECT 84.660 194.365 84.995 194.635 ;
        RECT 86.095 194.365 86.445 194.615 ;
        RECT 83.275 193.405 83.580 193.895 ;
        RECT 82.305 193.225 83.580 193.405 ;
        RECT 83.795 193.055 84.055 194.195 ;
        RECT 84.225 193.225 84.555 194.205 ;
        RECT 86.615 194.195 86.785 194.795 ;
        RECT 86.955 194.365 87.305 194.615 ;
        RECT 89.060 194.230 89.400 195.060 ;
        RECT 92.995 194.835 96.505 195.605 ;
        RECT 84.725 193.055 85.005 194.195 ;
        RECT 86.105 193.055 86.435 194.195 ;
        RECT 86.615 194.025 87.295 194.195 ;
        RECT 86.965 193.240 87.295 194.025 ;
        RECT 90.880 193.490 91.230 194.740 ;
        RECT 92.995 194.315 94.645 194.835 ;
        RECT 94.815 194.145 96.505 194.665 ;
        RECT 87.475 193.055 92.820 193.490 ;
        RECT 92.995 193.055 96.505 194.145 ;
        RECT 96.685 193.235 96.945 195.425 ;
        RECT 97.205 195.235 97.875 195.605 ;
        RECT 98.055 195.055 98.365 195.425 ;
        RECT 97.135 194.855 98.365 195.055 ;
        RECT 97.135 194.185 97.425 194.855 ;
        RECT 98.545 194.675 98.775 195.315 ;
        RECT 98.955 194.875 99.245 195.605 ;
        RECT 99.435 194.805 100.130 195.435 ;
        RECT 100.335 194.805 100.645 195.605 ;
        RECT 100.815 194.805 101.510 195.435 ;
        RECT 101.715 194.805 102.025 195.605 ;
        RECT 102.195 194.835 105.705 195.605 ;
        RECT 105.875 194.880 106.165 195.605 ;
        RECT 106.335 194.835 109.845 195.605 ;
        RECT 97.605 194.365 98.070 194.675 ;
        RECT 98.250 194.365 98.775 194.675 ;
        RECT 98.955 194.365 99.255 194.695 ;
        RECT 99.455 194.365 99.790 194.615 ;
        RECT 99.960 194.245 100.130 194.805 ;
        RECT 100.300 194.365 100.635 194.635 ;
        RECT 100.835 194.365 101.170 194.615 ;
        RECT 99.955 194.205 100.130 194.245 ;
        RECT 101.340 194.205 101.510 194.805 ;
        RECT 101.680 194.365 102.015 194.635 ;
        RECT 102.195 194.315 103.845 194.835 ;
        RECT 97.135 193.965 97.905 194.185 ;
        RECT 97.115 193.055 97.455 193.785 ;
        RECT 97.635 193.235 97.905 193.965 ;
        RECT 98.085 193.945 99.245 194.185 ;
        RECT 98.085 193.235 98.315 193.945 ;
        RECT 98.485 193.055 98.815 193.765 ;
        RECT 98.985 193.235 99.245 193.945 ;
        RECT 99.435 193.055 99.695 194.195 ;
        RECT 99.865 193.225 100.195 194.205 ;
        RECT 100.365 193.055 100.645 194.195 ;
        RECT 100.815 193.055 101.075 194.195 ;
        RECT 101.245 193.225 101.575 194.205 ;
        RECT 101.745 193.055 102.025 194.195 ;
        RECT 104.015 194.145 105.705 194.665 ;
        RECT 106.335 194.315 107.985 194.835 ;
        RECT 110.015 194.785 110.275 195.605 ;
        RECT 110.445 194.785 110.775 195.205 ;
        RECT 110.955 195.120 111.745 195.385 ;
        RECT 110.525 194.695 110.775 194.785 ;
        RECT 102.195 193.055 105.705 194.145 ;
        RECT 105.875 193.055 106.165 194.220 ;
        RECT 108.155 194.145 109.845 194.665 ;
        RECT 106.335 193.055 109.845 194.145 ;
        RECT 110.015 193.735 110.355 194.615 ;
        RECT 110.525 194.445 111.320 194.695 ;
        RECT 110.015 193.055 110.275 193.565 ;
        RECT 110.525 193.225 110.695 194.445 ;
        RECT 111.490 194.265 111.745 195.120 ;
        RECT 111.915 194.965 112.115 195.385 ;
        RECT 112.305 195.145 112.635 195.605 ;
        RECT 111.915 194.445 112.325 194.965 ;
        RECT 112.805 194.955 113.065 195.435 ;
        RECT 112.495 194.265 112.725 194.695 ;
        RECT 110.935 194.095 112.725 194.265 ;
        RECT 110.935 193.730 111.185 194.095 ;
        RECT 111.355 193.735 111.685 193.925 ;
        RECT 111.905 193.800 112.620 194.095 ;
        RECT 112.895 193.925 113.065 194.955 ;
        RECT 111.355 193.560 111.550 193.735 ;
        RECT 110.935 193.055 111.550 193.560 ;
        RECT 111.720 193.225 112.195 193.565 ;
        RECT 112.365 193.055 112.580 193.600 ;
        RECT 112.790 193.225 113.065 193.925 ;
        RECT 114.155 195.020 114.465 195.435 ;
        RECT 114.660 195.225 114.990 195.605 ;
        RECT 115.160 195.265 116.565 195.435 ;
        RECT 115.160 195.035 115.330 195.265 ;
        RECT 114.155 193.905 114.325 195.020 ;
        RECT 114.635 194.865 115.330 195.035 ;
        RECT 116.395 195.035 116.565 195.265 ;
        RECT 116.835 195.205 117.165 195.605 ;
        RECT 117.405 195.035 117.575 195.435 ;
        RECT 114.635 194.695 114.805 194.865 ;
        RECT 114.495 194.365 114.805 194.695 ;
        RECT 114.975 194.365 115.310 194.695 ;
        RECT 115.580 194.365 115.775 194.940 ;
        RECT 116.035 194.695 116.225 194.925 ;
        RECT 116.395 194.865 117.575 195.035 ;
        RECT 117.835 194.835 121.345 195.605 ;
        RECT 116.035 194.365 116.380 194.695 ;
        RECT 116.690 194.365 117.165 194.695 ;
        RECT 117.420 194.365 117.605 194.695 ;
        RECT 114.635 194.195 114.805 194.365 ;
        RECT 117.835 194.315 119.485 194.835 ;
        RECT 121.515 194.805 121.825 195.605 ;
        RECT 122.030 194.805 122.725 195.435 ;
        RECT 122.955 195.125 123.235 195.605 ;
        RECT 123.405 194.955 123.665 195.345 ;
        RECT 123.840 195.125 124.095 195.605 ;
        RECT 124.265 194.955 124.560 195.345 ;
        RECT 124.740 195.125 125.015 195.605 ;
        RECT 125.185 195.105 125.485 195.435 ;
        RECT 125.675 195.120 126.465 195.385 ;
        RECT 122.030 194.755 122.205 194.805 ;
        RECT 122.910 194.785 124.560 194.955 ;
        RECT 114.635 194.025 117.575 194.195 ;
        RECT 119.655 194.145 121.345 194.665 ;
        RECT 121.525 194.365 121.860 194.635 ;
        RECT 122.030 194.205 122.200 194.755 ;
        RECT 122.370 194.365 122.705 194.615 ;
        RECT 122.910 194.275 123.315 194.785 ;
        RECT 123.485 194.445 124.625 194.615 ;
        RECT 114.155 193.265 114.495 193.905 ;
        RECT 115.085 193.685 116.645 193.855 ;
        RECT 114.665 193.055 114.910 193.515 ;
        RECT 115.085 193.225 115.335 193.685 ;
        RECT 115.525 193.055 116.195 193.435 ;
        RECT 116.395 193.225 116.645 193.685 ;
        RECT 117.405 193.225 117.575 194.025 ;
        RECT 117.835 193.055 121.345 194.145 ;
        RECT 121.515 193.055 121.795 194.195 ;
        RECT 121.965 193.225 122.295 194.205 ;
        RECT 122.465 193.055 122.725 194.195 ;
        RECT 122.910 194.105 123.665 194.275 ;
        RECT 122.950 193.055 123.235 193.925 ;
        RECT 123.405 193.855 123.665 194.105 ;
        RECT 124.455 194.195 124.625 194.445 ;
        RECT 124.795 194.365 125.145 194.935 ;
        RECT 125.315 194.195 125.485 195.105 ;
        RECT 125.655 194.445 126.040 194.925 ;
        RECT 126.210 194.265 126.465 195.120 ;
        RECT 126.635 194.940 126.865 195.385 ;
        RECT 127.045 195.110 127.375 195.605 ;
        RECT 127.550 194.975 127.800 195.435 ;
        RECT 126.635 194.445 127.045 194.940 ;
        RECT 127.630 194.765 127.800 194.975 ;
        RECT 127.970 194.945 128.245 195.605 ;
        RECT 128.505 194.925 128.675 195.300 ;
        RECT 127.230 194.265 127.460 194.695 ;
        RECT 124.455 194.025 125.485 194.195 ;
        RECT 123.405 193.685 124.525 193.855 ;
        RECT 123.405 193.225 123.665 193.685 ;
        RECT 123.840 193.055 124.095 193.515 ;
        RECT 124.265 193.225 124.525 193.685 ;
        RECT 124.695 193.055 125.005 193.855 ;
        RECT 125.175 193.225 125.485 194.025 ;
        RECT 125.670 194.095 127.460 194.265 ;
        RECT 127.630 194.245 128.245 194.765 ;
        RECT 128.475 194.755 128.675 194.925 ;
        RECT 128.865 195.075 129.095 195.380 ;
        RECT 129.265 195.245 129.595 195.605 ;
        RECT 129.790 195.075 130.080 195.425 ;
        RECT 128.865 194.905 130.080 195.075 ;
        RECT 128.505 194.735 128.675 194.755 ;
        RECT 130.255 194.855 131.465 195.605 ;
        RECT 131.635 194.880 131.925 195.605 ;
        RECT 128.505 194.565 129.025 194.735 ;
        RECT 125.670 193.730 125.925 194.095 ;
        RECT 126.095 193.735 126.425 193.925 ;
        RECT 126.650 193.800 126.900 194.095 ;
        RECT 127.645 193.905 127.815 194.245 ;
        RECT 126.095 193.560 126.285 193.735 ;
        RECT 125.655 193.055 126.285 193.560 ;
        RECT 126.465 193.225 126.940 193.565 ;
        RECT 127.125 193.055 127.340 193.900 ;
        RECT 127.555 193.895 127.815 193.905 ;
        RECT 127.540 193.225 127.815 193.895 ;
        RECT 127.985 193.055 128.245 194.065 ;
        RECT 128.420 194.035 128.665 194.395 ;
        RECT 128.855 194.185 129.025 194.565 ;
        RECT 129.195 194.365 129.580 194.695 ;
        RECT 129.760 194.585 130.020 194.695 ;
        RECT 129.760 194.415 130.025 194.585 ;
        RECT 129.760 194.365 130.020 194.415 ;
        RECT 128.855 193.905 129.205 194.185 ;
        RECT 128.420 193.055 128.675 193.855 ;
        RECT 128.875 193.225 129.205 193.905 ;
        RECT 129.385 193.315 129.580 194.365 ;
        RECT 130.255 194.315 130.775 194.855 ;
        RECT 132.095 194.805 132.435 195.435 ;
        RECT 132.605 194.805 132.855 195.605 ;
        RECT 133.045 194.955 133.375 195.435 ;
        RECT 133.545 195.145 133.770 195.605 ;
        RECT 133.940 194.955 134.270 195.435 ;
        RECT 129.760 193.055 130.080 194.195 ;
        RECT 130.945 194.145 131.465 194.685 ;
        RECT 130.255 193.055 131.465 194.145 ;
        RECT 131.635 193.055 131.925 194.220 ;
        RECT 132.095 194.195 132.270 194.805 ;
        RECT 133.045 194.785 134.270 194.955 ;
        RECT 134.900 194.825 135.400 195.435 ;
        RECT 132.440 194.445 133.135 194.615 ;
        RECT 132.965 194.195 133.135 194.445 ;
        RECT 133.310 194.415 133.730 194.615 ;
        RECT 133.900 194.415 134.230 194.615 ;
        RECT 134.400 194.415 134.730 194.615 ;
        RECT 134.900 194.195 135.070 194.825 ;
        RECT 135.775 194.805 136.470 195.435 ;
        RECT 136.675 194.805 136.985 195.605 ;
        RECT 137.155 194.835 139.745 195.605 ;
        RECT 140.005 195.055 140.175 195.435 ;
        RECT 140.390 195.225 140.720 195.605 ;
        RECT 140.005 194.885 140.720 195.055 ;
        RECT 135.255 194.365 135.605 194.615 ;
        RECT 135.795 194.365 136.130 194.615 ;
        RECT 136.300 194.205 136.470 194.805 ;
        RECT 136.640 194.365 136.975 194.635 ;
        RECT 137.155 194.315 138.365 194.835 ;
        RECT 132.095 193.225 132.435 194.195 ;
        RECT 132.605 193.055 132.775 194.195 ;
        RECT 132.965 194.025 135.400 194.195 ;
        RECT 133.045 193.055 133.295 193.855 ;
        RECT 133.940 193.225 134.270 194.025 ;
        RECT 134.570 193.055 134.900 193.855 ;
        RECT 135.070 193.225 135.400 194.025 ;
        RECT 135.775 193.055 136.035 194.195 ;
        RECT 136.205 193.225 136.535 194.205 ;
        RECT 136.705 193.055 136.985 194.195 ;
        RECT 138.535 194.145 139.745 194.665 ;
        RECT 139.915 194.335 140.270 194.705 ;
        RECT 140.550 194.695 140.720 194.885 ;
        RECT 140.890 194.860 141.145 195.435 ;
        RECT 140.550 194.365 140.805 194.695 ;
        RECT 140.550 194.155 140.720 194.365 ;
        RECT 137.155 193.055 139.745 194.145 ;
        RECT 140.005 193.985 140.720 194.155 ;
        RECT 140.975 194.130 141.145 194.860 ;
        RECT 141.320 194.765 141.580 195.605 ;
        RECT 141.755 194.855 142.965 195.605 ;
        RECT 141.755 194.315 142.275 194.855 ;
        RECT 143.145 194.795 143.415 195.605 ;
        RECT 143.585 194.795 143.915 195.435 ;
        RECT 144.085 194.795 144.325 195.605 ;
        RECT 140.005 193.225 140.175 193.985 ;
        RECT 140.390 193.055 140.720 193.815 ;
        RECT 140.890 193.225 141.145 194.130 ;
        RECT 141.320 193.055 141.580 194.205 ;
        RECT 142.445 194.145 142.965 194.685 ;
        RECT 143.135 194.365 143.485 194.615 ;
        RECT 143.655 194.195 143.825 194.795 ;
        RECT 144.515 194.620 144.785 195.435 ;
        RECT 144.955 194.865 145.625 195.605 ;
        RECT 145.795 195.035 146.090 195.380 ;
        RECT 146.270 195.205 146.645 195.605 ;
        RECT 146.860 195.035 147.190 195.380 ;
        RECT 145.795 194.865 147.190 195.035 ;
        RECT 147.440 194.865 148.025 195.435 ;
        RECT 148.195 195.060 153.540 195.605 ;
        RECT 143.995 194.365 144.345 194.615 ;
        RECT 141.755 193.055 142.965 194.145 ;
        RECT 143.145 193.055 143.475 194.195 ;
        RECT 143.655 194.025 144.335 194.195 ;
        RECT 144.005 193.240 144.335 194.025 ;
        RECT 144.515 193.225 144.865 194.620 ;
        RECT 145.035 194.195 145.205 194.695 ;
        RECT 145.375 194.365 145.710 194.695 ;
        RECT 145.880 194.365 146.220 194.695 ;
        RECT 145.035 194.025 145.780 194.195 ;
        RECT 145.035 193.055 145.440 193.855 ;
        RECT 145.610 193.395 145.780 194.025 ;
        RECT 145.950 193.620 146.220 194.365 ;
        RECT 146.410 194.365 146.700 194.695 ;
        RECT 146.870 194.365 147.270 194.695 ;
        RECT 146.410 193.620 146.645 194.365 ;
        RECT 147.440 194.195 147.610 194.865 ;
        RECT 147.780 194.365 148.025 194.695 ;
        RECT 149.780 194.230 150.120 195.060 ;
        RECT 153.715 194.835 156.305 195.605 ;
        RECT 156.935 194.855 158.145 195.605 ;
        RECT 146.815 194.025 148.025 194.195 ;
        RECT 146.815 193.395 147.145 194.025 ;
        RECT 145.610 193.225 147.145 193.395 ;
        RECT 147.330 193.055 147.565 193.855 ;
        RECT 147.735 193.225 148.025 194.025 ;
        RECT 151.600 193.490 151.950 194.740 ;
        RECT 153.715 194.315 154.925 194.835 ;
        RECT 155.095 194.145 156.305 194.665 ;
        RECT 148.195 193.055 153.540 193.490 ;
        RECT 153.715 193.055 156.305 194.145 ;
        RECT 156.935 194.145 157.455 194.685 ;
        RECT 157.625 194.315 158.145 194.855 ;
        RECT 156.935 193.055 158.145 194.145 ;
        RECT 2.750 192.885 158.230 193.055 ;
        RECT 2.835 191.795 4.045 192.885 ;
        RECT 4.215 191.795 5.885 192.885 ;
        RECT 2.835 191.085 3.355 191.625 ;
        RECT 3.525 191.255 4.045 191.795 ;
        RECT 4.215 191.105 4.965 191.625 ;
        RECT 5.135 191.275 5.885 191.795 ;
        RECT 6.055 191.810 6.325 192.715 ;
        RECT 6.495 192.125 6.825 192.885 ;
        RECT 7.005 191.955 7.175 192.715 ;
        RECT 2.835 190.335 4.045 191.085 ;
        RECT 4.215 190.335 5.885 191.105 ;
        RECT 6.055 191.010 6.225 191.810 ;
        RECT 6.510 191.785 7.175 191.955 ;
        RECT 6.510 191.640 6.680 191.785 ;
        RECT 6.395 191.310 6.680 191.640 ;
        RECT 7.440 191.745 7.775 192.715 ;
        RECT 7.945 191.745 8.115 192.885 ;
        RECT 8.285 192.545 10.315 192.715 ;
        RECT 6.510 191.055 6.680 191.310 ;
        RECT 6.915 191.235 7.245 191.605 ;
        RECT 7.440 191.075 7.610 191.745 ;
        RECT 8.285 191.575 8.455 192.545 ;
        RECT 7.780 191.245 8.035 191.575 ;
        RECT 8.260 191.245 8.455 191.575 ;
        RECT 8.625 192.205 9.750 192.375 ;
        RECT 7.865 191.075 8.035 191.245 ;
        RECT 8.625 191.075 8.795 192.205 ;
        RECT 6.055 190.505 6.315 191.010 ;
        RECT 6.510 190.885 7.175 191.055 ;
        RECT 6.495 190.335 6.825 190.715 ;
        RECT 7.005 190.505 7.175 190.885 ;
        RECT 7.440 190.505 7.695 191.075 ;
        RECT 7.865 190.905 8.795 191.075 ;
        RECT 8.965 191.865 9.975 192.035 ;
        RECT 8.965 191.065 9.135 191.865 ;
        RECT 9.340 191.525 9.615 191.665 ;
        RECT 9.335 191.355 9.615 191.525 ;
        RECT 8.620 190.870 8.795 190.905 ;
        RECT 7.865 190.335 8.195 190.735 ;
        RECT 8.620 190.505 9.150 190.870 ;
        RECT 9.340 190.505 9.615 191.355 ;
        RECT 9.785 190.505 9.975 191.865 ;
        RECT 10.145 191.880 10.315 192.545 ;
        RECT 10.485 192.125 10.655 192.885 ;
        RECT 10.890 192.125 11.405 192.535 ;
        RECT 10.145 191.690 10.895 191.880 ;
        RECT 11.065 191.315 11.405 192.125 ;
        RECT 10.175 191.145 11.405 191.315 ;
        RECT 11.580 191.745 11.915 192.715 ;
        RECT 12.085 191.745 12.255 192.885 ;
        RECT 12.425 192.545 14.455 192.715 ;
        RECT 10.155 190.335 10.665 190.870 ;
        RECT 10.885 190.540 11.130 191.145 ;
        RECT 11.580 191.075 11.750 191.745 ;
        RECT 12.425 191.575 12.595 192.545 ;
        RECT 11.920 191.245 12.175 191.575 ;
        RECT 12.400 191.245 12.595 191.575 ;
        RECT 12.765 192.205 13.890 192.375 ;
        RECT 12.005 191.075 12.175 191.245 ;
        RECT 12.765 191.075 12.935 192.205 ;
        RECT 11.580 190.505 11.835 191.075 ;
        RECT 12.005 190.905 12.935 191.075 ;
        RECT 13.105 191.865 14.115 192.035 ;
        RECT 13.105 191.065 13.275 191.865 ;
        RECT 13.480 191.525 13.755 191.665 ;
        RECT 13.475 191.355 13.755 191.525 ;
        RECT 12.760 190.870 12.935 190.905 ;
        RECT 12.005 190.335 12.335 190.735 ;
        RECT 12.760 190.505 13.290 190.870 ;
        RECT 13.480 190.505 13.755 191.355 ;
        RECT 13.925 190.505 14.115 191.865 ;
        RECT 14.285 191.880 14.455 192.545 ;
        RECT 14.625 192.125 14.795 192.885 ;
        RECT 15.030 192.125 15.545 192.535 ;
        RECT 14.285 191.690 15.035 191.880 ;
        RECT 15.205 191.315 15.545 192.125 ;
        RECT 15.715 191.720 16.005 192.885 ;
        RECT 16.640 191.745 16.975 192.715 ;
        RECT 17.145 191.745 17.315 192.885 ;
        RECT 17.485 192.545 19.515 192.715 ;
        RECT 14.315 191.145 15.545 191.315 ;
        RECT 14.295 190.335 14.805 190.870 ;
        RECT 15.025 190.540 15.270 191.145 ;
        RECT 16.640 191.075 16.810 191.745 ;
        RECT 17.485 191.575 17.655 192.545 ;
        RECT 16.980 191.245 17.235 191.575 ;
        RECT 17.460 191.245 17.655 191.575 ;
        RECT 17.825 192.205 18.950 192.375 ;
        RECT 17.065 191.075 17.235 191.245 ;
        RECT 17.825 191.075 17.995 192.205 ;
        RECT 15.715 190.335 16.005 191.060 ;
        RECT 16.640 190.505 16.895 191.075 ;
        RECT 17.065 190.905 17.995 191.075 ;
        RECT 18.165 191.865 19.175 192.035 ;
        RECT 18.165 191.065 18.335 191.865 ;
        RECT 18.540 191.525 18.815 191.665 ;
        RECT 18.535 191.355 18.815 191.525 ;
        RECT 17.820 190.870 17.995 190.905 ;
        RECT 17.065 190.335 17.395 190.735 ;
        RECT 17.820 190.505 18.350 190.870 ;
        RECT 18.540 190.505 18.815 191.355 ;
        RECT 18.985 190.505 19.175 191.865 ;
        RECT 19.345 191.880 19.515 192.545 ;
        RECT 19.685 192.125 19.855 192.885 ;
        RECT 20.090 192.125 20.605 192.535 ;
        RECT 19.345 191.690 20.095 191.880 ;
        RECT 20.265 191.315 20.605 192.125 ;
        RECT 19.375 191.145 20.605 191.315 ;
        RECT 20.775 192.125 21.290 192.535 ;
        RECT 21.525 192.125 21.695 192.885 ;
        RECT 21.865 192.545 23.895 192.715 ;
        RECT 20.775 191.315 21.115 192.125 ;
        RECT 21.865 191.880 22.035 192.545 ;
        RECT 22.430 192.205 23.555 192.375 ;
        RECT 21.285 191.690 22.035 191.880 ;
        RECT 22.205 191.865 23.215 192.035 ;
        RECT 20.775 191.145 22.005 191.315 ;
        RECT 19.355 190.335 19.865 190.870 ;
        RECT 20.085 190.540 20.330 191.145 ;
        RECT 21.050 190.540 21.295 191.145 ;
        RECT 21.515 190.335 22.025 190.870 ;
        RECT 22.205 190.505 22.395 191.865 ;
        RECT 22.565 190.845 22.840 191.665 ;
        RECT 23.045 191.065 23.215 191.865 ;
        RECT 23.385 191.075 23.555 192.205 ;
        RECT 23.725 191.575 23.895 192.545 ;
        RECT 24.065 191.745 24.235 192.885 ;
        RECT 24.405 191.745 24.740 192.715 ;
        RECT 23.725 191.245 23.920 191.575 ;
        RECT 24.145 191.245 24.400 191.575 ;
        RECT 24.145 191.075 24.315 191.245 ;
        RECT 24.570 191.075 24.740 191.745 ;
        RECT 24.915 192.125 25.430 192.535 ;
        RECT 25.665 192.125 25.835 192.885 ;
        RECT 26.005 192.545 28.035 192.715 ;
        RECT 24.915 191.315 25.255 192.125 ;
        RECT 26.005 191.880 26.175 192.545 ;
        RECT 26.570 192.205 27.695 192.375 ;
        RECT 25.425 191.690 26.175 191.880 ;
        RECT 26.345 191.865 27.355 192.035 ;
        RECT 24.915 191.145 26.145 191.315 ;
        RECT 23.385 190.905 24.315 191.075 ;
        RECT 23.385 190.870 23.560 190.905 ;
        RECT 22.565 190.675 22.845 190.845 ;
        RECT 22.565 190.505 22.840 190.675 ;
        RECT 23.030 190.505 23.560 190.870 ;
        RECT 23.985 190.335 24.315 190.735 ;
        RECT 24.485 190.505 24.740 191.075 ;
        RECT 25.190 190.540 25.435 191.145 ;
        RECT 25.655 190.335 26.165 190.870 ;
        RECT 26.345 190.505 26.535 191.865 ;
        RECT 26.705 191.525 26.980 191.665 ;
        RECT 26.705 191.355 26.985 191.525 ;
        RECT 26.705 190.505 26.980 191.355 ;
        RECT 27.185 191.065 27.355 191.865 ;
        RECT 27.525 191.075 27.695 192.205 ;
        RECT 27.865 191.575 28.035 192.545 ;
        RECT 28.205 191.745 28.375 192.885 ;
        RECT 28.545 191.745 28.880 192.715 ;
        RECT 29.060 192.215 29.315 192.715 ;
        RECT 29.485 192.385 29.815 192.885 ;
        RECT 29.060 192.045 29.810 192.215 ;
        RECT 27.865 191.245 28.060 191.575 ;
        RECT 28.285 191.245 28.540 191.575 ;
        RECT 28.285 191.075 28.455 191.245 ;
        RECT 28.710 191.075 28.880 191.745 ;
        RECT 29.060 191.225 29.410 191.875 ;
        RECT 27.525 190.905 28.455 191.075 ;
        RECT 27.525 190.870 27.700 190.905 ;
        RECT 27.170 190.505 27.700 190.870 ;
        RECT 28.125 190.335 28.455 190.735 ;
        RECT 28.625 190.505 28.880 191.075 ;
        RECT 29.580 191.055 29.810 192.045 ;
        RECT 29.060 190.885 29.810 191.055 ;
        RECT 29.060 190.595 29.315 190.885 ;
        RECT 29.485 190.335 29.815 190.715 ;
        RECT 29.985 190.595 30.155 192.715 ;
        RECT 30.325 191.915 30.650 192.700 ;
        RECT 30.820 192.425 31.070 192.885 ;
        RECT 31.240 192.385 31.490 192.715 ;
        RECT 31.705 192.385 32.385 192.715 ;
        RECT 31.240 192.255 31.410 192.385 ;
        RECT 31.015 192.085 31.410 192.255 ;
        RECT 30.385 190.865 30.845 191.915 ;
        RECT 31.015 190.725 31.185 192.085 ;
        RECT 31.580 191.825 32.045 192.215 ;
        RECT 31.355 191.015 31.705 191.635 ;
        RECT 31.875 191.235 32.045 191.825 ;
        RECT 32.215 191.605 32.385 192.385 ;
        RECT 32.555 192.285 32.725 192.625 ;
        RECT 32.960 192.455 33.290 192.885 ;
        RECT 33.460 192.285 33.630 192.625 ;
        RECT 33.925 192.425 34.295 192.885 ;
        RECT 32.555 192.115 33.630 192.285 ;
        RECT 34.465 192.255 34.635 192.715 ;
        RECT 34.870 192.375 35.740 192.715 ;
        RECT 35.910 192.425 36.160 192.885 ;
        RECT 34.075 192.085 34.635 192.255 ;
        RECT 34.075 191.945 34.245 192.085 ;
        RECT 32.745 191.775 34.245 191.945 ;
        RECT 34.940 191.915 35.400 192.205 ;
        RECT 32.215 191.435 33.905 191.605 ;
        RECT 31.875 191.015 32.230 191.235 ;
        RECT 32.400 190.725 32.570 191.435 ;
        RECT 32.775 191.015 33.565 191.265 ;
        RECT 33.735 191.255 33.905 191.435 ;
        RECT 34.075 191.085 34.245 191.775 ;
        RECT 30.515 190.335 30.845 190.695 ;
        RECT 31.015 190.555 31.510 190.725 ;
        RECT 31.715 190.555 32.570 190.725 ;
        RECT 33.445 190.335 33.775 190.795 ;
        RECT 33.985 190.695 34.245 191.085 ;
        RECT 34.435 191.905 35.400 191.915 ;
        RECT 35.570 191.995 35.740 192.375 ;
        RECT 36.330 192.335 36.500 192.625 ;
        RECT 36.680 192.505 37.010 192.885 ;
        RECT 36.330 192.165 37.130 192.335 ;
        RECT 34.435 191.745 35.110 191.905 ;
        RECT 35.570 191.825 36.790 191.995 ;
        RECT 34.435 190.955 34.645 191.745 ;
        RECT 35.570 191.735 35.740 191.825 ;
        RECT 34.815 190.955 35.165 191.575 ;
        RECT 35.335 191.565 35.740 191.735 ;
        RECT 35.335 190.785 35.505 191.565 ;
        RECT 35.675 191.115 35.895 191.395 ;
        RECT 36.075 191.285 36.615 191.655 ;
        RECT 36.960 191.575 37.130 192.165 ;
        RECT 37.350 191.745 37.655 192.885 ;
        RECT 37.825 191.695 38.080 192.575 ;
        RECT 39.375 192.215 39.655 192.885 ;
        RECT 39.825 191.995 40.125 192.545 ;
        RECT 40.325 192.165 40.655 192.885 ;
        RECT 40.845 192.165 41.305 192.715 ;
        RECT 36.960 191.545 37.700 191.575 ;
        RECT 35.675 190.945 36.205 191.115 ;
        RECT 33.985 190.525 34.335 190.695 ;
        RECT 34.555 190.505 35.505 190.785 ;
        RECT 35.675 190.335 35.865 190.775 ;
        RECT 36.035 190.715 36.205 190.945 ;
        RECT 36.375 190.885 36.615 191.285 ;
        RECT 36.785 191.245 37.700 191.545 ;
        RECT 36.785 191.070 37.110 191.245 ;
        RECT 36.785 190.715 37.105 191.070 ;
        RECT 37.870 191.045 38.080 191.695 ;
        RECT 39.190 191.575 39.455 191.935 ;
        RECT 39.825 191.825 40.765 191.995 ;
        RECT 40.595 191.575 40.765 191.825 ;
        RECT 39.190 191.325 39.865 191.575 ;
        RECT 40.085 191.325 40.425 191.575 ;
        RECT 40.595 191.245 40.885 191.575 ;
        RECT 40.595 191.155 40.765 191.245 ;
        RECT 36.035 190.545 37.105 190.715 ;
        RECT 37.350 190.335 37.655 190.795 ;
        RECT 37.825 190.515 38.080 191.045 ;
        RECT 39.375 190.965 40.765 191.155 ;
        RECT 39.375 190.605 39.705 190.965 ;
        RECT 41.055 190.795 41.305 192.165 ;
        RECT 41.475 191.720 41.765 192.885 ;
        RECT 41.940 191.745 42.275 192.715 ;
        RECT 42.445 191.745 42.615 192.885 ;
        RECT 42.785 192.545 44.815 192.715 ;
        RECT 41.940 191.075 42.110 191.745 ;
        RECT 42.785 191.575 42.955 192.545 ;
        RECT 42.280 191.245 42.535 191.575 ;
        RECT 42.760 191.245 42.955 191.575 ;
        RECT 43.125 192.205 44.250 192.375 ;
        RECT 42.365 191.075 42.535 191.245 ;
        RECT 43.125 191.075 43.295 192.205 ;
        RECT 40.325 190.335 40.575 190.795 ;
        RECT 40.745 190.505 41.305 190.795 ;
        RECT 41.475 190.335 41.765 191.060 ;
        RECT 41.940 190.505 42.195 191.075 ;
        RECT 42.365 190.905 43.295 191.075 ;
        RECT 43.465 191.865 44.475 192.035 ;
        RECT 43.465 191.065 43.635 191.865 ;
        RECT 43.120 190.870 43.295 190.905 ;
        RECT 42.365 190.335 42.695 190.735 ;
        RECT 43.120 190.505 43.650 190.870 ;
        RECT 43.840 190.845 44.115 191.665 ;
        RECT 43.835 190.675 44.115 190.845 ;
        RECT 43.840 190.505 44.115 190.675 ;
        RECT 44.285 190.505 44.475 191.865 ;
        RECT 44.645 191.880 44.815 192.545 ;
        RECT 44.985 192.125 45.155 192.885 ;
        RECT 45.390 192.125 45.905 192.535 ;
        RECT 46.080 192.460 46.415 192.885 ;
        RECT 46.585 192.280 46.770 192.685 ;
        RECT 44.645 191.690 45.395 191.880 ;
        RECT 45.565 191.315 45.905 192.125 ;
        RECT 44.675 191.145 45.905 191.315 ;
        RECT 46.105 192.105 46.770 192.280 ;
        RECT 46.975 192.105 47.305 192.885 ;
        RECT 44.655 190.335 45.165 190.870 ;
        RECT 45.385 190.540 45.630 191.145 ;
        RECT 46.105 191.075 46.445 192.105 ;
        RECT 47.475 191.915 47.745 192.685 ;
        RECT 47.920 192.215 48.175 192.715 ;
        RECT 48.345 192.385 48.675 192.885 ;
        RECT 47.920 192.045 48.670 192.215 ;
        RECT 46.615 191.745 47.745 191.915 ;
        RECT 46.615 191.245 46.865 191.745 ;
        RECT 46.105 190.905 46.790 191.075 ;
        RECT 47.045 190.995 47.405 191.575 ;
        RECT 46.080 190.335 46.415 190.735 ;
        RECT 46.585 190.505 46.790 190.905 ;
        RECT 47.575 190.835 47.745 191.745 ;
        RECT 47.920 191.225 48.270 191.875 ;
        RECT 48.440 191.055 48.670 192.045 ;
        RECT 47.000 190.335 47.275 190.815 ;
        RECT 47.485 190.505 47.745 190.835 ;
        RECT 47.920 190.885 48.670 191.055 ;
        RECT 47.920 190.595 48.175 190.885 ;
        RECT 48.345 190.335 48.675 190.715 ;
        RECT 48.845 190.595 49.015 192.715 ;
        RECT 49.185 191.915 49.510 192.700 ;
        RECT 49.680 192.425 49.930 192.885 ;
        RECT 50.100 192.385 50.350 192.715 ;
        RECT 50.565 192.385 51.245 192.715 ;
        RECT 50.100 192.255 50.270 192.385 ;
        RECT 49.875 192.085 50.270 192.255 ;
        RECT 49.245 190.865 49.705 191.915 ;
        RECT 49.875 190.725 50.045 192.085 ;
        RECT 50.440 191.825 50.905 192.215 ;
        RECT 50.215 191.015 50.565 191.635 ;
        RECT 50.735 191.235 50.905 191.825 ;
        RECT 51.075 191.605 51.245 192.385 ;
        RECT 51.415 192.285 51.585 192.625 ;
        RECT 51.820 192.455 52.150 192.885 ;
        RECT 52.320 192.285 52.490 192.625 ;
        RECT 52.785 192.425 53.155 192.885 ;
        RECT 51.415 192.115 52.490 192.285 ;
        RECT 53.325 192.255 53.495 192.715 ;
        RECT 53.730 192.375 54.600 192.715 ;
        RECT 54.770 192.425 55.020 192.885 ;
        RECT 52.935 192.085 53.495 192.255 ;
        RECT 52.935 191.945 53.105 192.085 ;
        RECT 51.605 191.775 53.105 191.945 ;
        RECT 53.800 191.915 54.260 192.205 ;
        RECT 51.075 191.435 52.765 191.605 ;
        RECT 50.735 191.015 51.090 191.235 ;
        RECT 51.260 190.725 51.430 191.435 ;
        RECT 51.635 191.015 52.425 191.265 ;
        RECT 52.595 191.255 52.765 191.435 ;
        RECT 52.935 191.085 53.105 191.775 ;
        RECT 49.375 190.335 49.705 190.695 ;
        RECT 49.875 190.555 50.370 190.725 ;
        RECT 50.575 190.555 51.430 190.725 ;
        RECT 52.305 190.335 52.635 190.795 ;
        RECT 52.845 190.695 53.105 191.085 ;
        RECT 53.295 191.905 54.260 191.915 ;
        RECT 54.430 191.995 54.600 192.375 ;
        RECT 55.190 192.335 55.360 192.625 ;
        RECT 55.540 192.505 55.870 192.885 ;
        RECT 55.190 192.165 55.990 192.335 ;
        RECT 53.295 191.745 53.970 191.905 ;
        RECT 54.430 191.825 55.650 191.995 ;
        RECT 53.295 190.955 53.505 191.745 ;
        RECT 54.430 191.735 54.600 191.825 ;
        RECT 53.675 190.955 54.025 191.575 ;
        RECT 54.195 191.565 54.600 191.735 ;
        RECT 54.195 190.785 54.365 191.565 ;
        RECT 54.535 191.115 54.755 191.395 ;
        RECT 54.935 191.285 55.475 191.655 ;
        RECT 55.820 191.575 55.990 192.165 ;
        RECT 56.210 191.745 56.515 192.885 ;
        RECT 56.685 191.695 56.940 192.575 ;
        RECT 55.820 191.545 56.560 191.575 ;
        RECT 54.535 190.945 55.065 191.115 ;
        RECT 52.845 190.525 53.195 190.695 ;
        RECT 53.415 190.505 54.365 190.785 ;
        RECT 54.535 190.335 54.725 190.775 ;
        RECT 54.895 190.715 55.065 190.945 ;
        RECT 55.235 190.885 55.475 191.285 ;
        RECT 55.645 191.245 56.560 191.545 ;
        RECT 55.645 191.070 55.970 191.245 ;
        RECT 55.645 190.715 55.965 191.070 ;
        RECT 56.730 191.045 56.940 191.695 ;
        RECT 54.895 190.545 55.965 190.715 ;
        RECT 56.210 190.335 56.515 190.795 ;
        RECT 56.685 190.515 56.940 191.045 ;
        RECT 57.120 191.745 57.455 192.715 ;
        RECT 57.625 191.745 57.795 192.885 ;
        RECT 57.965 192.545 59.995 192.715 ;
        RECT 57.120 191.075 57.290 191.745 ;
        RECT 57.965 191.575 58.135 192.545 ;
        RECT 57.460 191.245 57.715 191.575 ;
        RECT 57.940 191.245 58.135 191.575 ;
        RECT 58.305 192.205 59.430 192.375 ;
        RECT 57.545 191.075 57.715 191.245 ;
        RECT 58.305 191.075 58.475 192.205 ;
        RECT 57.120 190.505 57.375 191.075 ;
        RECT 57.545 190.905 58.475 191.075 ;
        RECT 58.645 191.865 59.655 192.035 ;
        RECT 58.645 191.065 58.815 191.865 ;
        RECT 59.020 191.525 59.295 191.665 ;
        RECT 59.015 191.355 59.295 191.525 ;
        RECT 58.300 190.870 58.475 190.905 ;
        RECT 57.545 190.335 57.875 190.735 ;
        RECT 58.300 190.505 58.830 190.870 ;
        RECT 59.020 190.505 59.295 191.355 ;
        RECT 59.465 190.505 59.655 191.865 ;
        RECT 59.825 191.880 59.995 192.545 ;
        RECT 60.165 192.125 60.335 192.885 ;
        RECT 60.570 192.125 61.085 192.535 ;
        RECT 59.825 191.690 60.575 191.880 ;
        RECT 60.745 191.315 61.085 192.125 ;
        RECT 61.265 191.915 61.595 192.700 ;
        RECT 61.265 191.745 61.945 191.915 ;
        RECT 62.125 191.745 62.455 192.885 ;
        RECT 63.555 191.745 63.815 192.715 ;
        RECT 64.010 192.475 64.340 192.885 ;
        RECT 64.540 192.295 64.710 192.715 ;
        RECT 64.925 192.475 65.595 192.885 ;
        RECT 65.830 192.295 66.000 192.715 ;
        RECT 66.305 192.445 66.635 192.885 ;
        RECT 63.985 192.125 66.000 192.295 ;
        RECT 66.805 192.265 66.980 192.715 ;
        RECT 61.255 191.325 61.605 191.575 ;
        RECT 59.855 191.145 61.085 191.315 ;
        RECT 61.775 191.145 61.945 191.745 ;
        RECT 62.115 191.325 62.465 191.575 ;
        RECT 59.835 190.335 60.345 190.870 ;
        RECT 60.565 190.540 60.810 191.145 ;
        RECT 61.275 190.335 61.515 191.145 ;
        RECT 61.685 190.505 62.015 191.145 ;
        RECT 62.185 190.335 62.455 191.145 ;
        RECT 63.555 191.055 63.725 191.745 ;
        RECT 63.985 191.575 64.155 192.125 ;
        RECT 63.895 191.245 64.155 191.575 ;
        RECT 63.555 190.590 63.895 191.055 ;
        RECT 64.325 190.915 64.665 191.945 ;
        RECT 64.855 190.845 65.125 191.945 ;
        RECT 63.560 190.545 63.895 190.590 ;
        RECT 64.065 190.335 64.395 190.715 ;
        RECT 64.855 190.675 65.165 190.845 ;
        RECT 64.855 190.670 65.125 190.675 ;
        RECT 65.350 190.670 65.630 191.945 ;
        RECT 65.830 190.835 66.000 192.125 ;
        RECT 66.350 192.095 66.980 192.265 ;
        RECT 66.350 191.575 66.520 192.095 ;
        RECT 66.170 191.245 66.520 191.575 ;
        RECT 66.700 191.245 67.065 191.925 ;
        RECT 67.235 191.720 67.525 192.885 ;
        RECT 67.695 191.795 71.205 192.885 ;
        RECT 71.375 191.795 72.585 192.885 ;
        RECT 66.350 191.075 66.520 191.245 ;
        RECT 67.695 191.105 69.345 191.625 ;
        RECT 69.515 191.275 71.205 191.795 ;
        RECT 66.350 190.905 66.980 191.075 ;
        RECT 65.830 190.505 66.060 190.835 ;
        RECT 66.305 190.335 66.635 190.715 ;
        RECT 66.805 190.505 66.980 190.905 ;
        RECT 67.235 190.335 67.525 191.060 ;
        RECT 67.695 190.335 71.205 191.105 ;
        RECT 71.375 191.085 71.895 191.625 ;
        RECT 72.065 191.255 72.585 191.795 ;
        RECT 72.755 191.745 73.015 192.885 ;
        RECT 73.185 191.735 73.515 192.715 ;
        RECT 73.685 191.745 73.965 192.885 ;
        RECT 74.145 191.915 74.475 192.700 ;
        RECT 74.145 191.745 74.825 191.915 ;
        RECT 75.005 191.745 75.335 192.885 ;
        RECT 75.515 192.450 80.860 192.885 ;
        RECT 72.775 191.325 73.110 191.575 ;
        RECT 73.280 191.135 73.450 191.735 ;
        RECT 73.620 191.305 73.955 191.575 ;
        RECT 74.135 191.325 74.485 191.575 ;
        RECT 74.655 191.145 74.825 191.745 ;
        RECT 74.995 191.325 75.345 191.575 ;
        RECT 71.375 190.335 72.585 191.085 ;
        RECT 72.755 190.505 73.450 191.135 ;
        RECT 73.655 190.335 73.965 191.135 ;
        RECT 74.155 190.335 74.395 191.145 ;
        RECT 74.565 190.505 74.895 191.145 ;
        RECT 75.065 190.335 75.335 191.145 ;
        RECT 77.100 190.880 77.440 191.710 ;
        RECT 78.920 191.200 79.270 192.450 ;
        RECT 81.035 191.795 84.545 192.885 ;
        RECT 84.715 191.795 85.925 192.885 ;
        RECT 81.035 191.105 82.685 191.625 ;
        RECT 82.855 191.275 84.545 191.795 ;
        RECT 75.515 190.335 80.860 190.880 ;
        RECT 81.035 190.335 84.545 191.105 ;
        RECT 84.715 191.085 85.235 191.625 ;
        RECT 85.405 191.255 85.925 191.795 ;
        RECT 86.095 191.745 86.385 192.885 ;
        RECT 87.180 192.545 88.545 192.715 ;
        RECT 87.180 192.335 87.510 192.545 ;
        RECT 86.555 192.085 87.510 192.335 ;
        RECT 86.095 191.245 86.370 191.575 ;
        RECT 84.715 190.335 85.925 191.085 ;
        RECT 86.555 191.075 86.725 192.085 ;
        RECT 86.895 191.245 87.250 191.910 ;
        RECT 87.435 191.245 87.710 191.910 ;
        RECT 87.880 191.575 88.205 192.375 ;
        RECT 88.375 191.915 88.545 192.545 ;
        RECT 88.715 192.085 89.005 192.885 ;
        RECT 88.375 191.745 89.050 191.915 ;
        RECT 89.220 191.745 89.605 192.705 ;
        RECT 89.775 191.795 92.365 192.885 ;
        RECT 88.880 191.575 89.050 191.745 ;
        RECT 87.880 191.245 88.225 191.575 ;
        RECT 88.435 191.325 88.685 191.575 ;
        RECT 88.880 191.325 89.245 191.575 ;
        RECT 88.515 191.245 88.685 191.325 ;
        RECT 89.055 191.245 89.245 191.325 ;
        RECT 89.430 191.075 89.605 191.745 ;
        RECT 86.095 190.715 86.385 190.985 ;
        RECT 86.555 190.885 86.980 191.075 ;
        RECT 87.150 190.905 88.550 191.075 ;
        RECT 87.150 190.715 87.480 190.905 ;
        RECT 86.095 190.505 87.480 190.715 ;
        RECT 87.715 190.335 88.045 190.735 ;
        RECT 88.220 190.505 88.550 190.905 ;
        RECT 88.755 190.335 88.925 190.895 ;
        RECT 89.095 190.505 89.605 191.075 ;
        RECT 89.775 191.105 90.985 191.625 ;
        RECT 91.155 191.275 92.365 191.795 ;
        RECT 92.995 191.720 93.285 192.885 ;
        RECT 93.660 191.915 93.990 192.715 ;
        RECT 94.160 192.085 94.490 192.885 ;
        RECT 94.790 191.915 95.120 192.715 ;
        RECT 95.765 192.085 96.015 192.885 ;
        RECT 93.660 191.745 96.095 191.915 ;
        RECT 96.285 191.745 96.455 192.885 ;
        RECT 96.625 191.745 96.965 192.715 ;
        RECT 93.455 191.325 93.805 191.575 ;
        RECT 93.990 191.115 94.160 191.745 ;
        RECT 94.330 191.325 94.660 191.525 ;
        RECT 94.830 191.325 95.160 191.525 ;
        RECT 95.330 191.325 95.750 191.525 ;
        RECT 95.925 191.495 96.095 191.745 ;
        RECT 95.925 191.325 96.620 191.495 ;
        RECT 89.775 190.335 92.365 191.105 ;
        RECT 92.995 190.335 93.285 191.060 ;
        RECT 93.660 190.505 94.160 191.115 ;
        RECT 94.790 190.985 96.015 191.155 ;
        RECT 96.790 191.135 96.965 191.745 ;
        RECT 94.790 190.505 95.120 190.985 ;
        RECT 95.290 190.335 95.515 190.795 ;
        RECT 95.685 190.505 96.015 190.985 ;
        RECT 96.205 190.335 96.455 191.135 ;
        RECT 96.625 190.505 96.965 191.135 ;
        RECT 97.140 192.165 97.475 192.675 ;
        RECT 97.140 190.810 97.395 192.165 ;
        RECT 97.725 192.085 98.055 192.885 ;
        RECT 98.300 192.295 98.585 192.715 ;
        RECT 98.840 192.465 99.170 192.885 ;
        RECT 99.395 192.545 100.555 192.715 ;
        RECT 99.395 192.295 99.725 192.545 ;
        RECT 98.300 192.125 99.725 192.295 ;
        RECT 99.955 191.915 100.125 192.375 ;
        RECT 100.385 192.045 100.555 192.545 ;
        RECT 97.755 191.745 100.125 191.915 ;
        RECT 97.755 191.575 97.925 191.745 ;
        RECT 100.375 191.695 100.585 191.865 ;
        RECT 100.815 191.795 102.025 192.885 ;
        RECT 100.375 191.575 100.580 191.695 ;
        RECT 97.620 191.245 97.925 191.575 ;
        RECT 98.120 191.245 98.370 191.575 ;
        RECT 98.580 191.525 98.850 191.575 ;
        RECT 99.040 191.525 99.330 191.575 ;
        RECT 98.575 191.355 98.850 191.525 ;
        RECT 99.035 191.355 99.330 191.525 ;
        RECT 97.755 191.075 97.925 191.245 ;
        RECT 97.755 190.905 98.315 191.075 ;
        RECT 98.580 190.915 98.850 191.355 ;
        RECT 99.040 190.915 99.330 191.355 ;
        RECT 99.500 190.910 99.920 191.575 ;
        RECT 100.230 191.245 100.580 191.575 ;
        RECT 100.815 191.085 101.335 191.625 ;
        RECT 101.505 191.255 102.025 191.795 ;
        RECT 102.195 191.745 102.455 192.885 ;
        RECT 102.625 191.915 102.955 192.715 ;
        RECT 103.125 192.085 103.295 192.885 ;
        RECT 103.465 191.915 103.795 192.715 ;
        RECT 103.965 192.085 104.220 192.885 ;
        RECT 102.625 191.745 104.325 191.915 ;
        RECT 104.495 191.795 105.705 192.885 ;
        RECT 105.880 192.375 107.535 192.665 ;
        RECT 102.195 191.325 102.955 191.575 ;
        RECT 103.125 191.325 103.875 191.575 ;
        RECT 104.045 191.155 104.325 191.745 ;
        RECT 97.140 190.550 97.475 190.810 ;
        RECT 98.145 190.735 98.315 190.905 ;
        RECT 97.645 190.335 97.975 190.735 ;
        RECT 98.145 190.565 99.760 190.735 ;
        RECT 100.305 190.335 100.635 191.055 ;
        RECT 100.815 190.335 102.025 191.085 ;
        RECT 102.195 190.965 103.295 191.135 ;
        RECT 102.195 190.505 102.535 190.965 ;
        RECT 102.705 190.335 102.875 190.795 ;
        RECT 103.045 190.715 103.295 190.965 ;
        RECT 103.465 190.905 104.325 191.155 ;
        RECT 104.495 191.085 105.015 191.625 ;
        RECT 105.185 191.255 105.705 191.795 ;
        RECT 105.880 192.035 107.470 192.205 ;
        RECT 107.705 192.085 107.985 192.885 ;
        RECT 105.880 191.745 106.200 192.035 ;
        RECT 107.300 191.915 107.470 192.035 ;
        RECT 106.395 191.695 107.110 191.865 ;
        RECT 107.300 191.745 108.025 191.915 ;
        RECT 108.195 191.745 108.465 192.715 ;
        RECT 108.635 191.795 112.145 192.885 ;
        RECT 103.885 190.715 104.215 190.735 ;
        RECT 103.045 190.505 104.215 190.715 ;
        RECT 104.495 190.335 105.705 191.085 ;
        RECT 105.880 191.005 106.230 191.575 ;
        RECT 106.400 191.245 107.110 191.695 ;
        RECT 107.855 191.575 108.025 191.745 ;
        RECT 107.280 191.245 107.685 191.575 ;
        RECT 107.855 191.245 108.125 191.575 ;
        RECT 107.855 191.075 108.025 191.245 ;
        RECT 106.415 190.905 108.025 191.075 ;
        RECT 108.295 191.010 108.465 191.745 ;
        RECT 105.885 190.335 106.215 190.835 ;
        RECT 106.415 190.555 106.585 190.905 ;
        RECT 106.785 190.335 107.115 190.735 ;
        RECT 107.285 190.555 107.455 190.905 ;
        RECT 107.625 190.335 108.005 190.735 ;
        RECT 108.195 190.665 108.465 191.010 ;
        RECT 108.635 191.105 110.285 191.625 ;
        RECT 110.455 191.275 112.145 191.795 ;
        RECT 112.780 191.745 113.110 192.885 ;
        RECT 113.280 192.255 113.455 192.665 ;
        RECT 113.625 192.425 113.955 192.885 ;
        RECT 114.160 192.255 114.385 192.665 ;
        RECT 113.280 192.085 114.385 192.255 ;
        RECT 114.565 191.915 114.900 192.695 ;
        RECT 113.760 191.865 114.145 191.915 ;
        RECT 113.755 191.695 114.145 191.865 ;
        RECT 112.775 191.245 113.055 191.575 ;
        RECT 113.300 191.185 113.745 191.525 ;
        RECT 113.960 191.245 114.145 191.695 ;
        RECT 114.315 191.745 114.900 191.915 ;
        RECT 115.075 191.795 118.585 192.885 ;
        RECT 108.635 190.335 112.145 191.105 ;
        RECT 112.780 190.335 113.120 191.065 ;
        RECT 113.295 191.015 113.745 191.185 ;
        RECT 114.315 191.075 114.485 191.745 ;
        RECT 114.655 191.245 114.905 191.575 ;
        RECT 113.300 190.585 113.745 191.015 ;
        RECT 114.070 190.965 114.485 191.075 ;
        RECT 115.075 191.105 116.725 191.625 ;
        RECT 116.895 191.275 118.585 191.795 ;
        RECT 118.755 191.720 119.045 192.885 ;
        RECT 119.215 191.745 119.485 192.715 ;
        RECT 119.695 192.085 119.975 192.885 ;
        RECT 120.145 192.375 121.800 192.665 ;
        RECT 121.975 192.450 127.320 192.885 ;
        RECT 127.495 192.450 132.840 192.885 ;
        RECT 120.210 192.035 121.800 192.205 ;
        RECT 120.210 191.915 120.380 192.035 ;
        RECT 119.655 191.745 120.380 191.915 ;
        RECT 114.070 190.545 114.475 190.965 ;
        RECT 114.645 190.335 114.905 190.815 ;
        RECT 115.075 190.335 118.585 191.105 ;
        RECT 118.755 190.335 119.045 191.060 ;
        RECT 119.215 191.010 119.385 191.745 ;
        RECT 119.655 191.575 119.825 191.745 ;
        RECT 119.555 191.245 119.825 191.575 ;
        RECT 119.995 191.245 120.400 191.575 ;
        RECT 120.570 191.245 121.280 191.865 ;
        RECT 121.480 191.745 121.800 192.035 ;
        RECT 119.655 191.075 119.825 191.245 ;
        RECT 119.215 190.665 119.485 191.010 ;
        RECT 119.655 190.905 121.265 191.075 ;
        RECT 121.450 191.005 121.800 191.575 ;
        RECT 119.675 190.335 120.055 190.735 ;
        RECT 120.225 190.555 120.395 190.905 ;
        RECT 120.565 190.335 120.895 190.735 ;
        RECT 121.095 190.555 121.265 190.905 ;
        RECT 123.560 190.880 123.900 191.710 ;
        RECT 125.380 191.200 125.730 192.450 ;
        RECT 129.080 190.880 129.420 191.710 ;
        RECT 130.900 191.200 131.250 192.450 ;
        RECT 133.015 191.795 134.685 192.885 ;
        RECT 133.015 191.105 133.765 191.625 ;
        RECT 133.935 191.275 134.685 191.795 ;
        RECT 134.860 191.745 135.115 192.885 ;
        RECT 135.285 191.845 135.595 192.715 ;
        RECT 135.795 192.425 136.085 192.885 ;
        RECT 136.255 192.505 137.565 192.675 ;
        RECT 136.255 192.255 136.425 192.505 ;
        RECT 138.095 192.425 138.315 192.885 ;
        RECT 138.485 192.255 138.820 192.715 ;
        RECT 138.995 192.450 144.340 192.885 ;
        RECT 135.765 192.085 136.425 192.255 ;
        RECT 136.595 192.085 138.820 192.255 ;
        RECT 121.465 190.335 121.795 190.835 ;
        RECT 121.975 190.335 127.320 190.880 ;
        RECT 127.495 190.335 132.840 190.880 ;
        RECT 133.015 190.335 134.685 191.105 ;
        RECT 134.860 190.335 135.115 191.135 ;
        RECT 135.285 191.000 135.455 191.845 ;
        RECT 135.765 191.575 135.935 192.085 ;
        RECT 136.595 191.915 136.765 192.085 ;
        RECT 135.625 191.245 135.935 191.575 ;
        RECT 136.105 191.745 136.765 191.915 ;
        RECT 136.105 191.245 136.275 191.745 ;
        RECT 137.045 191.565 137.860 191.875 ;
        RECT 137.045 191.530 137.215 191.565 ;
        RECT 135.765 191.055 135.935 191.245 ;
        RECT 135.285 190.505 135.535 191.000 ;
        RECT 135.765 190.885 136.375 191.055 ;
        RECT 136.585 191.015 137.215 191.530 ;
        RECT 137.395 190.985 137.860 191.275 ;
        RECT 138.130 191.005 138.320 191.875 ;
        RECT 136.205 190.715 136.375 190.885 ;
        RECT 135.705 190.335 136.035 190.715 ;
        RECT 136.205 190.545 137.500 190.715 ;
        RECT 137.670 190.670 137.860 190.985 ;
        RECT 138.120 190.335 138.320 190.835 ;
        RECT 138.490 190.505 138.820 192.085 ;
        RECT 140.580 190.880 140.920 191.710 ;
        RECT 142.400 191.200 142.750 192.450 ;
        RECT 144.515 191.720 144.805 192.885 ;
        RECT 144.975 192.450 150.320 192.885 ;
        RECT 138.995 190.335 144.340 190.880 ;
        RECT 144.515 190.335 144.805 191.060 ;
        RECT 146.560 190.880 146.900 191.710 ;
        RECT 148.380 191.200 148.730 192.450 ;
        RECT 150.955 191.745 151.225 192.715 ;
        RECT 151.435 192.085 151.715 192.885 ;
        RECT 151.885 192.375 153.540 192.665 ;
        RECT 151.950 192.035 153.540 192.205 ;
        RECT 151.950 191.915 152.120 192.035 ;
        RECT 151.395 191.745 152.120 191.915 ;
        RECT 150.955 191.010 151.125 191.745 ;
        RECT 151.395 191.575 151.565 191.745 ;
        RECT 151.295 191.245 151.565 191.575 ;
        RECT 151.735 191.245 152.140 191.575 ;
        RECT 152.310 191.245 153.020 191.865 ;
        RECT 153.220 191.745 153.540 192.035 ;
        RECT 153.715 191.795 156.305 192.885 ;
        RECT 151.395 191.075 151.565 191.245 ;
        RECT 144.975 190.335 150.320 190.880 ;
        RECT 150.955 190.665 151.225 191.010 ;
        RECT 151.395 190.905 153.005 191.075 ;
        RECT 153.190 191.005 153.540 191.575 ;
        RECT 153.715 191.105 154.925 191.625 ;
        RECT 155.095 191.275 156.305 191.795 ;
        RECT 156.935 191.795 158.145 192.885 ;
        RECT 156.935 191.255 157.455 191.795 ;
        RECT 151.415 190.335 151.795 190.735 ;
        RECT 151.965 190.555 152.135 190.905 ;
        RECT 152.305 190.335 152.635 190.735 ;
        RECT 152.835 190.555 153.005 190.905 ;
        RECT 153.205 190.335 153.535 190.835 ;
        RECT 153.715 190.335 156.305 191.105 ;
        RECT 157.625 191.085 158.145 191.625 ;
        RECT 156.935 190.335 158.145 191.085 ;
        RECT 2.750 190.165 158.230 190.335 ;
        RECT 2.835 189.415 4.045 190.165 ;
        RECT 4.765 189.615 4.935 189.995 ;
        RECT 5.115 189.785 5.445 190.165 ;
        RECT 4.765 189.445 5.430 189.615 ;
        RECT 5.625 189.490 5.885 189.995 ;
        RECT 2.835 188.875 3.355 189.415 ;
        RECT 3.525 188.705 4.045 189.245 ;
        RECT 4.695 188.895 5.025 189.265 ;
        RECT 5.260 189.190 5.430 189.445 ;
        RECT 5.260 188.860 5.545 189.190 ;
        RECT 5.260 188.715 5.430 188.860 ;
        RECT 2.835 187.615 4.045 188.705 ;
        RECT 4.765 188.545 5.430 188.715 ;
        RECT 5.715 188.690 5.885 189.490 ;
        RECT 6.060 189.615 6.315 189.905 ;
        RECT 6.485 189.785 6.815 190.165 ;
        RECT 6.060 189.445 6.810 189.615 ;
        RECT 4.765 187.785 4.935 188.545 ;
        RECT 5.115 187.615 5.445 188.375 ;
        RECT 5.615 187.785 5.885 188.690 ;
        RECT 6.060 188.625 6.410 189.275 ;
        RECT 6.580 188.455 6.810 189.445 ;
        RECT 6.060 188.285 6.810 188.455 ;
        RECT 6.060 187.785 6.315 188.285 ;
        RECT 6.485 187.615 6.815 188.115 ;
        RECT 6.985 187.785 7.155 189.905 ;
        RECT 7.515 189.805 7.845 190.165 ;
        RECT 8.015 189.775 8.510 189.945 ;
        RECT 8.715 189.775 9.570 189.945 ;
        RECT 7.385 188.585 7.845 189.635 ;
        RECT 7.325 187.800 7.650 188.585 ;
        RECT 8.015 188.415 8.185 189.775 ;
        RECT 8.355 188.865 8.705 189.485 ;
        RECT 8.875 189.265 9.230 189.485 ;
        RECT 8.875 188.675 9.045 189.265 ;
        RECT 9.400 189.065 9.570 189.775 ;
        RECT 10.445 189.705 10.775 190.165 ;
        RECT 10.985 189.805 11.335 189.975 ;
        RECT 9.775 189.235 10.565 189.485 ;
        RECT 10.985 189.415 11.245 189.805 ;
        RECT 11.555 189.715 12.505 189.995 ;
        RECT 12.675 189.725 12.865 190.165 ;
        RECT 13.035 189.785 14.105 189.955 ;
        RECT 10.735 189.065 10.905 189.245 ;
        RECT 8.015 188.245 8.410 188.415 ;
        RECT 8.580 188.285 9.045 188.675 ;
        RECT 9.215 188.895 10.905 189.065 ;
        RECT 8.240 188.115 8.410 188.245 ;
        RECT 9.215 188.115 9.385 188.895 ;
        RECT 11.075 188.725 11.245 189.415 ;
        RECT 9.745 188.555 11.245 188.725 ;
        RECT 11.435 188.755 11.645 189.545 ;
        RECT 11.815 188.925 12.165 189.545 ;
        RECT 12.335 188.935 12.505 189.715 ;
        RECT 13.035 189.555 13.205 189.785 ;
        RECT 12.675 189.385 13.205 189.555 ;
        RECT 12.675 189.105 12.895 189.385 ;
        RECT 13.375 189.215 13.615 189.615 ;
        RECT 12.335 188.765 12.740 188.935 ;
        RECT 13.075 188.845 13.615 189.215 ;
        RECT 13.785 189.430 14.105 189.785 ;
        RECT 14.350 189.705 14.655 190.165 ;
        RECT 14.825 189.455 15.080 189.985 ;
        RECT 13.785 189.255 14.110 189.430 ;
        RECT 13.785 188.955 14.700 189.255 ;
        RECT 13.960 188.925 14.700 188.955 ;
        RECT 11.435 188.595 12.110 188.755 ;
        RECT 12.570 188.675 12.740 188.765 ;
        RECT 11.435 188.585 12.400 188.595 ;
        RECT 11.075 188.415 11.245 188.555 ;
        RECT 7.820 187.615 8.070 188.075 ;
        RECT 8.240 187.785 8.490 188.115 ;
        RECT 8.705 187.785 9.385 188.115 ;
        RECT 9.555 188.215 10.630 188.385 ;
        RECT 11.075 188.245 11.635 188.415 ;
        RECT 11.940 188.295 12.400 188.585 ;
        RECT 12.570 188.505 13.790 188.675 ;
        RECT 9.555 187.875 9.725 188.215 ;
        RECT 9.960 187.615 10.290 188.045 ;
        RECT 10.460 187.875 10.630 188.215 ;
        RECT 10.925 187.615 11.295 188.075 ;
        RECT 11.465 187.785 11.635 188.245 ;
        RECT 12.570 188.125 12.740 188.505 ;
        RECT 13.960 188.335 14.130 188.925 ;
        RECT 14.870 188.805 15.080 189.455 ;
        RECT 15.805 189.615 15.975 189.995 ;
        RECT 16.155 189.785 16.485 190.165 ;
        RECT 15.805 189.445 16.470 189.615 ;
        RECT 16.665 189.490 16.925 189.995 ;
        RECT 15.735 188.895 16.065 189.265 ;
        RECT 16.300 189.190 16.470 189.445 ;
        RECT 11.870 187.785 12.740 188.125 ;
        RECT 13.330 188.165 14.130 188.335 ;
        RECT 12.910 187.615 13.160 188.075 ;
        RECT 13.330 187.875 13.500 188.165 ;
        RECT 13.680 187.615 14.010 187.995 ;
        RECT 14.350 187.615 14.655 188.755 ;
        RECT 14.825 187.925 15.080 188.805 ;
        RECT 16.300 188.860 16.585 189.190 ;
        RECT 16.300 188.715 16.470 188.860 ;
        RECT 15.805 188.545 16.470 188.715 ;
        RECT 16.755 188.690 16.925 189.490 ;
        RECT 17.100 189.615 17.355 189.905 ;
        RECT 17.525 189.785 17.855 190.165 ;
        RECT 17.100 189.445 17.850 189.615 ;
        RECT 15.805 187.785 15.975 188.545 ;
        RECT 16.155 187.615 16.485 188.375 ;
        RECT 16.655 187.785 16.925 188.690 ;
        RECT 17.100 188.625 17.450 189.275 ;
        RECT 17.620 188.455 17.850 189.445 ;
        RECT 17.100 188.285 17.850 188.455 ;
        RECT 17.100 187.785 17.355 188.285 ;
        RECT 17.525 187.615 17.855 188.115 ;
        RECT 18.025 187.785 18.195 189.905 ;
        RECT 18.555 189.805 18.885 190.165 ;
        RECT 19.055 189.775 19.550 189.945 ;
        RECT 19.755 189.775 20.610 189.945 ;
        RECT 18.425 188.585 18.885 189.635 ;
        RECT 18.365 187.800 18.690 188.585 ;
        RECT 19.055 188.415 19.225 189.775 ;
        RECT 19.395 188.865 19.745 189.485 ;
        RECT 19.915 189.265 20.270 189.485 ;
        RECT 19.915 188.675 20.085 189.265 ;
        RECT 20.440 189.065 20.610 189.775 ;
        RECT 21.485 189.705 21.815 190.165 ;
        RECT 22.025 189.805 22.375 189.975 ;
        RECT 20.815 189.235 21.605 189.485 ;
        RECT 22.025 189.415 22.285 189.805 ;
        RECT 22.595 189.715 23.545 189.995 ;
        RECT 23.715 189.725 23.905 190.165 ;
        RECT 24.075 189.785 25.145 189.955 ;
        RECT 21.775 189.065 21.945 189.245 ;
        RECT 19.055 188.245 19.450 188.415 ;
        RECT 19.620 188.285 20.085 188.675 ;
        RECT 20.255 188.895 21.945 189.065 ;
        RECT 19.280 188.115 19.450 188.245 ;
        RECT 20.255 188.115 20.425 188.895 ;
        RECT 22.115 188.725 22.285 189.415 ;
        RECT 20.785 188.555 22.285 188.725 ;
        RECT 22.475 188.755 22.685 189.545 ;
        RECT 22.855 188.925 23.205 189.545 ;
        RECT 23.375 188.935 23.545 189.715 ;
        RECT 24.075 189.555 24.245 189.785 ;
        RECT 23.715 189.385 24.245 189.555 ;
        RECT 23.715 189.105 23.935 189.385 ;
        RECT 24.415 189.215 24.655 189.615 ;
        RECT 23.375 188.765 23.780 188.935 ;
        RECT 24.115 188.845 24.655 189.215 ;
        RECT 24.825 189.430 25.145 189.785 ;
        RECT 25.390 189.705 25.695 190.165 ;
        RECT 25.865 189.455 26.115 189.985 ;
        RECT 24.825 189.255 25.150 189.430 ;
        RECT 24.825 188.955 25.740 189.255 ;
        RECT 25.000 188.925 25.740 188.955 ;
        RECT 22.475 188.595 23.150 188.755 ;
        RECT 23.610 188.675 23.780 188.765 ;
        RECT 22.475 188.585 23.440 188.595 ;
        RECT 22.115 188.415 22.285 188.555 ;
        RECT 18.860 187.615 19.110 188.075 ;
        RECT 19.280 187.785 19.530 188.115 ;
        RECT 19.745 187.785 20.425 188.115 ;
        RECT 20.595 188.215 21.670 188.385 ;
        RECT 22.115 188.245 22.675 188.415 ;
        RECT 22.980 188.295 23.440 188.585 ;
        RECT 23.610 188.505 24.830 188.675 ;
        RECT 20.595 187.875 20.765 188.215 ;
        RECT 21.000 187.615 21.330 188.045 ;
        RECT 21.500 187.875 21.670 188.215 ;
        RECT 21.965 187.615 22.335 188.075 ;
        RECT 22.505 187.785 22.675 188.245 ;
        RECT 23.610 188.125 23.780 188.505 ;
        RECT 25.000 188.335 25.170 188.925 ;
        RECT 25.910 188.805 26.115 189.455 ;
        RECT 26.285 189.410 26.535 190.165 ;
        RECT 26.755 189.395 28.425 190.165 ;
        RECT 28.595 189.440 28.885 190.165 ;
        RECT 29.055 189.395 31.645 190.165 ;
        RECT 26.755 188.875 27.505 189.395 ;
        RECT 22.910 187.785 23.780 188.125 ;
        RECT 24.370 188.165 25.170 188.335 ;
        RECT 23.950 187.615 24.200 188.075 ;
        RECT 24.370 187.875 24.540 188.165 ;
        RECT 24.720 187.615 25.050 187.995 ;
        RECT 25.390 187.615 25.695 188.755 ;
        RECT 25.865 187.925 26.115 188.805 ;
        RECT 26.285 187.615 26.535 188.755 ;
        RECT 27.675 188.705 28.425 189.225 ;
        RECT 29.055 188.875 30.265 189.395 ;
        RECT 32.285 189.355 32.555 190.165 ;
        RECT 32.725 189.355 33.055 189.995 ;
        RECT 33.225 189.355 33.465 190.165 ;
        RECT 33.660 189.765 33.995 190.165 ;
        RECT 34.165 189.595 34.370 189.995 ;
        RECT 34.580 189.685 34.855 190.165 ;
        RECT 35.065 189.665 35.325 189.995 ;
        RECT 36.505 189.685 36.805 190.165 ;
        RECT 33.685 189.425 34.370 189.595 ;
        RECT 26.755 187.615 28.425 188.705 ;
        RECT 28.595 187.615 28.885 188.780 ;
        RECT 30.435 188.705 31.645 189.225 ;
        RECT 32.275 188.925 32.625 189.175 ;
        RECT 32.795 188.755 32.965 189.355 ;
        RECT 33.135 188.925 33.485 189.175 ;
        RECT 29.055 187.615 31.645 188.705 ;
        RECT 32.285 187.615 32.615 188.755 ;
        RECT 32.795 188.585 33.475 188.755 ;
        RECT 33.145 187.800 33.475 188.585 ;
        RECT 33.685 188.395 34.025 189.425 ;
        RECT 34.195 188.755 34.445 189.255 ;
        RECT 34.625 188.925 34.985 189.505 ;
        RECT 35.155 188.755 35.325 189.665 ;
        RECT 36.975 189.515 37.235 189.970 ;
        RECT 37.405 189.685 37.665 190.165 ;
        RECT 37.845 189.515 38.105 189.970 ;
        RECT 38.275 189.685 38.525 190.165 ;
        RECT 38.705 189.515 38.965 189.970 ;
        RECT 39.135 189.685 39.385 190.165 ;
        RECT 39.565 189.515 39.825 189.970 ;
        RECT 39.995 189.685 40.240 190.165 ;
        RECT 40.410 189.515 40.685 189.970 ;
        RECT 40.855 189.685 41.100 190.165 ;
        RECT 41.270 189.515 41.530 189.970 ;
        RECT 41.700 189.685 41.960 190.165 ;
        RECT 42.130 189.515 42.390 189.970 ;
        RECT 42.560 189.685 42.820 190.165 ;
        RECT 42.990 189.515 43.250 189.970 ;
        RECT 43.420 189.605 43.680 190.165 ;
        RECT 36.505 189.485 43.250 189.515 ;
        RECT 36.475 189.345 43.250 189.485 ;
        RECT 36.475 189.315 37.670 189.345 ;
        RECT 34.195 188.585 35.325 188.755 ;
        RECT 33.685 188.220 34.350 188.395 ;
        RECT 33.660 187.615 33.995 188.040 ;
        RECT 34.165 187.815 34.350 188.220 ;
        RECT 34.555 187.615 34.885 188.395 ;
        RECT 35.055 187.815 35.325 188.585 ;
        RECT 36.505 188.755 37.670 189.315 ;
        RECT 43.850 189.175 44.100 189.985 ;
        RECT 44.280 189.640 44.540 190.165 ;
        RECT 44.710 189.175 44.960 189.985 ;
        RECT 45.140 189.655 45.445 190.165 ;
        RECT 37.840 188.925 44.960 189.175 ;
        RECT 45.130 188.925 45.445 189.485 ;
        RECT 45.615 189.345 46.300 189.985 ;
        RECT 46.470 189.345 46.640 190.165 ;
        RECT 46.810 189.515 47.140 189.980 ;
        RECT 47.310 189.695 47.480 190.165 ;
        RECT 47.740 189.775 48.925 189.945 ;
        RECT 49.095 189.605 49.425 189.995 ;
        RECT 48.125 189.515 48.510 189.605 ;
        RECT 46.810 189.345 48.510 189.515 ;
        RECT 48.915 189.425 49.425 189.605 ;
        RECT 50.790 189.535 51.075 189.995 ;
        RECT 51.245 189.705 51.515 190.165 ;
        RECT 36.505 188.530 43.250 188.755 ;
        RECT 36.505 187.615 36.775 188.360 ;
        RECT 36.945 187.790 37.235 188.530 ;
        RECT 37.845 188.515 43.250 188.530 ;
        RECT 37.405 187.620 37.660 188.345 ;
        RECT 37.845 187.790 38.105 188.515 ;
        RECT 38.275 187.620 38.520 188.345 ;
        RECT 38.705 187.790 38.965 188.515 ;
        RECT 39.135 187.620 39.380 188.345 ;
        RECT 39.565 187.790 39.825 188.515 ;
        RECT 39.995 187.620 40.240 188.345 ;
        RECT 40.410 187.790 40.670 188.515 ;
        RECT 40.840 187.620 41.100 188.345 ;
        RECT 41.270 187.790 41.530 188.515 ;
        RECT 41.700 187.620 41.960 188.345 ;
        RECT 42.130 187.790 42.390 188.515 ;
        RECT 42.560 187.620 42.820 188.345 ;
        RECT 42.990 187.790 43.250 188.515 ;
        RECT 43.420 187.620 43.680 188.415 ;
        RECT 43.850 187.790 44.100 188.925 ;
        RECT 37.405 187.615 43.680 187.620 ;
        RECT 44.280 187.615 44.540 188.425 ;
        RECT 44.715 187.785 44.960 188.925 ;
        RECT 45.140 187.615 45.435 188.425 ;
        RECT 45.615 188.375 45.865 189.345 ;
        RECT 46.035 188.965 46.370 189.175 ;
        RECT 46.540 188.965 46.990 189.175 ;
        RECT 47.180 188.965 47.665 189.175 ;
        RECT 46.200 188.795 46.370 188.965 ;
        RECT 47.290 188.805 47.665 188.965 ;
        RECT 47.855 188.925 48.235 189.175 ;
        RECT 48.415 188.965 48.745 189.175 ;
        RECT 46.200 188.625 47.120 188.795 ;
        RECT 45.615 187.785 46.280 188.375 ;
        RECT 46.450 187.615 46.780 188.455 ;
        RECT 46.950 188.375 47.120 188.625 ;
        RECT 47.290 188.635 47.685 188.805 ;
        RECT 47.290 188.545 47.665 188.635 ;
        RECT 47.855 188.545 48.175 188.925 ;
        RECT 48.915 188.795 49.085 189.425 ;
        RECT 50.790 189.365 51.745 189.535 ;
        RECT 49.255 188.965 49.585 189.255 ;
        RECT 48.345 188.625 49.430 188.795 ;
        RECT 50.675 188.635 51.365 189.195 ;
        RECT 48.345 188.375 48.515 188.625 ;
        RECT 46.950 188.205 48.515 188.375 ;
        RECT 47.290 187.785 48.095 188.205 ;
        RECT 48.685 187.615 48.935 188.455 ;
        RECT 49.130 187.785 49.430 188.625 ;
        RECT 51.535 188.465 51.745 189.365 ;
        RECT 50.790 188.245 51.745 188.465 ;
        RECT 51.915 189.195 52.315 189.995 ;
        RECT 52.505 189.535 52.785 189.995 ;
        RECT 53.305 189.705 53.630 190.165 ;
        RECT 52.505 189.365 53.630 189.535 ;
        RECT 53.800 189.425 54.185 189.995 ;
        RECT 54.355 189.440 54.645 190.165 ;
        RECT 53.180 189.255 53.630 189.365 ;
        RECT 51.915 188.635 53.010 189.195 ;
        RECT 53.180 188.925 53.735 189.255 ;
        RECT 50.790 187.785 51.075 188.245 ;
        RECT 51.245 187.615 51.515 188.075 ;
        RECT 51.915 187.785 52.315 188.635 ;
        RECT 53.180 188.465 53.630 188.925 ;
        RECT 53.905 188.755 54.185 189.425 ;
        RECT 54.835 189.355 55.075 190.165 ;
        RECT 55.245 189.355 55.575 189.995 ;
        RECT 55.745 189.355 56.015 190.165 ;
        RECT 56.470 189.355 56.715 189.960 ;
        RECT 56.935 189.630 57.445 190.165 ;
        RECT 54.815 188.925 55.165 189.175 ;
        RECT 52.505 188.245 53.630 188.465 ;
        RECT 52.505 187.785 52.785 188.245 ;
        RECT 53.305 187.615 53.630 188.075 ;
        RECT 53.800 187.785 54.185 188.755 ;
        RECT 54.355 187.615 54.645 188.780 ;
        RECT 55.335 188.755 55.505 189.355 ;
        RECT 56.195 189.185 57.425 189.355 ;
        RECT 55.675 188.925 56.025 189.175 ;
        RECT 54.825 188.585 55.505 188.755 ;
        RECT 54.825 187.800 55.155 188.585 ;
        RECT 55.685 187.615 56.015 188.755 ;
        RECT 56.195 188.375 56.535 189.185 ;
        RECT 56.705 188.620 57.455 188.810 ;
        RECT 56.195 187.965 56.710 188.375 ;
        RECT 56.945 187.615 57.115 188.375 ;
        RECT 57.285 187.955 57.455 188.620 ;
        RECT 57.625 188.635 57.815 189.995 ;
        RECT 57.985 189.145 58.260 189.995 ;
        RECT 58.450 189.630 58.980 189.995 ;
        RECT 59.405 189.765 59.735 190.165 ;
        RECT 58.805 189.595 58.980 189.630 ;
        RECT 57.985 188.975 58.265 189.145 ;
        RECT 57.985 188.835 58.260 188.975 ;
        RECT 58.465 188.635 58.635 189.435 ;
        RECT 57.625 188.465 58.635 188.635 ;
        RECT 58.805 189.425 59.735 189.595 ;
        RECT 59.905 189.425 60.160 189.995 ;
        RECT 58.805 188.295 58.975 189.425 ;
        RECT 59.565 189.255 59.735 189.425 ;
        RECT 57.850 188.125 58.975 188.295 ;
        RECT 59.145 188.925 59.340 189.255 ;
        RECT 59.565 188.925 59.820 189.255 ;
        RECT 59.145 187.955 59.315 188.925 ;
        RECT 59.990 188.755 60.160 189.425 ;
        RECT 57.285 187.785 59.315 187.955 ;
        RECT 59.485 187.615 59.655 188.755 ;
        RECT 59.825 187.785 60.160 188.755 ;
        RECT 60.335 189.515 60.595 189.995 ;
        RECT 60.765 189.625 61.015 190.165 ;
        RECT 60.335 188.485 60.505 189.515 ;
        RECT 61.185 189.485 61.405 189.945 ;
        RECT 61.155 189.460 61.405 189.485 ;
        RECT 60.675 188.865 60.905 189.260 ;
        RECT 61.075 189.035 61.405 189.460 ;
        RECT 61.575 189.785 62.465 189.955 ;
        RECT 61.575 189.060 61.745 189.785 ;
        RECT 61.915 189.230 62.465 189.615 ;
        RECT 62.635 189.490 62.910 189.835 ;
        RECT 63.100 189.765 63.480 190.165 ;
        RECT 63.650 189.595 63.820 189.945 ;
        RECT 63.990 189.765 64.320 190.165 ;
        RECT 64.495 189.595 64.665 189.945 ;
        RECT 64.865 189.665 65.195 190.165 ;
        RECT 61.575 188.990 62.465 189.060 ;
        RECT 61.570 188.965 62.465 188.990 ;
        RECT 61.560 188.950 62.465 188.965 ;
        RECT 61.555 188.935 62.465 188.950 ;
        RECT 61.545 188.930 62.465 188.935 ;
        RECT 61.540 188.920 62.465 188.930 ;
        RECT 61.535 188.910 62.465 188.920 ;
        RECT 61.525 188.905 62.465 188.910 ;
        RECT 61.515 188.895 62.465 188.905 ;
        RECT 61.505 188.890 62.465 188.895 ;
        RECT 61.505 188.885 61.840 188.890 ;
        RECT 61.490 188.880 61.840 188.885 ;
        RECT 61.475 188.870 61.840 188.880 ;
        RECT 61.450 188.865 61.840 188.870 ;
        RECT 60.675 188.860 61.840 188.865 ;
        RECT 60.675 188.825 61.810 188.860 ;
        RECT 60.675 188.800 61.775 188.825 ;
        RECT 60.675 188.770 61.745 188.800 ;
        RECT 60.675 188.740 61.725 188.770 ;
        RECT 60.675 188.710 61.705 188.740 ;
        RECT 60.675 188.700 61.635 188.710 ;
        RECT 60.675 188.690 61.610 188.700 ;
        RECT 60.675 188.675 61.590 188.690 ;
        RECT 60.675 188.660 61.570 188.675 ;
        RECT 60.780 188.650 61.565 188.660 ;
        RECT 60.780 188.615 61.550 188.650 ;
        RECT 60.335 187.785 60.610 188.485 ;
        RECT 60.780 188.365 61.535 188.615 ;
        RECT 61.705 188.295 62.035 188.540 ;
        RECT 62.205 188.440 62.465 188.890 ;
        RECT 62.635 188.755 62.805 189.490 ;
        RECT 63.080 189.425 64.665 189.595 ;
        RECT 63.080 189.255 63.250 189.425 ;
        RECT 65.390 189.255 65.635 189.945 ;
        RECT 65.805 189.665 66.145 190.165 ;
        RECT 66.315 189.665 66.615 189.995 ;
        RECT 66.785 189.685 67.060 190.165 ;
        RECT 62.975 188.925 63.250 189.255 ;
        RECT 63.420 188.925 63.800 189.255 ;
        RECT 63.080 188.755 63.250 188.925 ;
        RECT 61.850 188.270 62.035 188.295 ;
        RECT 61.850 188.170 62.465 188.270 ;
        RECT 60.780 187.615 61.035 188.160 ;
        RECT 61.205 187.785 61.685 188.125 ;
        RECT 61.860 187.615 62.465 188.170 ;
        RECT 62.635 187.785 62.910 188.755 ;
        RECT 63.080 188.585 63.740 188.755 ;
        RECT 63.970 188.635 64.710 189.255 ;
        RECT 64.980 188.925 65.635 189.255 ;
        RECT 65.805 188.925 66.145 189.495 ;
        RECT 63.570 188.465 63.740 188.585 ;
        RECT 64.880 188.465 65.200 188.755 ;
        RECT 63.120 187.615 63.400 188.415 ;
        RECT 63.570 188.295 65.200 188.465 ;
        RECT 65.395 188.330 65.635 188.925 ;
        RECT 66.315 188.755 66.485 189.665 ;
        RECT 67.240 189.515 67.535 189.905 ;
        RECT 67.705 189.685 67.960 190.165 ;
        RECT 68.135 189.515 68.395 189.905 ;
        RECT 68.565 189.685 68.845 190.165 ;
        RECT 66.655 188.925 67.005 189.495 ;
        RECT 67.240 189.345 68.890 189.515 ;
        RECT 67.175 189.005 68.315 189.175 ;
        RECT 67.175 188.755 67.345 189.005 ;
        RECT 68.485 188.835 68.890 189.345 ;
        RECT 69.075 189.395 70.745 190.165 ;
        RECT 71.005 189.615 71.175 189.995 ;
        RECT 71.390 189.785 71.720 190.165 ;
        RECT 71.005 189.445 71.720 189.615 ;
        RECT 69.075 188.875 69.825 189.395 ;
        RECT 63.570 187.955 65.625 188.125 ;
        RECT 63.570 187.835 65.620 187.955 ;
        RECT 65.805 187.615 66.145 188.690 ;
        RECT 66.315 188.585 67.345 188.755 ;
        RECT 68.135 188.665 68.890 188.835 ;
        RECT 69.995 188.705 70.745 189.225 ;
        RECT 70.915 188.895 71.270 189.265 ;
        RECT 71.550 189.255 71.720 189.445 ;
        RECT 71.890 189.420 72.145 189.995 ;
        RECT 71.550 188.925 71.805 189.255 ;
        RECT 71.550 188.715 71.720 188.925 ;
        RECT 66.315 187.785 66.625 188.585 ;
        RECT 68.135 188.415 68.395 188.665 ;
        RECT 66.795 187.615 67.105 188.415 ;
        RECT 67.275 188.245 68.395 188.415 ;
        RECT 67.275 187.785 67.535 188.245 ;
        RECT 67.705 187.615 67.960 188.075 ;
        RECT 68.135 187.785 68.395 188.245 ;
        RECT 68.565 187.615 68.850 188.485 ;
        RECT 69.075 187.615 70.745 188.705 ;
        RECT 71.005 188.545 71.720 188.715 ;
        RECT 71.975 188.690 72.145 189.420 ;
        RECT 72.320 189.325 72.580 190.165 ;
        RECT 73.840 189.655 74.080 190.165 ;
        RECT 74.260 189.655 74.540 189.985 ;
        RECT 74.770 189.655 74.985 190.165 ;
        RECT 73.735 188.925 74.090 189.485 ;
        RECT 71.005 187.785 71.175 188.545 ;
        RECT 71.390 187.615 71.720 188.375 ;
        RECT 71.890 187.785 72.145 188.690 ;
        RECT 72.320 187.615 72.580 188.765 ;
        RECT 74.260 188.755 74.430 189.655 ;
        RECT 74.600 188.925 74.865 189.485 ;
        RECT 75.155 189.425 75.770 189.995 ;
        RECT 76.025 189.695 76.315 190.165 ;
        RECT 76.485 189.525 76.815 189.995 ;
        RECT 76.985 189.695 77.155 190.165 ;
        RECT 77.325 189.525 77.655 189.995 ;
        RECT 76.485 189.515 77.655 189.525 ;
        RECT 75.115 188.755 75.285 189.255 ;
        RECT 73.860 188.585 75.285 188.755 ;
        RECT 73.860 188.410 74.250 188.585 ;
        RECT 74.735 187.615 75.065 188.415 ;
        RECT 75.455 188.405 75.770 189.425 ;
        RECT 76.055 189.345 77.655 189.515 ;
        RECT 77.825 189.345 78.100 190.165 ;
        RECT 78.275 189.395 79.945 190.165 ;
        RECT 80.115 189.440 80.405 190.165 ;
        RECT 76.055 188.805 76.270 189.345 ;
        RECT 76.440 188.975 77.210 189.175 ;
        RECT 77.380 188.975 78.100 189.175 ;
        RECT 78.275 188.875 79.025 189.395 ;
        RECT 76.055 188.585 76.815 188.805 ;
        RECT 75.235 187.785 75.770 188.405 ;
        RECT 76.015 187.955 76.315 188.415 ;
        RECT 76.485 188.125 76.815 188.585 ;
        RECT 76.985 188.585 78.100 188.795 ;
        RECT 79.195 188.705 79.945 189.225 ;
        RECT 80.575 189.180 80.845 189.995 ;
        RECT 81.015 189.425 81.685 190.165 ;
        RECT 81.855 189.595 82.150 189.940 ;
        RECT 82.330 189.765 82.705 190.165 ;
        RECT 82.920 189.595 83.250 189.940 ;
        RECT 81.855 189.425 83.250 189.595 ;
        RECT 83.500 189.425 84.085 189.995 ;
        RECT 84.255 189.785 85.145 189.955 ;
        RECT 76.985 187.955 77.155 188.585 ;
        RECT 76.015 187.785 77.155 187.955 ;
        RECT 77.325 187.615 77.655 188.415 ;
        RECT 77.825 187.785 78.100 188.585 ;
        RECT 78.275 187.615 79.945 188.705 ;
        RECT 80.115 187.615 80.405 188.780 ;
        RECT 80.575 187.785 80.925 189.180 ;
        RECT 81.095 188.755 81.265 189.255 ;
        RECT 81.435 188.925 81.770 189.255 ;
        RECT 81.940 188.925 82.280 189.255 ;
        RECT 81.095 188.585 81.840 188.755 ;
        RECT 81.095 187.615 81.500 188.415 ;
        RECT 81.670 187.955 81.840 188.585 ;
        RECT 82.010 188.180 82.280 188.925 ;
        RECT 82.470 188.925 82.760 189.255 ;
        RECT 82.930 188.925 83.330 189.255 ;
        RECT 82.470 188.180 82.705 188.925 ;
        RECT 83.500 188.755 83.670 189.425 ;
        RECT 83.840 188.925 84.085 189.255 ;
        RECT 84.255 189.230 84.805 189.615 ;
        RECT 84.975 189.060 85.145 189.785 ;
        RECT 84.255 188.990 85.145 189.060 ;
        RECT 85.315 189.485 85.535 189.945 ;
        RECT 85.705 189.625 85.955 190.165 ;
        RECT 86.125 189.515 86.385 189.995 ;
        RECT 85.315 189.460 85.565 189.485 ;
        RECT 85.315 189.035 85.645 189.460 ;
        RECT 84.255 188.965 85.150 188.990 ;
        RECT 84.255 188.950 85.160 188.965 ;
        RECT 84.255 188.935 85.165 188.950 ;
        RECT 84.255 188.930 85.175 188.935 ;
        RECT 84.255 188.920 85.180 188.930 ;
        RECT 84.255 188.910 85.185 188.920 ;
        RECT 84.255 188.905 85.195 188.910 ;
        RECT 84.255 188.895 85.205 188.905 ;
        RECT 84.255 188.890 85.215 188.895 ;
        RECT 82.875 188.585 84.085 188.755 ;
        RECT 82.875 187.955 83.205 188.585 ;
        RECT 81.670 187.785 83.205 187.955 ;
        RECT 83.390 187.615 83.625 188.415 ;
        RECT 83.795 187.785 84.085 188.585 ;
        RECT 84.255 188.440 84.515 188.890 ;
        RECT 84.880 188.885 85.215 188.890 ;
        RECT 84.880 188.880 85.230 188.885 ;
        RECT 84.880 188.870 85.245 188.880 ;
        RECT 84.880 188.865 85.270 188.870 ;
        RECT 85.815 188.865 86.045 189.260 ;
        RECT 84.880 188.860 86.045 188.865 ;
        RECT 84.910 188.825 86.045 188.860 ;
        RECT 84.945 188.800 86.045 188.825 ;
        RECT 84.975 188.770 86.045 188.800 ;
        RECT 84.995 188.740 86.045 188.770 ;
        RECT 85.015 188.710 86.045 188.740 ;
        RECT 85.085 188.700 86.045 188.710 ;
        RECT 85.110 188.690 86.045 188.700 ;
        RECT 85.130 188.675 86.045 188.690 ;
        RECT 85.150 188.660 86.045 188.675 ;
        RECT 85.155 188.650 85.940 188.660 ;
        RECT 85.170 188.615 85.940 188.650 ;
        RECT 84.685 188.295 85.015 188.540 ;
        RECT 85.185 188.365 85.940 188.615 ;
        RECT 86.215 188.485 86.385 189.515 ;
        RECT 86.555 189.395 90.065 190.165 ;
        RECT 90.695 189.440 91.035 190.165 ;
        RECT 86.555 188.875 88.205 189.395 ;
        RECT 91.205 189.255 91.410 189.855 ;
        RECT 91.640 189.650 92.590 189.835 ;
        RECT 88.375 188.705 90.065 189.225 ;
        RECT 84.685 188.270 84.870 188.295 ;
        RECT 84.255 188.170 84.870 188.270 ;
        RECT 84.255 187.615 84.860 188.170 ;
        RECT 85.035 187.785 85.515 188.125 ;
        RECT 85.685 187.615 85.940 188.160 ;
        RECT 86.110 187.785 86.385 188.485 ;
        RECT 86.555 187.615 90.065 188.705 ;
        RECT 90.720 188.625 90.975 189.255 ;
        RECT 91.205 188.625 91.585 189.255 ;
        RECT 91.845 188.925 92.065 189.650 ;
        RECT 92.760 189.515 93.175 189.950 ;
        RECT 93.365 189.685 93.695 190.165 ;
        RECT 93.865 189.690 94.205 189.950 ;
        RECT 92.760 189.440 93.775 189.515 ;
        RECT 92.955 189.345 93.775 189.440 ;
        RECT 92.375 189.145 92.755 189.255 ;
        RECT 92.375 188.975 92.765 189.145 ;
        RECT 92.375 188.925 92.755 188.975 ;
        RECT 92.455 188.630 92.755 188.925 ;
        RECT 92.955 188.615 93.285 189.175 ;
        RECT 90.785 188.285 92.755 188.455 ;
        RECT 93.605 188.425 93.775 189.345 ;
        RECT 90.785 187.785 90.955 188.285 ;
        RECT 91.195 187.615 91.445 188.075 ;
        RECT 91.745 187.785 91.915 188.285 ;
        RECT 92.125 187.615 92.375 188.075 ;
        RECT 92.585 187.785 92.755 188.285 ;
        RECT 92.925 188.255 93.775 188.425 ;
        RECT 92.925 187.825 93.255 188.255 ;
        RECT 93.945 188.085 94.205 189.690 ;
        RECT 94.385 189.655 94.835 190.165 ;
        RECT 95.110 189.745 96.415 189.995 ;
        RECT 96.595 189.765 96.925 190.165 ;
        RECT 96.235 189.595 96.415 189.745 ;
        RECT 94.415 188.975 94.865 189.485 ;
        RECT 95.280 189.175 95.530 189.575 ;
        RECT 95.055 188.975 95.530 189.175 ;
        RECT 95.780 189.175 95.990 189.575 ;
        RECT 96.235 189.425 96.965 189.595 ;
        RECT 95.780 188.975 96.130 189.175 ;
        RECT 96.300 188.925 96.625 189.255 ;
        RECT 93.445 187.615 93.695 188.075 ;
        RECT 93.865 187.825 94.205 188.085 ;
        RECT 94.385 188.755 96.130 188.805 ;
        RECT 96.795 188.755 96.965 189.425 ;
        RECT 97.135 189.365 97.830 189.995 ;
        RECT 98.035 189.365 98.345 190.165 ;
        RECT 98.515 189.395 102.025 190.165 ;
        RECT 103.225 189.785 104.395 189.995 ;
        RECT 103.225 189.765 103.555 189.785 ;
        RECT 97.155 188.925 97.490 189.175 ;
        RECT 97.660 188.765 97.830 189.365 ;
        RECT 98.000 188.925 98.335 189.195 ;
        RECT 98.515 188.875 100.165 189.395 ;
        RECT 103.115 189.345 103.975 189.595 ;
        RECT 104.145 189.535 104.395 189.785 ;
        RECT 104.565 189.705 104.735 190.165 ;
        RECT 104.905 189.535 105.245 189.995 ;
        RECT 104.145 189.365 105.245 189.535 ;
        RECT 105.875 189.440 106.165 190.165 ;
        RECT 106.335 189.395 109.845 190.165 ;
        RECT 110.955 189.595 111.210 189.945 ;
        RECT 111.380 189.765 111.710 190.165 ;
        RECT 111.880 189.595 112.050 189.945 ;
        RECT 112.220 189.765 112.600 190.165 ;
        RECT 110.955 189.425 112.620 189.595 ;
        RECT 112.790 189.490 113.065 189.835 ;
        RECT 94.385 188.625 96.965 188.755 ;
        RECT 94.385 187.955 94.715 188.625 ;
        RECT 95.905 188.585 96.965 188.625 ;
        RECT 94.885 188.415 95.765 188.455 ;
        RECT 94.885 188.215 96.415 188.415 ;
        RECT 94.885 188.165 95.500 188.215 ;
        RECT 94.885 188.125 95.115 188.165 ;
        RECT 96.245 188.085 96.415 188.215 ;
        RECT 95.225 187.955 95.555 187.995 ;
        RECT 94.385 187.785 95.555 187.955 ;
        RECT 95.725 187.615 96.100 187.995 ;
        RECT 96.650 187.615 96.915 188.395 ;
        RECT 97.135 187.615 97.395 188.755 ;
        RECT 97.565 187.785 97.895 188.765 ;
        RECT 98.065 187.615 98.345 188.755 ;
        RECT 100.335 188.705 102.025 189.225 ;
        RECT 98.515 187.615 102.025 188.705 ;
        RECT 103.115 188.755 103.395 189.345 ;
        RECT 103.565 188.925 104.315 189.175 ;
        RECT 104.485 188.925 105.245 189.175 ;
        RECT 106.335 188.875 107.985 189.395 ;
        RECT 112.450 189.255 112.620 189.425 ;
        RECT 103.115 188.585 104.815 188.755 ;
        RECT 103.220 187.615 103.475 188.415 ;
        RECT 103.645 187.785 103.975 188.585 ;
        RECT 104.145 187.615 104.315 188.415 ;
        RECT 104.485 187.785 104.815 188.585 ;
        RECT 104.985 187.615 105.245 188.755 ;
        RECT 105.875 187.615 106.165 188.780 ;
        RECT 108.155 188.705 109.845 189.225 ;
        RECT 110.935 188.925 111.285 189.255 ;
        RECT 111.455 188.925 112.280 189.255 ;
        RECT 112.450 188.925 112.725 189.255 ;
        RECT 106.335 187.615 109.845 188.705 ;
        RECT 110.955 188.465 111.285 188.755 ;
        RECT 111.455 188.635 111.680 188.925 ;
        RECT 112.450 188.755 112.620 188.925 ;
        RECT 112.895 188.755 113.065 189.490 ;
        RECT 113.235 189.335 113.525 190.165 ;
        RECT 113.715 189.355 113.955 190.165 ;
        RECT 114.125 189.355 114.455 189.995 ;
        RECT 114.625 189.355 114.895 190.165 ;
        RECT 115.075 189.395 118.585 190.165 ;
        RECT 119.305 189.515 119.475 189.995 ;
        RECT 119.645 189.685 119.975 190.165 ;
        RECT 120.200 189.745 121.735 189.995 ;
        RECT 120.200 189.515 120.370 189.745 ;
        RECT 113.695 188.925 114.045 189.175 ;
        RECT 111.950 188.585 112.620 188.755 ;
        RECT 111.950 188.465 112.120 188.585 ;
        RECT 110.955 188.295 112.120 188.465 ;
        RECT 110.935 187.835 112.130 188.125 ;
        RECT 112.300 187.615 112.580 188.415 ;
        RECT 112.790 187.785 113.065 188.755 ;
        RECT 113.235 187.615 113.525 188.820 ;
        RECT 114.215 188.755 114.385 189.355 ;
        RECT 114.555 188.925 114.905 189.175 ;
        RECT 115.075 188.875 116.725 189.395 ;
        RECT 119.305 189.345 120.370 189.515 ;
        RECT 113.705 188.585 114.385 188.755 ;
        RECT 113.705 187.800 114.035 188.585 ;
        RECT 114.565 187.615 114.895 188.755 ;
        RECT 116.895 188.705 118.585 189.225 ;
        RECT 120.550 189.175 120.830 189.575 ;
        RECT 119.220 188.965 119.570 189.175 ;
        RECT 119.740 188.975 120.185 189.175 ;
        RECT 120.355 188.975 120.830 189.175 ;
        RECT 121.100 189.175 121.385 189.575 ;
        RECT 121.565 189.515 121.735 189.745 ;
        RECT 121.905 189.685 122.235 190.165 ;
        RECT 122.450 189.665 122.705 189.995 ;
        RECT 122.495 189.655 122.705 189.665 ;
        RECT 122.520 189.585 122.705 189.655 ;
        RECT 121.565 189.345 122.365 189.515 ;
        RECT 121.100 188.975 121.430 189.175 ;
        RECT 121.600 189.145 121.965 189.175 ;
        RECT 121.600 188.975 121.975 189.145 ;
        RECT 122.195 188.795 122.365 189.345 ;
        RECT 115.075 187.615 118.585 188.705 ;
        RECT 119.305 188.625 122.365 188.795 ;
        RECT 119.305 187.785 119.475 188.625 ;
        RECT 122.535 188.455 122.705 189.585 ;
        RECT 122.895 189.415 124.105 190.165 ;
        RECT 124.335 189.685 124.615 190.165 ;
        RECT 124.785 189.515 125.045 189.905 ;
        RECT 125.220 189.685 125.475 190.165 ;
        RECT 125.645 189.515 125.940 189.905 ;
        RECT 126.120 189.685 126.395 190.165 ;
        RECT 126.565 189.665 126.865 189.995 ;
        RECT 122.895 188.875 123.415 189.415 ;
        RECT 124.290 189.345 125.940 189.515 ;
        RECT 123.585 188.705 124.105 189.245 ;
        RECT 119.645 187.955 119.975 188.455 ;
        RECT 120.145 188.215 121.780 188.455 ;
        RECT 120.145 188.125 120.375 188.215 ;
        RECT 120.485 187.955 120.815 187.995 ;
        RECT 119.645 187.785 120.815 187.955 ;
        RECT 121.005 187.615 121.360 188.035 ;
        RECT 121.530 187.785 121.780 188.215 ;
        RECT 121.950 187.615 122.280 188.375 ;
        RECT 122.450 187.785 122.705 188.455 ;
        RECT 122.895 187.615 124.105 188.705 ;
        RECT 124.290 188.835 124.695 189.345 ;
        RECT 124.865 189.005 126.005 189.175 ;
        RECT 124.290 188.665 125.045 188.835 ;
        RECT 124.330 187.615 124.615 188.485 ;
        RECT 124.785 188.415 125.045 188.665 ;
        RECT 125.835 188.755 126.005 189.005 ;
        RECT 126.175 188.925 126.525 189.495 ;
        RECT 126.695 188.755 126.865 189.665 ;
        RECT 127.040 189.635 127.330 189.985 ;
        RECT 127.525 189.805 127.855 190.165 ;
        RECT 128.025 189.635 128.255 189.940 ;
        RECT 127.040 189.465 128.255 189.635 ;
        RECT 128.445 189.485 128.615 189.860 ;
        RECT 128.445 189.315 128.645 189.485 ;
        RECT 128.895 189.435 129.185 190.165 ;
        RECT 128.445 189.295 128.615 189.315 ;
        RECT 127.100 188.925 127.360 189.255 ;
        RECT 127.540 188.925 127.925 189.255 ;
        RECT 128.095 189.125 128.615 189.295 ;
        RECT 125.835 188.585 126.865 188.755 ;
        RECT 124.785 188.245 125.905 188.415 ;
        RECT 124.785 187.785 125.045 188.245 ;
        RECT 125.220 187.615 125.475 188.075 ;
        RECT 125.645 187.785 125.905 188.245 ;
        RECT 126.075 187.615 126.385 188.415 ;
        RECT 126.555 187.785 126.865 188.585 ;
        RECT 127.040 187.615 127.360 188.755 ;
        RECT 127.540 187.875 127.735 188.925 ;
        RECT 128.095 188.745 128.265 189.125 ;
        RECT 127.915 188.465 128.265 188.745 ;
        RECT 128.455 188.595 128.700 188.955 ;
        RECT 128.885 188.925 129.185 189.255 ;
        RECT 129.365 189.235 129.595 189.875 ;
        RECT 129.775 189.615 130.085 189.985 ;
        RECT 130.265 189.795 130.935 190.165 ;
        RECT 129.775 189.415 131.005 189.615 ;
        RECT 129.365 188.925 129.890 189.235 ;
        RECT 130.070 188.925 130.535 189.235 ;
        RECT 130.715 188.745 131.005 189.415 ;
        RECT 128.895 188.505 130.055 188.745 ;
        RECT 127.915 187.785 128.245 188.465 ;
        RECT 128.445 187.615 128.700 188.415 ;
        RECT 128.895 187.795 129.155 188.505 ;
        RECT 129.325 187.615 129.655 188.325 ;
        RECT 129.825 187.795 130.055 188.505 ;
        RECT 130.235 188.525 131.005 188.745 ;
        RECT 130.235 187.795 130.505 188.525 ;
        RECT 130.685 187.615 131.025 188.345 ;
        RECT 131.195 187.795 131.455 189.985 ;
        RECT 131.635 189.440 131.925 190.165 ;
        RECT 133.175 189.605 133.505 189.995 ;
        RECT 133.675 189.775 134.860 189.945 ;
        RECT 135.120 189.695 135.290 190.165 ;
        RECT 133.175 189.425 133.685 189.605 ;
        RECT 133.015 188.965 133.345 189.255 ;
        RECT 133.515 188.795 133.685 189.425 ;
        RECT 134.090 189.515 134.475 189.605 ;
        RECT 135.460 189.515 135.790 189.980 ;
        RECT 134.090 189.345 135.790 189.515 ;
        RECT 135.960 189.345 136.130 190.165 ;
        RECT 136.300 189.345 136.985 189.985 ;
        RECT 137.160 189.400 137.615 190.165 ;
        RECT 137.890 189.785 139.190 189.995 ;
        RECT 139.445 189.805 139.775 190.165 ;
        RECT 139.020 189.635 139.190 189.785 ;
        RECT 139.945 189.665 140.205 189.995 ;
        RECT 139.975 189.655 140.205 189.665 ;
        RECT 133.855 188.965 134.185 189.175 ;
        RECT 134.365 188.925 134.745 189.175 ;
        RECT 131.635 187.615 131.925 188.780 ;
        RECT 133.170 188.625 134.255 188.795 ;
        RECT 133.170 187.785 133.470 188.625 ;
        RECT 133.665 187.615 133.915 188.455 ;
        RECT 134.085 188.375 134.255 188.625 ;
        RECT 134.425 188.545 134.745 188.925 ;
        RECT 134.935 188.965 135.420 189.175 ;
        RECT 135.610 188.965 136.060 189.175 ;
        RECT 136.230 188.965 136.565 189.175 ;
        RECT 134.935 188.805 135.310 188.965 ;
        RECT 134.915 188.635 135.310 188.805 ;
        RECT 136.230 188.795 136.400 188.965 ;
        RECT 134.935 188.545 135.310 188.635 ;
        RECT 135.480 188.625 136.400 188.795 ;
        RECT 135.480 188.375 135.650 188.625 ;
        RECT 134.085 188.205 135.650 188.375 ;
        RECT 134.505 187.785 135.310 188.205 ;
        RECT 135.820 187.615 136.150 188.455 ;
        RECT 136.735 188.375 136.985 189.345 ;
        RECT 138.090 189.175 138.310 189.575 ;
        RECT 137.155 188.975 137.645 189.175 ;
        RECT 137.835 188.965 138.310 189.175 ;
        RECT 138.555 189.175 138.765 189.575 ;
        RECT 139.020 189.510 139.775 189.635 ;
        RECT 139.020 189.465 139.865 189.510 ;
        RECT 139.595 189.345 139.865 189.465 ;
        RECT 138.555 188.965 138.885 189.175 ;
        RECT 139.055 188.905 139.465 189.210 ;
        RECT 136.320 187.785 136.985 188.375 ;
        RECT 137.160 188.735 138.335 188.795 ;
        RECT 139.695 188.770 139.865 189.345 ;
        RECT 139.665 188.735 139.865 188.770 ;
        RECT 137.160 188.625 139.865 188.735 ;
        RECT 137.160 188.005 137.415 188.625 ;
        RECT 138.005 188.565 139.805 188.625 ;
        RECT 138.005 188.535 138.335 188.565 ;
        RECT 140.035 188.465 140.205 189.655 ;
        RECT 140.395 189.435 140.685 190.165 ;
        RECT 140.385 188.925 140.685 189.255 ;
        RECT 140.865 189.235 141.095 189.875 ;
        RECT 141.275 189.615 141.585 189.985 ;
        RECT 141.765 189.795 142.435 190.165 ;
        RECT 141.275 189.415 142.505 189.615 ;
        RECT 140.865 188.925 141.390 189.235 ;
        RECT 141.570 188.925 142.035 189.235 ;
        RECT 142.215 188.745 142.505 189.415 ;
        RECT 137.665 188.365 137.850 188.455 ;
        RECT 138.440 188.365 139.275 188.375 ;
        RECT 137.665 188.165 139.275 188.365 ;
        RECT 137.665 188.125 137.895 188.165 ;
        RECT 137.160 187.785 137.495 188.005 ;
        RECT 138.500 187.615 138.855 187.995 ;
        RECT 139.025 187.785 139.275 188.165 ;
        RECT 139.525 187.615 139.775 188.395 ;
        RECT 139.945 187.785 140.205 188.465 ;
        RECT 140.395 188.505 141.555 188.745 ;
        RECT 140.395 187.795 140.655 188.505 ;
        RECT 140.825 187.615 141.155 188.325 ;
        RECT 141.325 187.795 141.555 188.505 ;
        RECT 141.735 188.525 142.505 188.745 ;
        RECT 141.735 187.795 142.005 188.525 ;
        RECT 142.185 187.615 142.525 188.345 ;
        RECT 142.695 187.795 142.955 189.985 ;
        RECT 143.135 189.395 144.805 190.165 ;
        RECT 143.135 188.875 143.885 189.395 ;
        RECT 144.975 189.365 145.315 189.995 ;
        RECT 145.485 189.365 145.735 190.165 ;
        RECT 145.925 189.515 146.255 189.995 ;
        RECT 146.425 189.705 146.650 190.165 ;
        RECT 146.820 189.515 147.150 189.995 ;
        RECT 144.055 188.705 144.805 189.225 ;
        RECT 143.135 187.615 144.805 188.705 ;
        RECT 144.975 188.805 145.150 189.365 ;
        RECT 145.925 189.345 147.150 189.515 ;
        RECT 147.780 189.385 148.280 189.995 ;
        RECT 149.585 189.440 149.915 189.950 ;
        RECT 150.085 189.765 150.415 190.165 ;
        RECT 151.465 189.595 151.795 189.935 ;
        RECT 151.965 189.765 152.295 190.165 ;
        RECT 145.320 189.005 146.015 189.175 ;
        RECT 144.975 188.755 145.205 188.805 ;
        RECT 145.845 188.755 146.015 189.005 ;
        RECT 146.190 188.975 146.610 189.175 ;
        RECT 146.780 188.975 147.110 189.175 ;
        RECT 147.280 188.975 147.610 189.175 ;
        RECT 147.780 188.755 147.950 189.385 ;
        RECT 148.135 188.925 148.485 189.175 ;
        RECT 144.975 187.785 145.315 188.755 ;
        RECT 145.485 187.615 145.655 188.755 ;
        RECT 145.845 188.585 148.280 188.755 ;
        RECT 145.925 187.615 146.175 188.415 ;
        RECT 146.820 187.785 147.150 188.585 ;
        RECT 147.450 187.615 147.780 188.415 ;
        RECT 147.950 187.785 148.280 188.585 ;
        RECT 149.585 188.675 149.775 189.440 ;
        RECT 150.085 189.425 152.450 189.595 ;
        RECT 150.085 189.255 150.255 189.425 ;
        RECT 149.945 188.925 150.255 189.255 ;
        RECT 150.425 188.925 150.730 189.255 ;
        RECT 149.585 187.825 149.915 188.675 ;
        RECT 150.085 187.615 150.335 188.755 ;
        RECT 150.515 188.595 150.730 188.925 ;
        RECT 150.905 188.595 151.190 189.255 ;
        RECT 151.385 188.595 151.650 189.255 ;
        RECT 151.865 188.595 152.110 189.255 ;
        RECT 152.280 188.425 152.450 189.425 ;
        RECT 152.795 189.395 156.305 190.165 ;
        RECT 156.935 189.415 158.145 190.165 ;
        RECT 152.795 188.875 154.445 189.395 ;
        RECT 154.615 188.705 156.305 189.225 ;
        RECT 150.525 188.255 151.815 188.425 ;
        RECT 150.525 187.835 150.775 188.255 ;
        RECT 151.005 187.615 151.335 188.085 ;
        RECT 151.565 187.835 151.815 188.255 ;
        RECT 151.995 188.255 152.450 188.425 ;
        RECT 151.995 187.825 152.325 188.255 ;
        RECT 152.795 187.615 156.305 188.705 ;
        RECT 156.935 188.705 157.455 189.245 ;
        RECT 157.625 188.875 158.145 189.415 ;
        RECT 156.935 187.615 158.145 188.705 ;
        RECT 2.750 187.445 158.230 187.615 ;
        RECT 2.835 186.355 4.045 187.445 ;
        RECT 4.305 186.775 4.475 187.275 ;
        RECT 4.645 186.945 4.975 187.445 ;
        RECT 4.305 186.605 4.970 186.775 ;
        RECT 2.835 185.645 3.355 186.185 ;
        RECT 3.525 185.815 4.045 186.355 ;
        RECT 4.220 185.785 4.570 186.435 ;
        RECT 2.835 184.895 4.045 185.645 ;
        RECT 4.740 185.615 4.970 186.605 ;
        RECT 4.305 185.445 4.970 185.615 ;
        RECT 4.305 185.155 4.475 185.445 ;
        RECT 4.645 184.895 4.975 185.275 ;
        RECT 5.145 185.155 5.370 187.275 ;
        RECT 5.585 186.945 5.915 187.445 ;
        RECT 6.085 186.775 6.255 187.275 ;
        RECT 6.490 187.060 7.320 187.230 ;
        RECT 7.560 187.065 7.940 187.445 ;
        RECT 5.560 186.605 6.255 186.775 ;
        RECT 5.560 185.635 5.730 186.605 ;
        RECT 5.900 185.815 6.310 186.435 ;
        RECT 6.480 186.385 6.980 186.765 ;
        RECT 5.560 185.445 6.255 185.635 ;
        RECT 6.480 185.515 6.700 186.385 ;
        RECT 7.150 186.215 7.320 187.060 ;
        RECT 8.120 186.895 8.290 187.185 ;
        RECT 8.460 187.065 8.790 187.445 ;
        RECT 9.260 186.975 9.890 187.225 ;
        RECT 10.070 187.065 10.490 187.445 ;
        RECT 9.720 186.895 9.890 186.975 ;
        RECT 10.690 186.895 10.930 187.185 ;
        RECT 7.490 186.645 8.860 186.895 ;
        RECT 7.490 186.385 7.740 186.645 ;
        RECT 8.250 186.215 8.500 186.375 ;
        RECT 7.150 186.045 8.500 186.215 ;
        RECT 7.150 186.005 7.570 186.045 ;
        RECT 6.880 185.455 7.230 185.825 ;
        RECT 5.585 184.895 5.915 185.275 ;
        RECT 6.085 185.115 6.255 185.445 ;
        RECT 7.400 185.275 7.570 186.005 ;
        RECT 8.670 185.875 8.860 186.645 ;
        RECT 7.740 185.545 8.150 185.875 ;
        RECT 8.440 185.535 8.860 185.875 ;
        RECT 9.030 186.465 9.550 186.775 ;
        RECT 9.720 186.725 10.930 186.895 ;
        RECT 11.160 186.755 11.490 187.445 ;
        RECT 9.030 185.705 9.200 186.465 ;
        RECT 9.370 185.875 9.550 186.285 ;
        RECT 9.720 186.215 9.890 186.725 ;
        RECT 11.660 186.575 11.830 187.185 ;
        RECT 12.100 186.725 12.430 187.235 ;
        RECT 11.660 186.555 11.980 186.575 ;
        RECT 10.060 186.385 11.980 186.555 ;
        RECT 9.720 186.045 11.620 186.215 ;
        RECT 9.950 185.705 10.280 185.825 ;
        RECT 9.030 185.535 10.280 185.705 ;
        RECT 6.555 185.075 7.570 185.275 ;
        RECT 7.740 184.895 8.150 185.335 ;
        RECT 8.440 185.105 8.690 185.535 ;
        RECT 8.890 184.895 9.210 185.355 ;
        RECT 10.450 185.285 10.620 186.045 ;
        RECT 11.290 185.985 11.620 186.045 ;
        RECT 10.810 185.815 11.140 185.875 ;
        RECT 10.810 185.545 11.470 185.815 ;
        RECT 11.790 185.490 11.980 186.385 ;
        RECT 9.770 185.115 10.620 185.285 ;
        RECT 10.820 184.895 11.480 185.375 ;
        RECT 11.660 185.160 11.980 185.490 ;
        RECT 12.180 186.135 12.430 186.725 ;
        RECT 12.610 186.645 12.895 187.445 ;
        RECT 13.075 186.465 13.330 187.135 ;
        RECT 12.180 185.805 12.980 186.135 ;
        RECT 12.180 185.155 12.430 185.805 ;
        RECT 13.150 185.605 13.330 186.465 ;
        RECT 13.875 186.355 15.545 187.445 ;
        RECT 13.075 185.405 13.330 185.605 ;
        RECT 13.875 185.665 14.625 186.185 ;
        RECT 14.795 185.835 15.545 186.355 ;
        RECT 15.715 186.280 16.005 187.445 ;
        RECT 16.635 186.370 16.905 187.275 ;
        RECT 17.075 186.685 17.405 187.445 ;
        RECT 17.585 186.515 17.755 187.275 ;
        RECT 12.610 184.895 12.895 185.355 ;
        RECT 13.075 185.235 13.415 185.405 ;
        RECT 13.075 185.075 13.330 185.235 ;
        RECT 13.875 184.895 15.545 185.665 ;
        RECT 15.715 184.895 16.005 185.620 ;
        RECT 16.635 185.570 16.805 186.370 ;
        RECT 17.090 186.345 17.755 186.515 ;
        RECT 17.090 186.200 17.260 186.345 ;
        RECT 16.975 185.870 17.260 186.200 ;
        RECT 18.480 186.305 18.815 187.275 ;
        RECT 18.985 186.305 19.155 187.445 ;
        RECT 19.325 187.105 21.355 187.275 ;
        RECT 17.090 185.615 17.260 185.870 ;
        RECT 17.495 185.795 17.825 186.165 ;
        RECT 18.480 185.635 18.650 186.305 ;
        RECT 19.325 186.135 19.495 187.105 ;
        RECT 18.820 185.805 19.075 186.135 ;
        RECT 19.300 185.805 19.495 186.135 ;
        RECT 19.665 186.765 20.790 186.935 ;
        RECT 18.905 185.635 19.075 185.805 ;
        RECT 19.665 185.635 19.835 186.765 ;
        RECT 16.635 185.065 16.895 185.570 ;
        RECT 17.090 185.445 17.755 185.615 ;
        RECT 17.075 184.895 17.405 185.275 ;
        RECT 17.585 185.065 17.755 185.445 ;
        RECT 18.480 185.065 18.735 185.635 ;
        RECT 18.905 185.465 19.835 185.635 ;
        RECT 20.005 186.425 21.015 186.595 ;
        RECT 20.005 185.625 20.175 186.425 ;
        RECT 19.660 185.430 19.835 185.465 ;
        RECT 18.905 184.895 19.235 185.295 ;
        RECT 19.660 185.065 20.190 185.430 ;
        RECT 20.380 185.405 20.655 186.225 ;
        RECT 20.375 185.235 20.655 185.405 ;
        RECT 20.380 185.065 20.655 185.235 ;
        RECT 20.825 185.065 21.015 186.425 ;
        RECT 21.185 186.440 21.355 187.105 ;
        RECT 21.525 186.685 21.695 187.445 ;
        RECT 21.930 186.685 22.445 187.095 ;
        RECT 21.185 186.250 21.935 186.440 ;
        RECT 22.105 185.875 22.445 186.685 ;
        RECT 22.620 186.775 22.875 187.275 ;
        RECT 23.045 186.945 23.375 187.445 ;
        RECT 22.620 186.605 23.370 186.775 ;
        RECT 21.215 185.705 22.445 185.875 ;
        RECT 22.620 185.785 22.970 186.435 ;
        RECT 21.195 184.895 21.705 185.430 ;
        RECT 21.925 185.100 22.170 185.705 ;
        RECT 23.140 185.615 23.370 186.605 ;
        RECT 22.620 185.445 23.370 185.615 ;
        RECT 22.620 185.155 22.875 185.445 ;
        RECT 23.045 184.895 23.375 185.275 ;
        RECT 23.545 185.155 23.715 187.275 ;
        RECT 23.885 186.475 24.210 187.260 ;
        RECT 24.380 186.985 24.630 187.445 ;
        RECT 24.800 186.945 25.050 187.275 ;
        RECT 25.265 186.945 25.945 187.275 ;
        RECT 24.800 186.815 24.970 186.945 ;
        RECT 24.575 186.645 24.970 186.815 ;
        RECT 23.945 185.425 24.405 186.475 ;
        RECT 24.575 185.285 24.745 186.645 ;
        RECT 25.140 186.385 25.605 186.775 ;
        RECT 24.915 185.575 25.265 186.195 ;
        RECT 25.435 185.795 25.605 186.385 ;
        RECT 25.775 186.165 25.945 186.945 ;
        RECT 26.115 186.845 26.285 187.185 ;
        RECT 26.520 187.015 26.850 187.445 ;
        RECT 27.020 186.845 27.190 187.185 ;
        RECT 27.485 186.985 27.855 187.445 ;
        RECT 26.115 186.675 27.190 186.845 ;
        RECT 28.025 186.815 28.195 187.275 ;
        RECT 28.430 186.935 29.300 187.275 ;
        RECT 29.470 186.985 29.720 187.445 ;
        RECT 27.635 186.645 28.195 186.815 ;
        RECT 27.635 186.505 27.805 186.645 ;
        RECT 26.305 186.335 27.805 186.505 ;
        RECT 28.500 186.475 28.960 186.765 ;
        RECT 25.775 185.995 27.465 186.165 ;
        RECT 25.435 185.575 25.790 185.795 ;
        RECT 25.960 185.285 26.130 185.995 ;
        RECT 26.335 185.575 27.125 185.825 ;
        RECT 27.295 185.815 27.465 185.995 ;
        RECT 27.635 185.645 27.805 186.335 ;
        RECT 24.075 184.895 24.405 185.255 ;
        RECT 24.575 185.115 25.070 185.285 ;
        RECT 25.275 185.115 26.130 185.285 ;
        RECT 27.005 184.895 27.335 185.355 ;
        RECT 27.545 185.255 27.805 185.645 ;
        RECT 27.995 186.465 28.960 186.475 ;
        RECT 29.130 186.555 29.300 186.935 ;
        RECT 29.890 186.895 30.060 187.185 ;
        RECT 30.240 187.065 30.570 187.445 ;
        RECT 29.890 186.725 30.690 186.895 ;
        RECT 27.995 186.305 28.670 186.465 ;
        RECT 29.130 186.385 30.350 186.555 ;
        RECT 27.995 185.515 28.205 186.305 ;
        RECT 29.130 186.295 29.300 186.385 ;
        RECT 28.375 185.515 28.725 186.135 ;
        RECT 28.895 186.125 29.300 186.295 ;
        RECT 28.895 185.345 29.065 186.125 ;
        RECT 29.235 185.675 29.455 185.955 ;
        RECT 29.635 185.845 30.175 186.215 ;
        RECT 30.520 186.135 30.690 186.725 ;
        RECT 30.910 186.305 31.215 187.445 ;
        RECT 31.385 186.255 31.640 187.135 ;
        RECT 31.905 186.700 32.175 187.445 ;
        RECT 32.805 187.440 39.080 187.445 ;
        RECT 32.345 186.530 32.635 187.270 ;
        RECT 32.805 186.715 33.060 187.440 ;
        RECT 33.245 186.545 33.505 187.270 ;
        RECT 33.675 186.715 33.920 187.440 ;
        RECT 34.105 186.545 34.365 187.270 ;
        RECT 34.535 186.715 34.780 187.440 ;
        RECT 34.965 186.545 35.225 187.270 ;
        RECT 35.395 186.715 35.640 187.440 ;
        RECT 35.810 186.545 36.070 187.270 ;
        RECT 36.240 186.715 36.500 187.440 ;
        RECT 36.670 186.545 36.930 187.270 ;
        RECT 37.100 186.715 37.360 187.440 ;
        RECT 37.530 186.545 37.790 187.270 ;
        RECT 37.960 186.715 38.220 187.440 ;
        RECT 38.390 186.545 38.650 187.270 ;
        RECT 38.820 186.645 39.080 187.440 ;
        RECT 33.245 186.530 38.650 186.545 ;
        RECT 30.520 186.105 31.260 186.135 ;
        RECT 29.235 185.505 29.765 185.675 ;
        RECT 27.545 185.085 27.895 185.255 ;
        RECT 28.115 185.065 29.065 185.345 ;
        RECT 29.235 184.895 29.425 185.335 ;
        RECT 29.595 185.275 29.765 185.505 ;
        RECT 29.935 185.445 30.175 185.845 ;
        RECT 30.345 185.805 31.260 186.105 ;
        RECT 30.345 185.630 30.670 185.805 ;
        RECT 30.345 185.275 30.665 185.630 ;
        RECT 31.430 185.605 31.640 186.255 ;
        RECT 29.595 185.105 30.665 185.275 ;
        RECT 30.910 184.895 31.215 185.355 ;
        RECT 31.385 185.075 31.640 185.605 ;
        RECT 31.905 186.305 38.650 186.530 ;
        RECT 31.905 185.715 33.070 186.305 ;
        RECT 39.250 186.135 39.500 187.270 ;
        RECT 39.680 186.635 39.940 187.445 ;
        RECT 40.115 186.135 40.360 187.275 ;
        RECT 40.540 186.635 40.835 187.445 ;
        RECT 41.475 186.280 41.765 187.445 ;
        RECT 41.940 186.305 42.275 187.275 ;
        RECT 42.445 186.305 42.615 187.445 ;
        RECT 42.785 187.105 44.815 187.275 ;
        RECT 33.240 185.885 40.360 186.135 ;
        RECT 31.905 185.545 38.650 185.715 ;
        RECT 31.905 184.895 32.205 185.375 ;
        RECT 32.375 185.090 32.635 185.545 ;
        RECT 32.805 184.895 33.065 185.375 ;
        RECT 33.245 185.090 33.505 185.545 ;
        RECT 33.675 184.895 33.925 185.375 ;
        RECT 34.105 185.090 34.365 185.545 ;
        RECT 34.535 184.895 34.785 185.375 ;
        RECT 34.965 185.090 35.225 185.545 ;
        RECT 35.395 184.895 35.640 185.375 ;
        RECT 35.810 185.090 36.085 185.545 ;
        RECT 36.255 184.895 36.500 185.375 ;
        RECT 36.670 185.090 36.930 185.545 ;
        RECT 37.100 184.895 37.360 185.375 ;
        RECT 37.530 185.090 37.790 185.545 ;
        RECT 37.960 184.895 38.220 185.375 ;
        RECT 38.390 185.090 38.650 185.545 ;
        RECT 38.820 184.895 39.080 185.455 ;
        RECT 39.250 185.075 39.500 185.885 ;
        RECT 39.680 184.895 39.940 185.420 ;
        RECT 40.110 185.075 40.360 185.885 ;
        RECT 40.530 185.575 40.845 186.135 ;
        RECT 41.940 185.635 42.110 186.305 ;
        RECT 42.785 186.135 42.955 187.105 ;
        RECT 42.280 185.805 42.535 186.135 ;
        RECT 42.760 185.805 42.955 186.135 ;
        RECT 43.125 186.765 44.250 186.935 ;
        RECT 42.365 185.635 42.535 185.805 ;
        RECT 43.125 185.635 43.295 186.765 ;
        RECT 40.540 184.895 40.845 185.405 ;
        RECT 41.475 184.895 41.765 185.620 ;
        RECT 41.940 185.065 42.195 185.635 ;
        RECT 42.365 185.465 43.295 185.635 ;
        RECT 43.465 186.425 44.475 186.595 ;
        RECT 43.465 185.625 43.635 186.425 ;
        RECT 43.840 186.085 44.115 186.225 ;
        RECT 43.835 185.915 44.115 186.085 ;
        RECT 43.120 185.430 43.295 185.465 ;
        RECT 42.365 184.895 42.695 185.295 ;
        RECT 43.120 185.065 43.650 185.430 ;
        RECT 43.840 185.065 44.115 185.915 ;
        RECT 44.285 185.065 44.475 186.425 ;
        RECT 44.645 186.440 44.815 187.105 ;
        RECT 44.985 186.685 45.155 187.445 ;
        RECT 45.390 186.685 45.905 187.095 ;
        RECT 44.645 186.250 45.395 186.440 ;
        RECT 45.565 185.875 45.905 186.685 ;
        RECT 46.085 186.475 46.415 187.260 ;
        RECT 46.085 186.305 46.765 186.475 ;
        RECT 46.945 186.305 47.275 187.445 ;
        RECT 47.610 186.435 47.910 187.275 ;
        RECT 48.105 186.605 48.355 187.445 ;
        RECT 48.945 186.855 49.750 187.275 ;
        RECT 48.525 186.685 50.090 186.855 ;
        RECT 48.525 186.435 48.695 186.685 ;
        RECT 46.075 185.885 46.425 186.135 ;
        RECT 44.675 185.705 45.905 185.875 ;
        RECT 46.595 185.705 46.765 186.305 ;
        RECT 47.610 186.265 48.695 186.435 ;
        RECT 46.935 185.885 47.285 186.135 ;
        RECT 47.455 185.805 47.785 186.095 ;
        RECT 44.655 184.895 45.165 185.430 ;
        RECT 45.385 185.100 45.630 185.705 ;
        RECT 46.095 184.895 46.335 185.705 ;
        RECT 46.505 185.065 46.835 185.705 ;
        RECT 47.005 184.895 47.275 185.705 ;
        RECT 47.955 185.635 48.125 186.265 ;
        RECT 48.865 186.135 49.185 186.515 ;
        RECT 48.295 185.885 48.625 186.095 ;
        RECT 48.805 185.885 49.185 186.135 ;
        RECT 49.375 186.095 49.750 186.515 ;
        RECT 49.920 186.435 50.090 186.685 ;
        RECT 50.260 186.605 50.590 187.445 ;
        RECT 50.760 186.685 51.425 187.275 ;
        RECT 49.920 186.265 50.840 186.435 ;
        RECT 50.670 186.095 50.840 186.265 ;
        RECT 49.375 186.085 49.860 186.095 ;
        RECT 49.355 185.915 49.860 186.085 ;
        RECT 49.375 185.885 49.860 185.915 ;
        RECT 50.050 185.885 50.500 186.095 ;
        RECT 50.670 185.885 51.005 186.095 ;
        RECT 51.175 185.715 51.425 186.685 ;
        RECT 51.600 186.775 51.855 187.275 ;
        RECT 52.025 186.945 52.355 187.445 ;
        RECT 51.600 186.605 52.350 186.775 ;
        RECT 51.600 185.785 51.950 186.435 ;
        RECT 47.615 185.455 48.125 185.635 ;
        RECT 48.530 185.545 50.230 185.715 ;
        RECT 48.530 185.455 48.915 185.545 ;
        RECT 47.615 185.065 47.945 185.455 ;
        RECT 48.115 185.115 49.300 185.285 ;
        RECT 49.560 184.895 49.730 185.365 ;
        RECT 49.900 185.080 50.230 185.545 ;
        RECT 50.400 184.895 50.570 185.715 ;
        RECT 50.740 185.075 51.425 185.715 ;
        RECT 52.120 185.615 52.350 186.605 ;
        RECT 51.600 185.445 52.350 185.615 ;
        RECT 51.600 185.155 51.855 185.445 ;
        RECT 52.025 184.895 52.355 185.275 ;
        RECT 52.525 185.155 52.695 187.275 ;
        RECT 52.865 186.475 53.190 187.260 ;
        RECT 53.360 186.985 53.610 187.445 ;
        RECT 53.780 186.945 54.030 187.275 ;
        RECT 54.245 186.945 54.925 187.275 ;
        RECT 53.780 186.815 53.950 186.945 ;
        RECT 53.555 186.645 53.950 186.815 ;
        RECT 52.925 185.425 53.385 186.475 ;
        RECT 53.555 185.285 53.725 186.645 ;
        RECT 54.120 186.385 54.585 186.775 ;
        RECT 53.895 185.575 54.245 186.195 ;
        RECT 54.415 185.795 54.585 186.385 ;
        RECT 54.755 186.165 54.925 186.945 ;
        RECT 55.095 186.845 55.265 187.185 ;
        RECT 55.500 187.015 55.830 187.445 ;
        RECT 56.000 186.845 56.170 187.185 ;
        RECT 56.465 186.985 56.835 187.445 ;
        RECT 55.095 186.675 56.170 186.845 ;
        RECT 57.005 186.815 57.175 187.275 ;
        RECT 57.410 186.935 58.280 187.275 ;
        RECT 58.450 186.985 58.700 187.445 ;
        RECT 56.615 186.645 57.175 186.815 ;
        RECT 56.615 186.505 56.785 186.645 ;
        RECT 55.285 186.335 56.785 186.505 ;
        RECT 57.480 186.475 57.940 186.765 ;
        RECT 54.755 185.995 56.445 186.165 ;
        RECT 54.415 185.575 54.770 185.795 ;
        RECT 54.940 185.285 55.110 185.995 ;
        RECT 55.315 185.575 56.105 185.825 ;
        RECT 56.275 185.815 56.445 185.995 ;
        RECT 56.615 185.645 56.785 186.335 ;
        RECT 53.055 184.895 53.385 185.255 ;
        RECT 53.555 185.115 54.050 185.285 ;
        RECT 54.255 185.115 55.110 185.285 ;
        RECT 55.985 184.895 56.315 185.355 ;
        RECT 56.525 185.255 56.785 185.645 ;
        RECT 56.975 186.465 57.940 186.475 ;
        RECT 58.110 186.555 58.280 186.935 ;
        RECT 58.870 186.895 59.040 187.185 ;
        RECT 59.220 187.065 59.550 187.445 ;
        RECT 58.870 186.725 59.670 186.895 ;
        RECT 56.975 186.305 57.650 186.465 ;
        RECT 58.110 186.385 59.330 186.555 ;
        RECT 56.975 185.515 57.185 186.305 ;
        RECT 58.110 186.295 58.280 186.385 ;
        RECT 57.355 185.515 57.705 186.135 ;
        RECT 57.875 186.125 58.280 186.295 ;
        RECT 57.875 185.345 58.045 186.125 ;
        RECT 58.215 185.675 58.435 185.955 ;
        RECT 58.615 185.845 59.155 186.215 ;
        RECT 59.500 186.135 59.670 186.725 ;
        RECT 59.890 186.305 60.195 187.445 ;
        RECT 60.365 186.255 60.620 187.135 ;
        RECT 61.500 186.690 61.830 187.445 ;
        RECT 62.000 186.895 62.190 187.275 ;
        RECT 62.360 187.065 62.690 187.445 ;
        RECT 62.860 186.895 63.070 187.275 ;
        RECT 63.240 187.005 63.520 187.445 ;
        RECT 63.690 187.085 65.670 187.275 ;
        RECT 62.000 186.835 63.070 186.895 ;
        RECT 65.480 186.895 65.670 187.085 ;
        RECT 65.840 187.065 66.170 187.445 ;
        RECT 66.340 186.895 66.575 187.275 ;
        RECT 62.000 186.665 65.310 186.835 ;
        RECT 65.480 186.725 66.575 186.895 ;
        RECT 62.000 186.510 63.215 186.665 ;
        RECT 66.745 186.630 67.030 187.445 ;
        RECT 59.500 186.105 60.240 186.135 ;
        RECT 58.215 185.505 58.745 185.675 ;
        RECT 56.525 185.085 56.875 185.255 ;
        RECT 57.095 185.065 58.045 185.345 ;
        RECT 58.215 184.895 58.405 185.335 ;
        RECT 58.575 185.275 58.745 185.505 ;
        RECT 58.915 185.445 59.155 185.845 ;
        RECT 59.325 185.805 60.240 186.105 ;
        RECT 59.325 185.630 59.650 185.805 ;
        RECT 59.325 185.275 59.645 185.630 ;
        RECT 60.410 185.605 60.620 186.255 ;
        RECT 58.575 185.105 59.645 185.275 ;
        RECT 59.890 184.895 60.195 185.355 ;
        RECT 60.365 185.075 60.620 185.605 ;
        RECT 61.315 186.255 63.215 186.510 ;
        RECT 63.455 186.325 66.575 186.495 ;
        RECT 61.315 185.655 61.725 186.255 ;
        RECT 61.895 185.825 63.245 186.085 ;
        RECT 63.455 185.800 63.705 186.325 ;
        RECT 63.875 185.880 65.165 186.155 ;
        RECT 65.675 186.130 66.575 186.325 ;
        RECT 67.235 186.280 67.525 187.445 ;
        RECT 67.695 186.745 68.055 187.445 ;
        RECT 68.585 186.915 68.915 187.255 ;
        RECT 69.445 187.085 70.115 187.445 ;
        RECT 70.285 186.915 70.475 187.275 ;
        RECT 70.645 187.065 70.995 187.445 ;
        RECT 68.585 186.895 70.475 186.915 ;
        RECT 68.585 186.685 71.005 186.895 ;
        RECT 70.285 186.640 71.005 186.685 ;
        RECT 67.730 186.305 69.650 186.515 ;
        RECT 65.675 185.825 67.025 186.130 ;
        RECT 67.730 185.805 68.100 186.305 ;
        RECT 68.440 185.805 68.990 186.135 ;
        RECT 69.345 185.800 69.650 186.305 ;
        RECT 69.975 185.885 70.645 186.425 ;
        RECT 70.815 186.145 71.005 186.640 ;
        RECT 71.175 186.510 71.355 187.275 ;
        RECT 71.525 186.680 71.855 187.445 ;
        RECT 72.025 186.510 72.215 187.275 ;
        RECT 72.385 186.680 72.715 187.445 ;
        RECT 71.175 186.340 73.040 186.510 ;
        RECT 70.815 185.805 72.640 186.145 ;
        RECT 70.815 185.680 71.015 185.805 ;
        RECT 61.315 185.425 63.120 185.655 ;
        RECT 63.290 185.425 67.030 185.630 ;
        RECT 63.290 185.255 63.520 185.425 ;
        RECT 61.500 185.065 63.520 185.255 ;
        RECT 63.690 184.895 64.020 185.255 ;
        RECT 64.550 184.895 64.880 185.255 ;
        RECT 65.410 184.895 65.740 185.255 ;
        RECT 66.270 184.895 66.600 185.255 ;
        RECT 67.235 184.895 67.525 185.620 ;
        RECT 67.725 185.425 69.855 185.595 ;
        RECT 70.035 185.465 71.015 185.680 ;
        RECT 72.810 185.615 73.040 186.340 ;
        RECT 73.225 186.465 73.555 187.275 ;
        RECT 73.725 186.645 73.965 187.445 ;
        RECT 73.225 186.295 73.940 186.465 ;
        RECT 73.220 185.885 73.600 186.125 ;
        RECT 73.770 186.055 73.940 186.295 ;
        RECT 74.145 186.425 74.315 187.275 ;
        RECT 74.485 186.645 74.815 187.445 ;
        RECT 74.985 186.425 75.155 187.275 ;
        RECT 74.145 186.255 75.155 186.425 ;
        RECT 75.325 186.295 75.655 187.445 ;
        RECT 75.975 186.305 76.265 187.445 ;
        RECT 76.435 186.725 76.885 187.275 ;
        RECT 77.075 186.725 77.405 187.445 ;
        RECT 73.770 185.885 74.270 186.055 ;
        RECT 73.770 185.715 73.940 185.885 ;
        RECT 74.660 185.715 75.155 186.255 ;
        RECT 71.415 185.445 73.040 185.615 ;
        RECT 73.305 185.545 73.940 185.715 ;
        RECT 74.145 185.545 75.155 185.715 ;
        RECT 71.415 185.425 72.535 185.445 ;
        RECT 69.525 185.295 69.855 185.425 ;
        RECT 68.155 184.895 68.485 185.255 ;
        RECT 69.015 184.895 69.355 185.255 ;
        RECT 69.525 185.065 70.795 185.295 ;
        RECT 70.985 184.895 71.315 185.275 ;
        RECT 71.845 184.895 72.175 185.255 ;
        RECT 72.705 184.895 73.035 185.275 ;
        RECT 73.305 185.065 73.475 185.545 ;
        RECT 73.655 184.895 73.895 185.375 ;
        RECT 74.145 185.065 74.315 185.545 ;
        RECT 74.485 184.895 74.815 185.375 ;
        RECT 74.985 185.065 75.155 185.545 ;
        RECT 75.325 184.895 75.655 185.695 ;
        RECT 75.975 184.895 76.265 185.695 ;
        RECT 76.435 185.355 76.685 186.725 ;
        RECT 77.615 186.555 77.915 187.105 ;
        RECT 78.085 186.775 78.365 187.445 ;
        RECT 76.975 186.385 77.915 186.555 ;
        RECT 76.975 186.135 77.145 186.385 ;
        RECT 78.250 186.135 78.565 186.575 ;
        RECT 76.855 185.805 77.145 186.135 ;
        RECT 77.315 185.885 77.645 186.135 ;
        RECT 77.875 185.885 78.565 186.135 ;
        RECT 78.735 186.475 79.045 187.275 ;
        RECT 79.215 186.645 79.525 187.445 ;
        RECT 79.695 186.815 79.955 187.275 ;
        RECT 80.125 186.985 80.380 187.445 ;
        RECT 80.555 186.815 80.815 187.275 ;
        RECT 79.695 186.645 80.815 186.815 ;
        RECT 78.735 186.305 79.765 186.475 ;
        RECT 76.975 185.715 77.145 185.805 ;
        RECT 76.975 185.525 78.365 185.715 ;
        RECT 76.435 185.065 76.985 185.355 ;
        RECT 77.155 184.895 77.405 185.355 ;
        RECT 78.035 185.165 78.365 185.525 ;
        RECT 78.735 185.395 78.905 186.305 ;
        RECT 79.075 185.565 79.425 186.135 ;
        RECT 79.595 186.055 79.765 186.305 ;
        RECT 80.555 186.395 80.815 186.645 ;
        RECT 80.985 186.575 81.270 187.445 ;
        RECT 81.495 186.475 81.805 187.275 ;
        RECT 81.975 186.645 82.285 187.445 ;
        RECT 82.455 186.815 82.715 187.275 ;
        RECT 82.885 186.985 83.140 187.445 ;
        RECT 83.315 186.815 83.575 187.275 ;
        RECT 82.455 186.645 83.575 186.815 ;
        RECT 80.555 186.225 81.310 186.395 ;
        RECT 79.595 185.885 80.735 186.055 ;
        RECT 80.905 185.715 81.310 186.225 ;
        RECT 79.660 185.545 81.310 185.715 ;
        RECT 81.495 186.305 82.525 186.475 ;
        RECT 78.735 185.065 79.035 185.395 ;
        RECT 79.205 184.895 79.480 185.375 ;
        RECT 79.660 185.155 79.955 185.545 ;
        RECT 80.125 184.895 80.380 185.375 ;
        RECT 80.555 185.155 80.815 185.545 ;
        RECT 81.495 185.395 81.665 186.305 ;
        RECT 81.835 185.565 82.185 186.135 ;
        RECT 82.355 186.055 82.525 186.305 ;
        RECT 83.315 186.395 83.575 186.645 ;
        RECT 83.745 186.575 84.030 187.445 ;
        RECT 84.255 187.010 89.600 187.445 ;
        RECT 83.315 186.225 84.070 186.395 ;
        RECT 82.355 185.885 83.495 186.055 ;
        RECT 83.665 185.715 84.070 186.225 ;
        RECT 82.420 185.545 84.070 185.715 ;
        RECT 80.985 184.895 81.265 185.375 ;
        RECT 81.495 185.065 81.795 185.395 ;
        RECT 81.965 184.895 82.240 185.375 ;
        RECT 82.420 185.155 82.715 185.545 ;
        RECT 82.885 184.895 83.140 185.375 ;
        RECT 83.315 185.155 83.575 185.545 ;
        RECT 85.840 185.440 86.180 186.270 ;
        RECT 87.660 185.760 88.010 187.010 ;
        RECT 89.775 186.355 92.365 187.445 ;
        RECT 89.775 185.665 90.985 186.185 ;
        RECT 91.155 185.835 92.365 186.355 ;
        RECT 92.995 186.280 93.285 187.445 ;
        RECT 93.510 186.575 93.795 187.445 ;
        RECT 93.965 186.815 94.225 187.275 ;
        RECT 94.400 186.985 94.655 187.445 ;
        RECT 94.825 186.815 95.085 187.275 ;
        RECT 93.965 186.645 95.085 186.815 ;
        RECT 95.255 186.645 95.565 187.445 ;
        RECT 93.965 186.395 94.225 186.645 ;
        RECT 95.735 186.475 96.045 187.275 ;
        RECT 93.470 186.225 94.225 186.395 ;
        RECT 95.015 186.305 96.045 186.475 ;
        RECT 96.215 186.355 97.425 187.445 ;
        RECT 97.595 186.890 98.200 187.445 ;
        RECT 98.375 186.935 98.855 187.275 ;
        RECT 99.025 186.900 99.280 187.445 ;
        RECT 97.595 186.790 98.210 186.890 ;
        RECT 98.025 186.765 98.210 186.790 ;
        RECT 93.470 185.715 93.875 186.225 ;
        RECT 95.015 186.055 95.185 186.305 ;
        RECT 94.045 185.885 95.185 186.055 ;
        RECT 83.745 184.895 84.025 185.375 ;
        RECT 84.255 184.895 89.600 185.440 ;
        RECT 89.775 184.895 92.365 185.665 ;
        RECT 92.995 184.895 93.285 185.620 ;
        RECT 93.470 185.545 95.120 185.715 ;
        RECT 95.355 185.565 95.705 186.135 ;
        RECT 93.515 184.895 93.795 185.375 ;
        RECT 93.965 185.155 94.225 185.545 ;
        RECT 94.400 184.895 94.655 185.375 ;
        RECT 94.825 185.155 95.120 185.545 ;
        RECT 95.875 185.395 96.045 186.305 ;
        RECT 95.300 184.895 95.575 185.375 ;
        RECT 95.745 185.065 96.045 185.395 ;
        RECT 96.215 185.645 96.735 186.185 ;
        RECT 96.905 185.815 97.425 186.355 ;
        RECT 97.595 186.170 97.855 186.620 ;
        RECT 98.025 186.520 98.355 186.765 ;
        RECT 98.525 186.445 99.280 186.695 ;
        RECT 99.450 186.575 99.725 187.275 ;
        RECT 98.510 186.410 99.280 186.445 ;
        RECT 98.495 186.400 99.280 186.410 ;
        RECT 98.490 186.385 99.385 186.400 ;
        RECT 98.470 186.370 99.385 186.385 ;
        RECT 98.450 186.360 99.385 186.370 ;
        RECT 98.425 186.350 99.385 186.360 ;
        RECT 98.355 186.320 99.385 186.350 ;
        RECT 98.335 186.290 99.385 186.320 ;
        RECT 98.315 186.260 99.385 186.290 ;
        RECT 98.285 186.235 99.385 186.260 ;
        RECT 98.250 186.200 99.385 186.235 ;
        RECT 98.220 186.195 99.385 186.200 ;
        RECT 98.220 186.190 98.610 186.195 ;
        RECT 98.220 186.180 98.585 186.190 ;
        RECT 98.220 186.175 98.570 186.180 ;
        RECT 98.220 186.170 98.555 186.175 ;
        RECT 97.595 186.165 98.555 186.170 ;
        RECT 97.595 186.155 98.545 186.165 ;
        RECT 97.595 186.150 98.535 186.155 ;
        RECT 97.595 186.140 98.525 186.150 ;
        RECT 97.595 186.130 98.520 186.140 ;
        RECT 97.595 186.125 98.515 186.130 ;
        RECT 97.595 186.110 98.505 186.125 ;
        RECT 97.595 186.095 98.500 186.110 ;
        RECT 97.595 186.070 98.490 186.095 ;
        RECT 97.595 186.000 98.485 186.070 ;
        RECT 96.215 184.895 97.425 185.645 ;
        RECT 97.595 185.445 98.145 185.830 ;
        RECT 98.315 185.275 98.485 186.000 ;
        RECT 97.595 185.105 98.485 185.275 ;
        RECT 98.655 185.600 98.985 186.025 ;
        RECT 99.155 185.800 99.385 186.195 ;
        RECT 98.655 185.115 98.875 185.600 ;
        RECT 99.555 185.545 99.725 186.575 ;
        RECT 99.045 184.895 99.295 185.435 ;
        RECT 99.465 185.065 99.725 185.545 ;
        RECT 99.905 185.075 100.165 187.265 ;
        RECT 100.335 186.715 100.675 187.445 ;
        RECT 100.855 186.535 101.125 187.265 ;
        RECT 100.355 186.315 101.125 186.535 ;
        RECT 101.305 186.555 101.535 187.265 ;
        RECT 101.705 186.735 102.035 187.445 ;
        RECT 102.205 186.555 102.465 187.265 ;
        RECT 101.305 186.315 102.465 186.555 ;
        RECT 102.655 186.355 104.325 187.445 ;
        RECT 100.355 185.645 100.645 186.315 ;
        RECT 100.825 185.825 101.290 186.135 ;
        RECT 101.470 185.825 101.995 186.135 ;
        RECT 100.355 185.445 101.585 185.645 ;
        RECT 100.425 184.895 101.095 185.265 ;
        RECT 101.275 185.075 101.585 185.445 ;
        RECT 101.765 185.185 101.995 185.825 ;
        RECT 102.175 185.805 102.475 186.135 ;
        RECT 102.655 185.665 103.405 186.185 ;
        RECT 103.575 185.835 104.325 186.355 ;
        RECT 104.965 186.835 105.295 187.265 ;
        RECT 105.475 187.005 105.670 187.445 ;
        RECT 105.840 186.835 106.170 187.265 ;
        RECT 104.965 186.665 106.170 186.835 ;
        RECT 104.965 186.335 105.860 186.665 ;
        RECT 106.340 186.495 106.615 187.265 ;
        RECT 106.030 186.305 106.615 186.495 ;
        RECT 106.795 186.355 110.305 187.445 ;
        RECT 110.475 186.355 111.685 187.445 ;
        RECT 111.860 186.935 113.515 187.225 ;
        RECT 104.970 185.805 105.265 186.135 ;
        RECT 105.445 185.805 105.860 186.135 ;
        RECT 102.175 184.895 102.465 185.625 ;
        RECT 102.655 184.895 104.325 185.665 ;
        RECT 104.965 184.895 105.265 185.625 ;
        RECT 105.445 185.185 105.675 185.805 ;
        RECT 106.030 185.635 106.205 186.305 ;
        RECT 105.875 185.455 106.205 185.635 ;
        RECT 106.375 185.485 106.615 186.135 ;
        RECT 106.795 185.665 108.445 186.185 ;
        RECT 108.615 185.835 110.305 186.355 ;
        RECT 105.875 185.075 106.100 185.455 ;
        RECT 106.270 184.895 106.600 185.285 ;
        RECT 106.795 184.895 110.305 185.665 ;
        RECT 110.475 185.645 110.995 186.185 ;
        RECT 111.165 185.815 111.685 186.355 ;
        RECT 111.860 186.595 113.450 186.765 ;
        RECT 113.685 186.645 113.965 187.445 ;
        RECT 111.860 186.305 112.180 186.595 ;
        RECT 113.280 186.475 113.450 186.595 ;
        RECT 110.475 184.895 111.685 185.645 ;
        RECT 111.860 185.565 112.210 186.135 ;
        RECT 112.380 185.805 113.090 186.425 ;
        RECT 113.280 186.305 114.005 186.475 ;
        RECT 114.175 186.305 114.445 187.275 ;
        RECT 114.625 186.495 114.900 187.265 ;
        RECT 115.070 186.835 115.400 187.265 ;
        RECT 115.570 187.005 115.765 187.445 ;
        RECT 115.945 186.835 116.275 187.265 ;
        RECT 115.070 186.665 116.275 186.835 ;
        RECT 114.625 186.305 115.210 186.495 ;
        RECT 115.380 186.335 116.275 186.665 ;
        RECT 116.455 186.305 116.715 187.445 ;
        RECT 113.835 186.135 114.005 186.305 ;
        RECT 113.260 185.805 113.665 186.135 ;
        RECT 113.835 185.805 114.105 186.135 ;
        RECT 113.835 185.635 114.005 185.805 ;
        RECT 112.395 185.465 114.005 185.635 ;
        RECT 114.275 185.570 114.445 186.305 ;
        RECT 111.865 184.895 112.195 185.395 ;
        RECT 112.395 185.115 112.565 185.465 ;
        RECT 112.765 184.895 113.095 185.295 ;
        RECT 113.265 185.115 113.435 185.465 ;
        RECT 113.605 184.895 113.985 185.295 ;
        RECT 114.175 185.225 114.445 185.570 ;
        RECT 114.625 185.485 114.865 186.135 ;
        RECT 115.035 185.635 115.210 186.305 ;
        RECT 116.885 186.295 117.215 187.275 ;
        RECT 117.385 186.305 117.665 187.445 ;
        RECT 115.380 185.805 115.795 186.135 ;
        RECT 115.975 185.805 116.270 186.135 ;
        RECT 116.475 185.885 116.810 186.135 ;
        RECT 115.035 185.455 115.365 185.635 ;
        RECT 114.640 184.895 114.970 185.285 ;
        RECT 115.140 185.075 115.365 185.455 ;
        RECT 115.565 185.185 115.795 185.805 ;
        RECT 116.980 185.745 117.150 186.295 ;
        RECT 118.755 186.280 119.045 187.445 ;
        RECT 119.215 186.355 120.885 187.445 ;
        RECT 121.060 187.065 121.395 187.445 ;
        RECT 117.320 185.865 117.655 186.135 ;
        RECT 116.975 185.695 117.150 185.745 ;
        RECT 115.975 184.895 116.275 185.625 ;
        RECT 116.455 185.065 117.150 185.695 ;
        RECT 117.355 184.895 117.665 185.695 ;
        RECT 119.215 185.665 119.965 186.185 ;
        RECT 120.135 185.835 120.885 186.355 ;
        RECT 118.755 184.895 119.045 185.620 ;
        RECT 119.215 184.895 120.885 185.665 ;
        RECT 121.055 185.575 121.295 186.885 ;
        RECT 121.565 186.475 121.815 187.275 ;
        RECT 122.035 186.725 122.365 187.445 ;
        RECT 122.550 186.475 122.800 187.275 ;
        RECT 123.265 186.645 123.595 187.445 ;
        RECT 123.765 187.015 124.105 187.275 ;
        RECT 121.465 186.305 123.655 186.475 ;
        RECT 121.465 185.395 121.635 186.305 ;
        RECT 123.340 186.135 123.655 186.305 ;
        RECT 121.140 185.065 121.635 185.395 ;
        RECT 121.855 185.170 122.205 186.135 ;
        RECT 122.385 185.165 122.685 186.135 ;
        RECT 122.865 185.165 123.145 186.135 ;
        RECT 123.340 185.885 123.670 186.135 ;
        RECT 123.325 184.895 123.595 185.695 ;
        RECT 123.845 185.615 124.105 187.015 ;
        RECT 125.205 186.645 125.535 187.445 ;
        RECT 125.715 187.105 127.145 187.275 ;
        RECT 125.715 186.475 125.965 187.105 ;
        RECT 123.765 185.105 124.105 185.615 ;
        RECT 125.195 186.305 125.965 186.475 ;
        RECT 125.195 185.635 125.365 186.305 ;
        RECT 125.535 185.805 125.940 186.135 ;
        RECT 126.155 185.805 126.405 186.935 ;
        RECT 126.605 186.135 126.805 186.935 ;
        RECT 126.975 186.425 127.145 187.105 ;
        RECT 127.315 186.595 127.630 187.445 ;
        RECT 127.805 186.645 128.245 187.275 ;
        RECT 128.415 187.010 133.760 187.445 ;
        RECT 126.975 186.255 127.765 186.425 ;
        RECT 126.605 185.805 126.850 186.135 ;
        RECT 127.035 185.805 127.425 186.085 ;
        RECT 127.595 185.805 127.765 186.255 ;
        RECT 127.935 185.635 128.245 186.645 ;
        RECT 125.195 185.065 125.685 185.635 ;
        RECT 125.855 185.465 127.015 185.635 ;
        RECT 125.855 185.065 126.085 185.465 ;
        RECT 126.255 184.895 126.675 185.295 ;
        RECT 126.845 185.065 127.015 185.465 ;
        RECT 127.185 184.895 127.635 185.635 ;
        RECT 127.805 185.075 128.245 185.635 ;
        RECT 130.000 185.440 130.340 186.270 ;
        RECT 131.820 185.760 132.170 187.010 ;
        RECT 133.945 186.475 134.275 187.260 ;
        RECT 133.945 186.305 134.625 186.475 ;
        RECT 134.805 186.305 135.135 187.445 ;
        RECT 135.315 186.355 138.825 187.445 ;
        RECT 138.995 186.355 140.205 187.445 ;
        RECT 140.375 186.890 140.980 187.445 ;
        RECT 141.155 186.935 141.635 187.275 ;
        RECT 141.805 186.900 142.060 187.445 ;
        RECT 140.375 186.790 140.990 186.890 ;
        RECT 140.805 186.765 140.990 186.790 ;
        RECT 133.935 185.885 134.285 186.135 ;
        RECT 134.455 185.705 134.625 186.305 ;
        RECT 134.795 185.885 135.145 186.135 ;
        RECT 128.415 184.895 133.760 185.440 ;
        RECT 133.955 184.895 134.195 185.705 ;
        RECT 134.365 185.065 134.695 185.705 ;
        RECT 134.865 184.895 135.135 185.705 ;
        RECT 135.315 185.665 136.965 186.185 ;
        RECT 137.135 185.835 138.825 186.355 ;
        RECT 135.315 184.895 138.825 185.665 ;
        RECT 138.995 185.645 139.515 186.185 ;
        RECT 139.685 185.815 140.205 186.355 ;
        RECT 140.375 186.170 140.635 186.620 ;
        RECT 140.805 186.520 141.135 186.765 ;
        RECT 141.305 186.445 142.060 186.695 ;
        RECT 142.230 186.575 142.505 187.275 ;
        RECT 141.290 186.410 142.060 186.445 ;
        RECT 141.275 186.400 142.060 186.410 ;
        RECT 141.270 186.385 142.165 186.400 ;
        RECT 141.250 186.370 142.165 186.385 ;
        RECT 141.230 186.360 142.165 186.370 ;
        RECT 141.205 186.350 142.165 186.360 ;
        RECT 141.135 186.320 142.165 186.350 ;
        RECT 141.115 186.290 142.165 186.320 ;
        RECT 141.095 186.260 142.165 186.290 ;
        RECT 141.065 186.235 142.165 186.260 ;
        RECT 141.030 186.200 142.165 186.235 ;
        RECT 141.000 186.195 142.165 186.200 ;
        RECT 141.000 186.190 141.390 186.195 ;
        RECT 141.000 186.180 141.365 186.190 ;
        RECT 141.000 186.175 141.350 186.180 ;
        RECT 141.000 186.170 141.335 186.175 ;
        RECT 140.375 186.165 141.335 186.170 ;
        RECT 140.375 186.155 141.325 186.165 ;
        RECT 140.375 186.150 141.315 186.155 ;
        RECT 140.375 186.140 141.305 186.150 ;
        RECT 140.375 186.130 141.300 186.140 ;
        RECT 140.375 186.125 141.295 186.130 ;
        RECT 140.375 186.110 141.285 186.125 ;
        RECT 140.375 186.095 141.280 186.110 ;
        RECT 140.375 186.070 141.270 186.095 ;
        RECT 140.375 186.000 141.265 186.070 ;
        RECT 138.995 184.895 140.205 185.645 ;
        RECT 140.375 185.445 140.925 185.830 ;
        RECT 141.095 185.275 141.265 186.000 ;
        RECT 140.375 185.105 141.265 185.275 ;
        RECT 141.435 185.600 141.765 186.025 ;
        RECT 141.935 185.800 142.165 186.195 ;
        RECT 141.435 185.115 141.655 185.600 ;
        RECT 142.335 185.545 142.505 186.575 ;
        RECT 142.675 186.355 144.345 187.445 ;
        RECT 141.825 184.895 142.075 185.435 ;
        RECT 142.245 185.065 142.505 185.545 ;
        RECT 142.675 185.665 143.425 186.185 ;
        RECT 143.595 185.835 144.345 186.355 ;
        RECT 144.515 186.280 144.805 187.445 ;
        RECT 144.975 187.010 150.320 187.445 ;
        RECT 142.675 184.895 144.345 185.665 ;
        RECT 144.515 184.895 144.805 185.620 ;
        RECT 146.560 185.440 146.900 186.270 ;
        RECT 148.380 185.760 148.730 187.010 ;
        RECT 150.495 186.355 152.165 187.445 ;
        RECT 150.495 185.665 151.245 186.185 ;
        RECT 151.415 185.835 152.165 186.355 ;
        RECT 152.335 186.475 152.645 187.275 ;
        RECT 152.815 186.645 153.125 187.445 ;
        RECT 153.295 186.815 153.555 187.275 ;
        RECT 153.725 186.985 153.980 187.445 ;
        RECT 154.155 186.815 154.415 187.275 ;
        RECT 153.295 186.645 154.415 186.815 ;
        RECT 152.335 186.305 153.365 186.475 ;
        RECT 144.975 184.895 150.320 185.440 ;
        RECT 150.495 184.895 152.165 185.665 ;
        RECT 152.335 185.395 152.505 186.305 ;
        RECT 152.675 185.565 153.025 186.135 ;
        RECT 153.195 186.055 153.365 186.305 ;
        RECT 154.155 186.395 154.415 186.645 ;
        RECT 154.585 186.575 154.870 187.445 ;
        RECT 154.155 186.225 154.910 186.395 ;
        RECT 155.095 186.355 156.765 187.445 ;
        RECT 153.195 185.885 154.335 186.055 ;
        RECT 154.505 185.715 154.910 186.225 ;
        RECT 153.260 185.545 154.910 185.715 ;
        RECT 155.095 185.665 155.845 186.185 ;
        RECT 156.015 185.835 156.765 186.355 ;
        RECT 156.935 186.355 158.145 187.445 ;
        RECT 156.935 185.815 157.455 186.355 ;
        RECT 152.335 185.065 152.635 185.395 ;
        RECT 152.805 184.895 153.080 185.375 ;
        RECT 153.260 185.155 153.555 185.545 ;
        RECT 153.725 184.895 153.980 185.375 ;
        RECT 154.155 185.155 154.415 185.545 ;
        RECT 154.585 184.895 154.865 185.375 ;
        RECT 155.095 184.895 156.765 185.665 ;
        RECT 157.625 185.645 158.145 186.185 ;
        RECT 156.935 184.895 158.145 185.645 ;
        RECT 2.750 184.725 158.230 184.895 ;
        RECT 2.835 183.975 4.045 184.725 ;
        RECT 2.835 183.435 3.355 183.975 ;
        RECT 4.215 183.955 6.805 184.725 ;
        RECT 6.975 184.050 7.235 184.555 ;
        RECT 7.415 184.345 7.745 184.725 ;
        RECT 7.925 184.175 8.095 184.555 ;
        RECT 3.525 183.265 4.045 183.805 ;
        RECT 4.215 183.435 5.425 183.955 ;
        RECT 5.595 183.265 6.805 183.785 ;
        RECT 2.835 182.175 4.045 183.265 ;
        RECT 4.215 182.175 6.805 183.265 ;
        RECT 6.975 183.250 7.145 184.050 ;
        RECT 7.430 184.005 8.095 184.175 ;
        RECT 7.430 183.750 7.600 184.005 ;
        RECT 8.360 183.985 8.615 184.555 ;
        RECT 8.785 184.325 9.115 184.725 ;
        RECT 9.540 184.190 10.070 184.555 ;
        RECT 9.540 184.155 9.715 184.190 ;
        RECT 8.785 183.985 9.715 184.155 ;
        RECT 7.315 183.420 7.600 183.750 ;
        RECT 7.835 183.455 8.165 183.825 ;
        RECT 7.430 183.275 7.600 183.420 ;
        RECT 8.360 183.315 8.530 183.985 ;
        RECT 8.785 183.815 8.955 183.985 ;
        RECT 8.700 183.485 8.955 183.815 ;
        RECT 9.180 183.485 9.375 183.815 ;
        RECT 6.975 182.345 7.245 183.250 ;
        RECT 7.430 183.105 8.095 183.275 ;
        RECT 7.415 182.175 7.745 182.935 ;
        RECT 7.925 182.345 8.095 183.105 ;
        RECT 8.360 182.345 8.695 183.315 ;
        RECT 8.865 182.175 9.035 183.315 ;
        RECT 9.205 182.515 9.375 183.485 ;
        RECT 9.545 182.855 9.715 183.985 ;
        RECT 9.885 183.195 10.055 183.995 ;
        RECT 10.260 183.705 10.535 184.555 ;
        RECT 10.255 183.535 10.535 183.705 ;
        RECT 10.260 183.395 10.535 183.535 ;
        RECT 10.705 183.195 10.895 184.555 ;
        RECT 11.075 184.190 11.585 184.725 ;
        RECT 11.805 183.915 12.050 184.520 ;
        RECT 12.770 183.915 13.015 184.520 ;
        RECT 13.235 184.190 13.745 184.725 ;
        RECT 11.095 183.745 12.325 183.915 ;
        RECT 9.885 183.025 10.895 183.195 ;
        RECT 11.065 183.180 11.815 183.370 ;
        RECT 9.545 182.685 10.670 182.855 ;
        RECT 11.065 182.515 11.235 183.180 ;
        RECT 11.985 182.935 12.325 183.745 ;
        RECT 9.205 182.345 11.235 182.515 ;
        RECT 11.405 182.175 11.575 182.935 ;
        RECT 11.810 182.525 12.325 182.935 ;
        RECT 12.495 183.745 13.725 183.915 ;
        RECT 12.495 182.935 12.835 183.745 ;
        RECT 13.005 183.180 13.755 183.370 ;
        RECT 12.495 182.525 13.010 182.935 ;
        RECT 13.245 182.175 13.415 182.935 ;
        RECT 13.585 182.515 13.755 183.180 ;
        RECT 13.925 183.195 14.115 184.555 ;
        RECT 14.285 183.705 14.560 184.555 ;
        RECT 14.750 184.190 15.280 184.555 ;
        RECT 15.705 184.325 16.035 184.725 ;
        RECT 15.105 184.155 15.280 184.190 ;
        RECT 14.285 183.535 14.565 183.705 ;
        RECT 14.285 183.395 14.560 183.535 ;
        RECT 14.765 183.195 14.935 183.995 ;
        RECT 13.925 183.025 14.935 183.195 ;
        RECT 15.105 183.985 16.035 184.155 ;
        RECT 16.205 183.985 16.460 184.555 ;
        RECT 15.105 182.855 15.275 183.985 ;
        RECT 15.865 183.815 16.035 183.985 ;
        RECT 14.150 182.685 15.275 182.855 ;
        RECT 15.445 183.485 15.640 183.815 ;
        RECT 15.865 183.485 16.120 183.815 ;
        RECT 15.445 182.515 15.615 183.485 ;
        RECT 16.290 183.315 16.460 183.985 ;
        RECT 16.685 183.970 16.935 184.725 ;
        RECT 17.105 184.015 17.355 184.545 ;
        RECT 17.525 184.265 17.830 184.725 ;
        RECT 18.075 184.345 19.145 184.515 ;
        RECT 17.105 183.365 17.310 184.015 ;
        RECT 18.075 183.990 18.395 184.345 ;
        RECT 18.070 183.815 18.395 183.990 ;
        RECT 17.480 183.515 18.395 183.815 ;
        RECT 18.565 183.775 18.805 184.175 ;
        RECT 18.975 184.115 19.145 184.345 ;
        RECT 19.315 184.285 19.505 184.725 ;
        RECT 19.675 184.275 20.625 184.555 ;
        RECT 20.845 184.365 21.195 184.535 ;
        RECT 18.975 183.945 19.505 184.115 ;
        RECT 17.480 183.485 18.220 183.515 ;
        RECT 13.585 182.345 15.615 182.515 ;
        RECT 15.785 182.175 15.955 183.315 ;
        RECT 16.125 182.345 16.460 183.315 ;
        RECT 16.685 182.175 16.935 183.315 ;
        RECT 17.105 182.485 17.355 183.365 ;
        RECT 17.525 182.175 17.830 183.315 ;
        RECT 18.050 182.895 18.220 183.485 ;
        RECT 18.565 183.405 19.105 183.775 ;
        RECT 19.285 183.665 19.505 183.945 ;
        RECT 19.675 183.495 19.845 184.275 ;
        RECT 19.440 183.325 19.845 183.495 ;
        RECT 20.015 183.485 20.365 184.105 ;
        RECT 19.440 183.235 19.610 183.325 ;
        RECT 20.535 183.315 20.745 184.105 ;
        RECT 18.390 183.065 19.610 183.235 ;
        RECT 20.070 183.155 20.745 183.315 ;
        RECT 18.050 182.725 18.850 182.895 ;
        RECT 18.170 182.175 18.500 182.555 ;
        RECT 18.680 182.435 18.850 182.725 ;
        RECT 19.440 182.685 19.610 183.065 ;
        RECT 19.780 183.145 20.745 183.155 ;
        RECT 20.935 183.975 21.195 184.365 ;
        RECT 21.405 184.265 21.735 184.725 ;
        RECT 22.610 184.335 23.465 184.505 ;
        RECT 23.670 184.335 24.165 184.505 ;
        RECT 24.335 184.365 24.665 184.725 ;
        RECT 20.935 183.285 21.105 183.975 ;
        RECT 21.275 183.625 21.445 183.805 ;
        RECT 21.615 183.795 22.405 184.045 ;
        RECT 22.610 183.625 22.780 184.335 ;
        RECT 22.950 183.825 23.305 184.045 ;
        RECT 21.275 183.455 22.965 183.625 ;
        RECT 19.780 182.855 20.240 183.145 ;
        RECT 20.935 183.115 22.435 183.285 ;
        RECT 20.935 182.975 21.105 183.115 ;
        RECT 20.545 182.805 21.105 182.975 ;
        RECT 19.020 182.175 19.270 182.635 ;
        RECT 19.440 182.345 20.310 182.685 ;
        RECT 20.545 182.345 20.715 182.805 ;
        RECT 21.550 182.775 22.625 182.945 ;
        RECT 20.885 182.175 21.255 182.635 ;
        RECT 21.550 182.435 21.720 182.775 ;
        RECT 21.890 182.175 22.220 182.605 ;
        RECT 22.455 182.435 22.625 182.775 ;
        RECT 22.795 182.675 22.965 183.455 ;
        RECT 23.135 183.235 23.305 183.825 ;
        RECT 23.475 183.425 23.825 184.045 ;
        RECT 23.135 182.845 23.600 183.235 ;
        RECT 23.995 182.975 24.165 184.335 ;
        RECT 24.335 183.145 24.795 184.195 ;
        RECT 23.770 182.805 24.165 182.975 ;
        RECT 23.770 182.675 23.940 182.805 ;
        RECT 22.795 182.345 23.475 182.675 ;
        RECT 23.690 182.345 23.940 182.675 ;
        RECT 24.110 182.175 24.360 182.635 ;
        RECT 24.530 182.360 24.855 183.145 ;
        RECT 25.025 182.345 25.195 184.465 ;
        RECT 25.365 184.345 25.695 184.725 ;
        RECT 25.865 184.175 26.120 184.465 ;
        RECT 25.370 184.005 26.120 184.175 ;
        RECT 27.215 184.050 27.475 184.555 ;
        RECT 27.655 184.345 27.985 184.725 ;
        RECT 28.165 184.175 28.335 184.555 ;
        RECT 25.370 183.015 25.600 184.005 ;
        RECT 25.770 183.185 26.120 183.835 ;
        RECT 27.215 183.250 27.385 184.050 ;
        RECT 27.670 184.005 28.335 184.175 ;
        RECT 27.670 183.750 27.840 184.005 ;
        RECT 28.595 184.000 28.885 184.725 ;
        RECT 29.060 183.985 29.315 184.555 ;
        RECT 29.485 184.325 29.815 184.725 ;
        RECT 30.240 184.190 30.770 184.555 ;
        RECT 30.240 184.155 30.415 184.190 ;
        RECT 29.485 183.985 30.415 184.155 ;
        RECT 27.555 183.420 27.840 183.750 ;
        RECT 28.075 183.455 28.405 183.825 ;
        RECT 27.670 183.275 27.840 183.420 ;
        RECT 25.370 182.845 26.120 183.015 ;
        RECT 25.365 182.175 25.695 182.675 ;
        RECT 25.865 182.345 26.120 182.845 ;
        RECT 27.215 182.345 27.485 183.250 ;
        RECT 27.670 183.105 28.335 183.275 ;
        RECT 27.655 182.175 27.985 182.935 ;
        RECT 28.165 182.345 28.335 183.105 ;
        RECT 28.595 182.175 28.885 183.340 ;
        RECT 29.060 183.315 29.230 183.985 ;
        RECT 29.485 183.815 29.655 183.985 ;
        RECT 29.400 183.485 29.655 183.815 ;
        RECT 29.880 183.485 30.075 183.815 ;
        RECT 29.060 182.345 29.395 183.315 ;
        RECT 29.565 182.175 29.735 183.315 ;
        RECT 29.905 182.515 30.075 183.485 ;
        RECT 30.245 182.855 30.415 183.985 ;
        RECT 30.585 183.195 30.755 183.995 ;
        RECT 30.960 183.705 31.235 184.555 ;
        RECT 30.955 183.535 31.235 183.705 ;
        RECT 30.960 183.395 31.235 183.535 ;
        RECT 31.405 183.195 31.595 184.555 ;
        RECT 31.775 184.190 32.285 184.725 ;
        RECT 32.505 183.915 32.750 184.520 ;
        RECT 33.470 183.915 33.715 184.520 ;
        RECT 33.935 184.190 34.445 184.725 ;
        RECT 31.795 183.745 33.025 183.915 ;
        RECT 30.585 183.025 31.595 183.195 ;
        RECT 31.765 183.180 32.515 183.370 ;
        RECT 30.245 182.685 31.370 182.855 ;
        RECT 31.765 182.515 31.935 183.180 ;
        RECT 32.685 182.935 33.025 183.745 ;
        RECT 29.905 182.345 31.935 182.515 ;
        RECT 32.105 182.175 32.275 182.935 ;
        RECT 32.510 182.525 33.025 182.935 ;
        RECT 33.195 183.745 34.425 183.915 ;
        RECT 33.195 182.935 33.535 183.745 ;
        RECT 33.705 183.180 34.455 183.370 ;
        RECT 33.195 182.525 33.710 182.935 ;
        RECT 33.945 182.175 34.115 182.935 ;
        RECT 34.285 182.515 34.455 183.180 ;
        RECT 34.625 183.195 34.815 184.555 ;
        RECT 34.985 184.385 35.260 184.555 ;
        RECT 34.985 184.215 35.265 184.385 ;
        RECT 34.985 183.395 35.260 184.215 ;
        RECT 35.450 184.190 35.980 184.555 ;
        RECT 36.405 184.325 36.735 184.725 ;
        RECT 35.805 184.155 35.980 184.190 ;
        RECT 35.465 183.195 35.635 183.995 ;
        RECT 34.625 183.025 35.635 183.195 ;
        RECT 35.805 183.985 36.735 184.155 ;
        RECT 36.905 183.985 37.160 184.555 ;
        RECT 35.805 182.855 35.975 183.985 ;
        RECT 36.565 183.815 36.735 183.985 ;
        RECT 34.850 182.685 35.975 182.855 ;
        RECT 36.145 183.485 36.340 183.815 ;
        RECT 36.565 183.485 36.820 183.815 ;
        RECT 36.145 182.515 36.315 183.485 ;
        RECT 36.990 183.315 37.160 183.985 ;
        RECT 37.610 183.915 37.855 184.520 ;
        RECT 38.075 184.190 38.585 184.725 ;
        RECT 34.285 182.345 36.315 182.515 ;
        RECT 36.485 182.175 36.655 183.315 ;
        RECT 36.825 182.345 37.160 183.315 ;
        RECT 37.335 183.745 38.565 183.915 ;
        RECT 37.335 182.935 37.675 183.745 ;
        RECT 37.845 183.180 38.595 183.370 ;
        RECT 37.335 182.525 37.850 182.935 ;
        RECT 38.085 182.175 38.255 182.935 ;
        RECT 38.425 182.515 38.595 183.180 ;
        RECT 38.765 183.195 38.955 184.555 ;
        RECT 39.125 183.705 39.400 184.555 ;
        RECT 39.590 184.190 40.120 184.555 ;
        RECT 40.545 184.325 40.875 184.725 ;
        RECT 39.945 184.155 40.120 184.190 ;
        RECT 39.125 183.535 39.405 183.705 ;
        RECT 39.125 183.395 39.400 183.535 ;
        RECT 39.605 183.195 39.775 183.995 ;
        RECT 38.765 183.025 39.775 183.195 ;
        RECT 39.945 183.985 40.875 184.155 ;
        RECT 41.045 183.985 41.300 184.555 ;
        RECT 39.945 182.855 40.115 183.985 ;
        RECT 40.705 183.815 40.875 183.985 ;
        RECT 38.990 182.685 40.115 182.855 ;
        RECT 40.285 183.485 40.480 183.815 ;
        RECT 40.705 183.485 40.960 183.815 ;
        RECT 40.285 182.515 40.455 183.485 ;
        RECT 41.130 183.315 41.300 183.985 ;
        RECT 41.675 184.095 42.005 184.455 ;
        RECT 42.625 184.265 42.875 184.725 ;
        RECT 43.045 184.265 43.605 184.555 ;
        RECT 41.675 183.905 43.065 184.095 ;
        RECT 42.895 183.815 43.065 183.905 ;
        RECT 38.425 182.345 40.455 182.515 ;
        RECT 40.625 182.175 40.795 183.315 ;
        RECT 40.965 182.345 41.300 183.315 ;
        RECT 41.490 183.485 42.165 183.735 ;
        RECT 42.385 183.485 42.725 183.735 ;
        RECT 42.895 183.485 43.185 183.815 ;
        RECT 41.490 183.125 41.755 183.485 ;
        RECT 42.895 183.235 43.065 183.485 ;
        RECT 42.125 183.065 43.065 183.235 ;
        RECT 41.675 182.175 41.955 182.845 ;
        RECT 42.125 182.515 42.425 183.065 ;
        RECT 43.355 182.895 43.605 184.265 ;
        RECT 43.865 184.075 44.035 184.555 ;
        RECT 44.205 184.245 44.535 184.725 ;
        RECT 44.760 184.305 46.295 184.555 ;
        RECT 44.760 184.075 44.930 184.305 ;
        RECT 43.865 183.905 44.930 184.075 ;
        RECT 45.110 183.735 45.390 184.135 ;
        RECT 43.780 183.525 44.130 183.735 ;
        RECT 44.300 183.535 44.745 183.735 ;
        RECT 44.915 183.535 45.390 183.735 ;
        RECT 45.660 183.735 45.945 184.135 ;
        RECT 46.125 184.075 46.295 184.305 ;
        RECT 46.465 184.245 46.795 184.725 ;
        RECT 47.010 184.225 47.265 184.555 ;
        RECT 47.055 184.215 47.265 184.225 ;
        RECT 47.080 184.145 47.265 184.215 ;
        RECT 46.125 183.905 46.925 184.075 ;
        RECT 45.660 183.535 45.990 183.735 ;
        RECT 46.160 183.705 46.525 183.735 ;
        RECT 46.160 183.535 46.535 183.705 ;
        RECT 46.755 183.355 46.925 183.905 ;
        RECT 42.625 182.175 42.955 182.895 ;
        RECT 43.145 182.345 43.605 182.895 ;
        RECT 43.865 183.185 46.925 183.355 ;
        RECT 43.865 182.345 44.035 183.185 ;
        RECT 47.095 183.015 47.265 184.145 ;
        RECT 47.455 183.905 47.715 184.725 ;
        RECT 47.885 183.905 48.215 184.325 ;
        RECT 48.395 184.240 49.185 184.505 ;
        RECT 47.965 183.815 48.215 183.905 ;
        RECT 44.205 182.515 44.535 183.015 ;
        RECT 44.705 182.775 46.340 183.015 ;
        RECT 44.705 182.685 44.935 182.775 ;
        RECT 45.045 182.515 45.375 182.555 ;
        RECT 44.205 182.345 45.375 182.515 ;
        RECT 45.565 182.175 45.920 182.595 ;
        RECT 46.090 182.345 46.340 182.775 ;
        RECT 46.510 182.175 46.840 182.935 ;
        RECT 47.010 182.345 47.265 183.015 ;
        RECT 47.455 182.855 47.795 183.735 ;
        RECT 47.965 183.565 48.760 183.815 ;
        RECT 47.455 182.175 47.715 182.685 ;
        RECT 47.965 182.345 48.135 183.565 ;
        RECT 48.930 183.385 49.185 184.240 ;
        RECT 49.355 184.085 49.555 184.505 ;
        RECT 49.745 184.265 50.075 184.725 ;
        RECT 49.355 183.565 49.765 184.085 ;
        RECT 50.245 184.075 50.505 184.555 ;
        RECT 49.935 183.385 50.165 183.815 ;
        RECT 48.375 183.215 50.165 183.385 ;
        RECT 48.375 182.850 48.625 183.215 ;
        RECT 48.795 182.855 49.125 183.045 ;
        RECT 49.345 182.920 50.060 183.215 ;
        RECT 50.335 183.045 50.505 184.075 ;
        RECT 48.795 182.680 48.990 182.855 ;
        RECT 48.375 182.175 48.990 182.680 ;
        RECT 49.160 182.345 49.635 182.685 ;
        RECT 49.805 182.175 50.020 182.720 ;
        RECT 50.230 182.345 50.505 183.045 ;
        RECT 50.675 183.985 51.060 184.555 ;
        RECT 51.230 184.265 51.555 184.725 ;
        RECT 52.075 184.095 52.355 184.555 ;
        RECT 50.675 183.315 50.955 183.985 ;
        RECT 51.230 183.925 52.355 184.095 ;
        RECT 51.230 183.815 51.680 183.925 ;
        RECT 51.125 183.485 51.680 183.815 ;
        RECT 52.545 183.755 52.945 184.555 ;
        RECT 53.345 184.265 53.615 184.725 ;
        RECT 53.785 184.095 54.070 184.555 ;
        RECT 50.675 182.345 51.060 183.315 ;
        RECT 51.230 183.025 51.680 183.485 ;
        RECT 51.850 183.195 52.945 183.755 ;
        RECT 51.230 182.805 52.355 183.025 ;
        RECT 51.230 182.175 51.555 182.635 ;
        RECT 52.075 182.345 52.355 182.805 ;
        RECT 52.545 182.345 52.945 183.195 ;
        RECT 53.115 183.925 54.070 184.095 ;
        RECT 54.355 184.000 54.645 184.725 ;
        RECT 55.895 184.165 56.225 184.555 ;
        RECT 56.395 184.335 57.580 184.505 ;
        RECT 57.840 184.255 58.010 184.725 ;
        RECT 55.895 183.985 56.405 184.165 ;
        RECT 53.115 183.025 53.325 183.925 ;
        RECT 53.495 183.195 54.185 183.755 ;
        RECT 55.735 183.525 56.065 183.815 ;
        RECT 56.235 183.355 56.405 183.985 ;
        RECT 56.810 184.075 57.195 184.165 ;
        RECT 58.180 184.075 58.510 184.540 ;
        RECT 56.810 183.905 58.510 184.075 ;
        RECT 58.680 183.905 58.850 184.725 ;
        RECT 59.020 183.905 59.705 184.545 ;
        RECT 61.255 184.345 61.585 184.725 ;
        RECT 60.810 184.175 61.085 184.315 ;
        RECT 61.755 184.175 61.965 184.345 ;
        RECT 60.810 183.985 61.965 184.175 ;
        RECT 62.135 184.175 62.465 184.555 ;
        RECT 62.655 184.345 62.985 184.725 ;
        RECT 62.135 183.970 62.985 184.175 ;
        RECT 56.575 183.525 56.905 183.735 ;
        RECT 57.085 183.485 57.465 183.735 ;
        RECT 57.655 183.705 58.140 183.735 ;
        RECT 57.635 183.535 58.140 183.705 ;
        RECT 53.115 182.805 54.070 183.025 ;
        RECT 53.345 182.175 53.615 182.635 ;
        RECT 53.785 182.345 54.070 182.805 ;
        RECT 54.355 182.175 54.645 183.340 ;
        RECT 55.890 183.185 56.975 183.355 ;
        RECT 55.890 182.345 56.190 183.185 ;
        RECT 56.385 182.175 56.635 183.015 ;
        RECT 56.805 182.935 56.975 183.185 ;
        RECT 57.145 183.105 57.465 183.485 ;
        RECT 57.655 183.525 58.140 183.535 ;
        RECT 58.330 183.525 58.780 183.735 ;
        RECT 58.950 183.525 59.285 183.735 ;
        RECT 57.655 183.105 58.030 183.525 ;
        RECT 58.950 183.355 59.120 183.525 ;
        RECT 58.200 183.185 59.120 183.355 ;
        RECT 58.200 182.935 58.370 183.185 ;
        RECT 56.805 182.765 58.370 182.935 ;
        RECT 57.225 182.345 58.030 182.765 ;
        RECT 58.540 182.175 58.870 183.015 ;
        RECT 59.455 182.935 59.705 183.905 ;
        RECT 60.805 183.360 61.065 183.815 ;
        RECT 61.320 183.410 61.905 183.785 ;
        RECT 59.040 182.345 59.705 182.935 ;
        RECT 60.810 182.175 61.135 183.160 ;
        RECT 61.320 183.025 61.525 183.410 ;
        RECT 62.075 183.195 62.485 183.800 ;
        RECT 62.655 183.480 62.985 183.970 ;
        RECT 62.655 183.025 62.825 183.480 ;
        RECT 61.315 182.855 61.525 183.025 ;
        RECT 61.320 182.825 61.525 182.855 ;
        RECT 61.705 182.805 62.825 183.025 ;
        RECT 61.705 182.345 61.965 182.805 ;
        RECT 62.135 182.175 62.985 182.625 ;
        RECT 63.155 182.345 63.400 184.555 ;
        RECT 63.585 183.925 63.825 184.725 ;
        RECT 64.260 184.365 66.280 184.555 ;
        RECT 66.450 184.365 66.780 184.725 ;
        RECT 67.310 184.365 67.640 184.725 ;
        RECT 68.170 184.365 68.500 184.725 ;
        RECT 69.030 184.365 69.360 184.725 ;
        RECT 66.050 184.195 66.280 184.365 ;
        RECT 70.395 184.345 70.725 184.725 ;
        RECT 70.895 184.195 71.085 184.555 ;
        RECT 71.255 184.365 71.585 184.725 ;
        RECT 71.755 184.195 71.935 184.555 ;
        RECT 72.130 184.365 72.465 184.725 ;
        RECT 72.635 184.195 72.880 184.555 ;
        RECT 73.050 184.365 73.380 184.725 ;
        RECT 73.550 184.195 73.930 184.555 ;
        RECT 74.100 184.365 74.470 184.725 ;
        RECT 75.070 184.195 75.400 184.535 ;
        RECT 64.075 183.965 65.880 184.195 ;
        RECT 66.050 183.990 69.790 184.195 ;
        RECT 70.895 184.175 71.935 184.195 ;
        RECT 64.075 183.365 64.485 183.965 ;
        RECT 69.995 183.935 71.935 184.175 ;
        RECT 72.105 184.005 75.400 184.195 ;
        RECT 75.925 184.005 76.255 184.725 ;
        RECT 76.480 184.365 76.810 184.725 ;
        RECT 76.980 184.195 77.310 184.555 ;
        RECT 77.480 184.285 77.715 184.725 ;
        RECT 78.305 184.345 78.640 184.725 ;
        RECT 79.600 184.385 79.935 184.555 ;
        RECT 76.490 184.025 77.310 184.195 ;
        RECT 64.655 183.535 66.005 183.795 ;
        RECT 63.585 182.175 63.840 183.175 ;
        RECT 64.075 183.110 65.975 183.365 ;
        RECT 66.215 183.295 66.465 183.820 ;
        RECT 66.635 183.465 67.925 183.740 ;
        RECT 68.435 183.490 69.785 183.795 ;
        RECT 68.435 183.295 69.335 183.490 ;
        RECT 66.215 183.125 69.335 183.295 ;
        RECT 69.995 183.315 70.250 183.935 ;
        RECT 72.105 183.765 72.280 184.005 ;
        RECT 70.435 183.485 72.280 183.765 ;
        RECT 72.450 183.485 72.715 183.825 ;
        RECT 72.885 183.535 73.555 183.825 ;
        RECT 73.755 183.705 74.085 183.825 ;
        RECT 73.735 183.535 74.085 183.705 ;
        RECT 64.760 182.955 65.975 183.110 ;
        RECT 69.995 183.105 71.550 183.315 ;
        RECT 72.095 183.305 72.280 183.485 ;
        RECT 72.535 183.365 72.715 183.485 ;
        RECT 73.755 183.365 74.085 183.535 ;
        RECT 72.095 183.135 72.365 183.305 ;
        RECT 64.260 182.175 64.590 182.930 ;
        RECT 64.760 182.785 68.070 182.955 ;
        RECT 64.760 182.725 65.830 182.785 ;
        RECT 64.760 182.345 64.950 182.725 ;
        RECT 65.120 182.175 65.450 182.555 ;
        RECT 65.620 182.345 65.830 182.725 ;
        RECT 68.240 182.725 69.335 182.895 ;
        RECT 66.000 182.175 66.280 182.615 ;
        RECT 68.240 182.535 68.430 182.725 ;
        RECT 66.450 182.345 68.430 182.535 ;
        RECT 68.600 182.175 68.930 182.555 ;
        RECT 69.100 182.345 69.335 182.725 ;
        RECT 69.505 182.175 69.790 182.990 ;
        RECT 70.000 182.175 70.335 182.935 ;
        RECT 70.505 182.345 70.690 183.105 ;
        RECT 70.860 182.175 71.190 182.935 ;
        RECT 71.360 182.345 71.550 183.105 ;
        RECT 71.720 182.175 71.970 182.975 ;
        RECT 72.190 182.940 72.365 183.135 ;
        RECT 72.535 183.110 74.085 183.365 ;
        RECT 74.405 183.300 74.735 183.790 ;
        RECT 74.945 183.480 75.290 183.790 ;
        RECT 75.545 183.490 76.135 183.790 ;
        RECT 75.545 183.300 75.755 183.490 ;
        RECT 74.405 183.110 75.755 183.300 ;
        RECT 72.190 182.770 73.420 182.940 ;
        RECT 75.925 182.930 76.255 183.275 ;
        RECT 74.030 182.705 76.255 182.930 ;
        RECT 76.490 182.905 76.685 184.025 ;
        RECT 77.880 183.985 79.150 184.175 ;
        RECT 79.320 183.985 79.935 184.385 ;
        RECT 80.115 184.000 80.405 184.725 ;
        RECT 76.855 183.485 77.535 183.815 ;
        RECT 77.705 183.485 78.040 183.815 ;
        RECT 78.210 183.705 78.500 183.815 ;
        RECT 78.210 183.535 78.505 183.705 ;
        RECT 78.210 183.485 78.500 183.535 ;
        RECT 78.790 183.485 79.150 183.815 ;
        RECT 77.365 183.300 77.535 183.485 ;
        RECT 79.320 183.300 79.500 183.985 ;
        RECT 80.575 183.925 81.270 184.555 ;
        RECT 81.475 183.925 81.785 184.725 ;
        RECT 82.415 184.250 82.755 184.510 ;
        RECT 79.670 183.485 79.945 183.815 ;
        RECT 80.595 183.485 80.930 183.735 ;
        RECT 77.365 183.045 79.940 183.300 ;
        RECT 76.490 182.735 77.220 182.905 ;
        RECT 74.030 182.600 74.360 182.705 ;
        RECT 72.230 182.345 74.360 182.600 ;
        RECT 74.530 182.175 74.860 182.535 ;
        RECT 75.070 182.345 75.330 182.705 ;
        RECT 75.500 182.175 75.830 182.535 ;
        RECT 76.000 182.345 76.255 182.705 ;
        RECT 76.530 182.175 76.860 182.555 ;
        RECT 77.030 182.345 77.220 182.735 ;
        RECT 77.400 182.175 77.830 182.875 ;
        RECT 78.335 182.345 79.005 183.045 ;
        RECT 79.175 182.175 79.505 182.875 ;
        RECT 79.675 182.345 79.940 183.045 ;
        RECT 80.115 182.175 80.405 183.340 ;
        RECT 81.100 183.325 81.270 183.925 ;
        RECT 81.440 183.485 81.775 183.755 ;
        RECT 80.575 182.175 80.835 183.315 ;
        RECT 81.005 182.345 81.335 183.325 ;
        RECT 81.505 182.175 81.785 183.315 ;
        RECT 82.415 182.645 82.675 184.250 ;
        RECT 82.925 184.245 83.255 184.725 ;
        RECT 83.445 184.075 83.860 184.510 ;
        RECT 84.030 184.210 84.980 184.395 ;
        RECT 82.845 184.000 83.860 184.075 ;
        RECT 82.845 183.905 83.665 184.000 ;
        RECT 82.845 182.985 83.015 183.905 ;
        RECT 83.335 183.175 83.665 183.735 ;
        RECT 83.865 183.485 84.245 183.815 ;
        RECT 84.555 183.485 84.775 184.210 ;
        RECT 85.210 183.815 85.415 184.415 ;
        RECT 85.585 184.000 85.925 184.725 ;
        RECT 86.295 184.095 86.625 184.455 ;
        RECT 87.255 184.265 87.505 184.725 ;
        RECT 87.675 184.265 88.225 184.555 ;
        RECT 86.295 183.905 87.685 184.095 ;
        RECT 87.515 183.815 87.685 183.905 ;
        RECT 83.865 183.365 84.165 183.485 ;
        RECT 83.855 183.195 84.165 183.365 ;
        RECT 83.865 183.190 84.165 183.195 ;
        RECT 85.035 183.185 85.415 183.815 ;
        RECT 85.645 183.185 85.900 183.815 ;
        RECT 86.095 183.485 86.785 183.735 ;
        RECT 87.015 183.485 87.345 183.735 ;
        RECT 87.515 183.485 87.805 183.815 ;
        RECT 86.095 183.045 86.410 183.485 ;
        RECT 87.515 183.235 87.685 183.485 ;
        RECT 86.745 183.065 87.685 183.235 ;
        RECT 82.845 182.815 83.695 182.985 ;
        RECT 82.415 182.385 82.755 182.645 ;
        RECT 82.925 182.175 83.175 182.635 ;
        RECT 83.365 182.385 83.695 182.815 ;
        RECT 83.865 182.845 85.835 183.015 ;
        RECT 83.865 182.345 84.035 182.845 ;
        RECT 84.245 182.175 84.495 182.635 ;
        RECT 84.705 182.345 84.875 182.845 ;
        RECT 85.175 182.175 85.425 182.635 ;
        RECT 85.665 182.345 85.835 182.845 ;
        RECT 86.295 182.175 86.575 182.845 ;
        RECT 86.745 182.515 87.045 183.065 ;
        RECT 87.975 182.895 88.225 184.265 ;
        RECT 88.395 183.925 88.685 184.725 ;
        RECT 89.315 183.925 89.625 184.725 ;
        RECT 89.830 183.925 90.525 184.555 ;
        RECT 90.700 184.250 91.035 184.510 ;
        RECT 91.205 184.325 91.535 184.725 ;
        RECT 91.705 184.325 93.320 184.495 ;
        RECT 89.830 183.875 90.005 183.925 ;
        RECT 89.325 183.485 89.660 183.755 ;
        RECT 89.830 183.325 90.000 183.875 ;
        RECT 90.170 183.485 90.505 183.735 ;
        RECT 87.255 182.175 87.585 182.895 ;
        RECT 87.775 182.345 88.225 182.895 ;
        RECT 88.395 182.175 88.685 183.315 ;
        RECT 89.315 182.175 89.595 183.315 ;
        RECT 89.765 182.345 90.095 183.325 ;
        RECT 90.265 182.175 90.525 183.315 ;
        RECT 90.700 182.895 90.955 184.250 ;
        RECT 91.705 184.155 91.875 184.325 ;
        RECT 91.315 183.985 91.875 184.155 ;
        RECT 92.140 184.045 92.410 184.145 ;
        RECT 91.315 183.815 91.485 183.985 ;
        RECT 92.135 183.875 92.410 184.045 ;
        RECT 91.180 183.485 91.485 183.815 ;
        RECT 91.680 183.705 91.930 183.815 ;
        RECT 91.675 183.535 91.930 183.705 ;
        RECT 91.680 183.485 91.930 183.535 ;
        RECT 92.140 183.485 92.410 183.875 ;
        RECT 92.600 183.705 92.890 184.145 ;
        RECT 92.595 183.535 92.890 183.705 ;
        RECT 92.600 183.485 92.890 183.535 ;
        RECT 93.060 183.485 93.480 184.150 ;
        RECT 93.865 184.005 94.195 184.725 ;
        RECT 95.295 184.105 95.560 184.555 ;
        RECT 95.730 184.275 96.020 184.725 ;
        RECT 96.190 184.105 96.480 184.555 ;
        RECT 95.295 183.935 96.480 184.105 ;
        RECT 96.660 183.815 96.905 184.420 ;
        RECT 93.790 183.485 94.140 183.815 ;
        RECT 91.315 183.315 91.485 183.485 ;
        RECT 93.935 183.365 94.140 183.485 ;
        RECT 91.315 183.145 93.685 183.315 ;
        RECT 93.935 183.195 94.145 183.365 ;
        RECT 95.315 183.150 95.645 183.735 ;
        RECT 95.815 183.485 96.300 183.735 ;
        RECT 96.645 183.485 96.905 183.815 ;
        RECT 97.155 183.485 97.425 184.420 ;
        RECT 97.605 183.735 97.815 184.420 ;
        RECT 97.985 184.075 98.325 184.555 ;
        RECT 98.505 184.245 98.815 184.725 ;
        RECT 97.985 183.905 98.655 184.075 ;
        RECT 98.485 183.815 98.655 183.905 ;
        RECT 97.605 183.485 98.085 183.735 ;
        RECT 98.485 183.485 98.825 183.815 ;
        RECT 90.700 182.385 91.035 182.895 ;
        RECT 91.285 182.175 91.615 182.975 ;
        RECT 91.860 182.765 93.285 182.935 ;
        RECT 91.860 182.345 92.145 182.765 ;
        RECT 92.400 182.175 92.730 182.595 ;
        RECT 92.955 182.515 93.285 182.765 ;
        RECT 93.515 182.685 93.685 183.145 ;
        RECT 93.945 182.515 94.115 183.015 ;
        RECT 92.955 182.345 94.115 182.515 ;
        RECT 95.295 182.175 95.620 182.975 ;
        RECT 95.815 182.395 96.000 183.485 ;
        RECT 98.485 183.315 98.655 183.485 ;
        RECT 96.170 183.145 98.655 183.315 ;
        RECT 96.170 182.345 96.420 183.145 ;
        RECT 96.590 182.175 97.330 182.975 ;
        RECT 97.515 182.345 97.845 183.145 ;
        RECT 98.015 182.175 98.825 182.975 ;
        RECT 98.995 182.345 99.255 184.555 ;
        RECT 99.435 183.955 102.025 184.725 ;
        RECT 102.670 184.155 102.925 184.505 ;
        RECT 103.095 184.325 103.425 184.725 ;
        RECT 103.595 184.155 103.765 184.505 ;
        RECT 103.935 184.325 104.315 184.725 ;
        RECT 102.670 183.985 104.335 184.155 ;
        RECT 104.505 184.050 104.780 184.395 ;
        RECT 99.435 183.435 100.645 183.955 ;
        RECT 104.165 183.815 104.335 183.985 ;
        RECT 100.815 183.265 102.025 183.785 ;
        RECT 102.655 183.485 103.000 183.815 ;
        RECT 103.170 183.485 103.995 183.815 ;
        RECT 104.165 183.485 104.440 183.815 ;
        RECT 99.435 182.175 102.025 183.265 ;
        RECT 102.675 183.025 103.000 183.315 ;
        RECT 103.170 183.195 103.365 183.485 ;
        RECT 104.165 183.315 104.335 183.485 ;
        RECT 104.610 183.315 104.780 184.050 ;
        RECT 105.875 184.000 106.165 184.725 ;
        RECT 107.255 184.250 107.595 184.510 ;
        RECT 103.675 183.145 104.335 183.315 ;
        RECT 103.675 183.025 103.845 183.145 ;
        RECT 102.675 182.855 103.845 183.025 ;
        RECT 102.655 182.395 103.845 182.685 ;
        RECT 104.015 182.175 104.295 182.975 ;
        RECT 104.505 182.345 104.780 183.315 ;
        RECT 105.875 182.175 106.165 183.340 ;
        RECT 107.255 182.645 107.515 184.250 ;
        RECT 107.765 184.245 108.095 184.725 ;
        RECT 108.285 184.075 108.700 184.510 ;
        RECT 108.870 184.210 109.820 184.395 ;
        RECT 107.685 184.000 108.700 184.075 ;
        RECT 107.685 183.905 108.505 184.000 ;
        RECT 107.685 182.985 107.855 183.905 ;
        RECT 108.175 183.175 108.505 183.735 ;
        RECT 108.705 183.485 109.085 183.815 ;
        RECT 109.395 183.485 109.615 184.210 ;
        RECT 110.050 183.815 110.255 184.415 ;
        RECT 110.425 184.000 110.765 184.725 ;
        RECT 110.935 184.180 116.280 184.725 ;
        RECT 108.705 183.365 109.005 183.485 ;
        RECT 108.695 183.195 109.005 183.365 ;
        RECT 108.705 183.190 109.005 183.195 ;
        RECT 109.875 183.185 110.255 183.815 ;
        RECT 110.485 183.185 110.740 183.815 ;
        RECT 112.520 183.350 112.860 184.180 ;
        RECT 116.455 183.955 118.125 184.725 ;
        RECT 118.765 183.985 119.095 184.725 ;
        RECT 119.275 184.195 119.595 184.555 ;
        RECT 119.800 184.365 120.130 184.725 ;
        RECT 120.590 184.195 120.935 184.555 ;
        RECT 119.275 184.025 120.935 184.195 ;
        RECT 107.685 182.815 108.535 182.985 ;
        RECT 107.255 182.385 107.595 182.645 ;
        RECT 107.765 182.175 108.015 182.635 ;
        RECT 108.205 182.385 108.535 182.815 ;
        RECT 108.705 182.845 110.675 183.015 ;
        RECT 108.705 182.345 108.875 182.845 ;
        RECT 109.085 182.175 109.335 182.635 ;
        RECT 109.545 182.345 109.715 182.845 ;
        RECT 110.015 182.175 110.265 182.635 ;
        RECT 110.505 182.345 110.675 182.845 ;
        RECT 114.340 182.610 114.690 183.860 ;
        RECT 116.455 183.435 117.205 183.955 ;
        RECT 117.375 183.265 118.125 183.785 ;
        RECT 110.935 182.175 116.280 182.610 ;
        RECT 116.455 182.175 118.125 183.265 ;
        RECT 118.815 183.185 119.090 183.815 ;
        RECT 118.800 182.525 119.105 183.015 ;
        RECT 119.275 182.695 119.575 184.025 ;
        RECT 121.495 183.945 121.790 184.725 ;
        RECT 122.435 184.245 122.765 184.725 ;
        RECT 119.955 183.565 120.285 183.735 ;
        RECT 119.960 183.315 120.285 183.565 ;
        RECT 120.465 183.485 121.075 183.815 ;
        RECT 121.245 183.315 121.745 183.775 ;
        RECT 122.445 183.485 122.760 184.060 ;
        RECT 122.950 183.485 123.330 184.445 ;
        RECT 123.705 184.155 123.895 184.555 ;
        RECT 124.115 184.365 124.445 184.725 ;
        RECT 124.615 184.175 124.805 184.555 ;
        RECT 124.975 184.345 125.305 184.725 ;
        RECT 123.705 183.985 124.445 184.155 ;
        RECT 124.615 183.985 125.015 184.175 ;
        RECT 125.665 183.995 125.965 184.725 ;
        RECT 124.275 183.815 124.445 183.985 ;
        RECT 123.780 183.400 124.105 183.815 ;
        RECT 119.960 183.135 121.745 183.315 ;
        RECT 119.745 182.785 121.780 182.955 ;
        RECT 119.745 182.525 120.075 182.785 ;
        RECT 120.670 182.705 121.780 182.785 ;
        RECT 118.800 182.345 120.075 182.525 ;
        RECT 120.245 182.175 120.415 182.615 ;
        RECT 120.670 182.345 120.840 182.705 ;
        RECT 121.020 182.175 121.350 182.535 ;
        RECT 121.520 182.345 121.780 182.705 ;
        RECT 122.495 182.875 123.610 183.140 ;
        RECT 124.275 183.120 124.615 183.815 ;
        RECT 122.495 182.345 122.715 182.875 ;
        RECT 122.885 182.175 123.215 182.685 ;
        RECT 123.385 182.345 123.610 182.875 ;
        RECT 123.780 182.890 124.615 183.120 ;
        RECT 123.780 182.345 124.095 182.890 ;
        RECT 124.285 182.175 124.615 182.590 ;
        RECT 124.785 182.345 125.015 183.985 ;
        RECT 126.145 183.815 126.375 184.435 ;
        RECT 126.575 184.165 126.800 184.545 ;
        RECT 126.970 184.335 127.300 184.725 ;
        RECT 126.575 183.985 126.905 184.165 ;
        RECT 125.670 183.485 125.965 183.815 ;
        RECT 126.145 183.485 126.560 183.815 ;
        RECT 126.730 183.315 126.905 183.985 ;
        RECT 127.075 183.485 127.315 184.135 ;
        RECT 127.495 183.955 129.165 184.725 ;
        RECT 129.340 183.995 129.680 184.725 ;
        RECT 127.495 183.435 128.245 183.955 ;
        RECT 125.185 182.175 125.475 183.145 ;
        RECT 125.665 182.955 126.560 183.285 ;
        RECT 126.730 183.125 127.315 183.315 ;
        RECT 128.415 183.265 129.165 183.785 ;
        RECT 129.335 183.485 129.615 183.815 ;
        RECT 129.860 183.705 130.305 184.475 ;
        RECT 130.630 184.095 131.035 184.515 ;
        RECT 131.205 184.245 131.465 184.725 ;
        RECT 130.630 183.985 131.045 184.095 ;
        RECT 131.635 184.000 131.925 184.725 ;
        RECT 129.855 183.535 130.305 183.705 ;
        RECT 130.520 183.365 130.705 183.815 ;
        RECT 125.665 182.785 126.870 182.955 ;
        RECT 125.665 182.355 125.995 182.785 ;
        RECT 126.175 182.175 126.370 182.615 ;
        RECT 126.540 182.355 126.870 182.785 ;
        RECT 127.040 182.355 127.315 183.125 ;
        RECT 127.495 182.175 129.165 183.265 ;
        RECT 129.340 182.175 129.670 183.315 ;
        RECT 130.315 183.195 130.705 183.365 ;
        RECT 130.320 183.145 130.705 183.195 ;
        RECT 130.875 183.315 131.045 183.985 ;
        RECT 131.215 183.485 131.465 183.815 ;
        RECT 133.015 183.780 133.355 184.555 ;
        RECT 133.525 184.265 133.695 184.725 ;
        RECT 133.935 184.290 134.295 184.555 ;
        RECT 133.935 184.285 134.290 184.290 ;
        RECT 133.935 184.275 134.285 184.285 ;
        RECT 133.935 184.270 134.280 184.275 ;
        RECT 133.935 184.260 134.275 184.270 ;
        RECT 134.925 184.265 135.095 184.725 ;
        RECT 133.935 184.255 134.270 184.260 ;
        RECT 133.935 184.245 134.260 184.255 ;
        RECT 133.935 184.235 134.250 184.245 ;
        RECT 133.935 184.095 134.235 184.235 ;
        RECT 133.525 183.905 134.235 184.095 ;
        RECT 134.425 184.095 134.755 184.175 ;
        RECT 135.265 184.095 135.605 184.555 ;
        RECT 134.425 183.905 135.605 184.095 ;
        RECT 135.775 183.975 136.985 184.725 ;
        RECT 130.875 183.145 131.460 183.315 ;
        RECT 129.840 182.805 130.945 182.975 ;
        RECT 129.840 182.395 130.015 182.805 ;
        RECT 130.185 182.175 130.515 182.635 ;
        RECT 130.720 182.395 130.945 182.805 ;
        RECT 131.125 182.365 131.460 183.145 ;
        RECT 131.635 182.175 131.925 183.340 ;
        RECT 133.015 182.345 133.295 183.780 ;
        RECT 133.525 183.335 133.810 183.905 ;
        RECT 133.995 183.505 134.465 183.735 ;
        RECT 134.635 183.715 134.965 183.735 ;
        RECT 134.635 183.535 135.085 183.715 ;
        RECT 135.275 183.535 135.605 183.735 ;
        RECT 133.525 183.120 134.675 183.335 ;
        RECT 133.465 182.175 134.175 182.950 ;
        RECT 134.345 182.345 134.675 183.120 ;
        RECT 134.870 182.420 135.085 183.535 ;
        RECT 135.375 183.195 135.605 183.535 ;
        RECT 135.775 183.435 136.295 183.975 ;
        RECT 136.465 183.265 136.985 183.805 ;
        RECT 135.265 182.175 135.595 182.895 ;
        RECT 135.775 182.175 136.985 183.265 ;
        RECT 137.160 183.125 137.495 184.545 ;
        RECT 137.675 184.355 138.420 184.725 ;
        RECT 138.985 184.185 139.240 184.545 ;
        RECT 139.420 184.355 139.750 184.725 ;
        RECT 139.930 184.185 140.155 184.545 ;
        RECT 137.670 183.995 140.155 184.185 ;
        RECT 137.670 183.305 137.895 183.995 ;
        RECT 140.375 183.955 142.045 184.725 ;
        RECT 142.215 184.095 142.555 184.555 ;
        RECT 142.725 184.265 142.895 184.725 ;
        RECT 143.065 184.345 144.235 184.555 ;
        RECT 143.065 184.095 143.315 184.345 ;
        RECT 143.905 184.325 144.235 184.345 ;
        RECT 138.095 183.485 138.375 183.815 ;
        RECT 138.555 183.485 139.130 183.815 ;
        RECT 139.310 183.485 139.745 183.815 ;
        RECT 139.925 183.485 140.195 183.815 ;
        RECT 140.375 183.435 141.125 183.955 ;
        RECT 142.215 183.925 143.315 184.095 ;
        RECT 143.485 183.905 144.345 184.155 ;
        RECT 137.670 183.125 140.165 183.305 ;
        RECT 141.295 183.265 142.045 183.785 ;
        RECT 142.215 183.485 142.975 183.735 ;
        RECT 143.145 183.485 143.895 183.735 ;
        RECT 144.065 183.315 144.345 183.905 ;
        RECT 144.515 183.955 148.025 184.725 ;
        RECT 144.515 183.435 146.165 183.955 ;
        RECT 148.655 183.925 148.965 184.725 ;
        RECT 149.170 183.925 149.865 184.555 ;
        RECT 150.045 184.000 150.375 184.510 ;
        RECT 150.545 184.325 150.875 184.725 ;
        RECT 151.925 184.155 152.255 184.495 ;
        RECT 152.425 184.325 152.755 184.725 ;
        RECT 153.255 184.225 153.555 184.555 ;
        RECT 153.725 184.245 154.000 184.725 ;
        RECT 137.160 182.355 137.425 183.125 ;
        RECT 137.595 182.175 137.925 182.895 ;
        RECT 138.115 182.715 139.305 182.945 ;
        RECT 138.115 182.355 138.375 182.715 ;
        RECT 138.545 182.175 138.875 182.545 ;
        RECT 139.045 182.355 139.305 182.715 ;
        RECT 139.875 182.355 140.165 183.125 ;
        RECT 140.375 182.175 142.045 183.265 ;
        RECT 142.215 182.175 142.475 183.315 ;
        RECT 142.645 183.145 144.345 183.315 ;
        RECT 146.335 183.265 148.025 183.785 ;
        RECT 148.665 183.485 149.000 183.755 ;
        RECT 149.170 183.325 149.340 183.925 ;
        RECT 149.510 183.485 149.845 183.735 ;
        RECT 142.645 182.345 142.975 183.145 ;
        RECT 143.145 182.175 143.315 182.975 ;
        RECT 143.485 182.345 143.815 183.145 ;
        RECT 143.985 182.175 144.240 182.975 ;
        RECT 144.515 182.175 148.025 183.265 ;
        RECT 148.655 182.175 148.935 183.315 ;
        RECT 149.105 182.345 149.435 183.325 ;
        RECT 149.605 182.175 149.865 183.315 ;
        RECT 150.045 183.235 150.235 184.000 ;
        RECT 150.545 183.985 152.910 184.155 ;
        RECT 150.545 183.815 150.715 183.985 ;
        RECT 150.405 183.485 150.715 183.815 ;
        RECT 150.885 183.485 151.190 183.815 ;
        RECT 150.045 182.385 150.375 183.235 ;
        RECT 150.545 182.175 150.795 183.315 ;
        RECT 150.975 183.155 151.190 183.485 ;
        RECT 151.365 183.155 151.650 183.815 ;
        RECT 151.845 183.155 152.110 183.815 ;
        RECT 152.325 183.155 152.570 183.815 ;
        RECT 152.740 182.985 152.910 183.985 ;
        RECT 150.985 182.815 152.275 182.985 ;
        RECT 150.985 182.395 151.235 182.815 ;
        RECT 151.465 182.175 151.795 182.645 ;
        RECT 152.025 182.395 152.275 182.815 ;
        RECT 152.455 182.815 152.910 182.985 ;
        RECT 153.255 183.315 153.425 184.225 ;
        RECT 154.180 184.075 154.475 184.465 ;
        RECT 154.645 184.245 154.900 184.725 ;
        RECT 155.075 184.075 155.335 184.465 ;
        RECT 155.505 184.245 155.785 184.725 ;
        RECT 153.595 183.485 153.945 184.055 ;
        RECT 154.180 183.905 155.830 184.075 ;
        RECT 156.935 183.975 158.145 184.725 ;
        RECT 154.115 183.565 155.255 183.735 ;
        RECT 154.115 183.315 154.285 183.565 ;
        RECT 155.425 183.395 155.830 183.905 ;
        RECT 153.255 183.145 154.285 183.315 ;
        RECT 155.075 183.225 155.830 183.395 ;
        RECT 156.935 183.265 157.455 183.805 ;
        RECT 157.625 183.435 158.145 183.975 ;
        RECT 152.455 182.385 152.785 182.815 ;
        RECT 153.255 182.345 153.565 183.145 ;
        RECT 155.075 182.975 155.335 183.225 ;
        RECT 153.735 182.175 154.045 182.975 ;
        RECT 154.215 182.805 155.335 182.975 ;
        RECT 154.215 182.345 154.475 182.805 ;
        RECT 154.645 182.175 154.900 182.635 ;
        RECT 155.075 182.345 155.335 182.805 ;
        RECT 155.505 182.175 155.790 183.045 ;
        RECT 156.935 182.175 158.145 183.265 ;
        RECT 2.750 182.005 158.230 182.175 ;
        RECT 2.835 180.915 4.045 182.005 ;
        RECT 4.305 181.335 4.475 181.835 ;
        RECT 4.645 181.505 4.975 182.005 ;
        RECT 4.305 181.165 4.970 181.335 ;
        RECT 2.835 180.205 3.355 180.745 ;
        RECT 3.525 180.375 4.045 180.915 ;
        RECT 4.220 180.345 4.570 180.995 ;
        RECT 2.835 179.455 4.045 180.205 ;
        RECT 4.740 180.175 4.970 181.165 ;
        RECT 4.305 180.005 4.970 180.175 ;
        RECT 4.305 179.715 4.475 180.005 ;
        RECT 4.645 179.455 4.975 179.835 ;
        RECT 5.145 179.715 5.370 181.835 ;
        RECT 5.585 181.505 5.915 182.005 ;
        RECT 6.085 181.335 6.255 181.835 ;
        RECT 6.490 181.620 7.320 181.790 ;
        RECT 7.560 181.625 7.940 182.005 ;
        RECT 5.560 181.165 6.255 181.335 ;
        RECT 5.560 180.195 5.730 181.165 ;
        RECT 5.900 180.375 6.310 180.995 ;
        RECT 6.480 180.945 6.980 181.325 ;
        RECT 5.560 180.005 6.255 180.195 ;
        RECT 6.480 180.075 6.700 180.945 ;
        RECT 7.150 180.775 7.320 181.620 ;
        RECT 8.120 181.455 8.290 181.745 ;
        RECT 8.460 181.625 8.790 182.005 ;
        RECT 9.260 181.535 9.890 181.785 ;
        RECT 10.070 181.625 10.490 182.005 ;
        RECT 9.720 181.455 9.890 181.535 ;
        RECT 10.690 181.455 10.930 181.745 ;
        RECT 7.490 181.205 8.860 181.455 ;
        RECT 7.490 180.945 7.740 181.205 ;
        RECT 8.250 180.775 8.500 180.935 ;
        RECT 7.150 180.605 8.500 180.775 ;
        RECT 7.150 180.565 7.570 180.605 ;
        RECT 6.880 180.015 7.230 180.385 ;
        RECT 5.585 179.455 5.915 179.835 ;
        RECT 6.085 179.675 6.255 180.005 ;
        RECT 7.400 179.835 7.570 180.565 ;
        RECT 8.670 180.435 8.860 181.205 ;
        RECT 7.740 180.105 8.150 180.435 ;
        RECT 8.440 180.095 8.860 180.435 ;
        RECT 9.030 181.025 9.550 181.335 ;
        RECT 9.720 181.285 10.930 181.455 ;
        RECT 11.160 181.315 11.490 182.005 ;
        RECT 9.030 180.265 9.200 181.025 ;
        RECT 9.370 180.435 9.550 180.845 ;
        RECT 9.720 180.775 9.890 181.285 ;
        RECT 11.660 181.135 11.830 181.745 ;
        RECT 12.100 181.285 12.430 181.795 ;
        RECT 11.660 181.115 11.980 181.135 ;
        RECT 10.060 180.945 11.980 181.115 ;
        RECT 9.720 180.605 11.620 180.775 ;
        RECT 9.950 180.265 10.280 180.385 ;
        RECT 9.030 180.095 10.280 180.265 ;
        RECT 6.555 179.635 7.570 179.835 ;
        RECT 7.740 179.455 8.150 179.895 ;
        RECT 8.440 179.665 8.690 180.095 ;
        RECT 8.890 179.455 9.210 179.915 ;
        RECT 10.450 179.845 10.620 180.605 ;
        RECT 11.290 180.545 11.620 180.605 ;
        RECT 10.810 180.375 11.140 180.435 ;
        RECT 10.810 180.105 11.470 180.375 ;
        RECT 11.790 180.050 11.980 180.945 ;
        RECT 9.770 179.675 10.620 179.845 ;
        RECT 10.820 179.455 11.480 179.935 ;
        RECT 11.660 179.720 11.980 180.050 ;
        RECT 12.180 180.695 12.430 181.285 ;
        RECT 12.610 181.205 12.895 182.005 ;
        RECT 13.075 181.025 13.330 181.695 ;
        RECT 12.180 180.365 12.980 180.695 ;
        RECT 12.180 179.715 12.430 180.365 ;
        RECT 13.150 180.165 13.330 181.025 ;
        RECT 14.425 181.075 14.595 181.835 ;
        RECT 14.775 181.245 15.105 182.005 ;
        RECT 14.425 180.905 15.090 181.075 ;
        RECT 15.275 180.930 15.545 181.835 ;
        RECT 14.920 180.760 15.090 180.905 ;
        RECT 14.355 180.355 14.685 180.725 ;
        RECT 14.920 180.430 15.205 180.760 ;
        RECT 14.920 180.175 15.090 180.430 ;
        RECT 13.075 179.965 13.330 180.165 ;
        RECT 14.425 180.005 15.090 180.175 ;
        RECT 15.375 180.130 15.545 180.930 ;
        RECT 15.715 180.840 16.005 182.005 ;
        RECT 16.550 181.665 16.805 181.695 ;
        RECT 16.465 181.495 16.805 181.665 ;
        RECT 16.550 181.025 16.805 181.495 ;
        RECT 16.985 181.205 17.270 182.005 ;
        RECT 17.450 181.285 17.780 181.795 ;
        RECT 12.610 179.455 12.895 179.915 ;
        RECT 13.075 179.795 13.415 179.965 ;
        RECT 13.075 179.635 13.330 179.795 ;
        RECT 14.425 179.625 14.595 180.005 ;
        RECT 14.775 179.455 15.105 179.835 ;
        RECT 15.285 179.625 15.545 180.130 ;
        RECT 15.715 179.455 16.005 180.180 ;
        RECT 16.550 180.165 16.730 181.025 ;
        RECT 17.450 180.695 17.700 181.285 ;
        RECT 18.050 181.135 18.220 181.745 ;
        RECT 18.390 181.315 18.720 182.005 ;
        RECT 18.950 181.455 19.190 181.745 ;
        RECT 19.390 181.625 19.810 182.005 ;
        RECT 19.990 181.535 20.620 181.785 ;
        RECT 21.090 181.625 21.420 182.005 ;
        RECT 19.990 181.455 20.160 181.535 ;
        RECT 21.590 181.455 21.760 181.745 ;
        RECT 21.940 181.625 22.320 182.005 ;
        RECT 22.560 181.620 23.390 181.790 ;
        RECT 18.950 181.285 20.160 181.455 ;
        RECT 16.900 180.365 17.700 180.695 ;
        RECT 16.550 179.635 16.805 180.165 ;
        RECT 16.985 179.455 17.270 179.915 ;
        RECT 17.450 179.715 17.700 180.365 ;
        RECT 17.900 181.115 18.220 181.135 ;
        RECT 17.900 180.945 19.820 181.115 ;
        RECT 17.900 180.050 18.090 180.945 ;
        RECT 19.990 180.775 20.160 181.285 ;
        RECT 20.330 181.025 20.850 181.335 ;
        RECT 18.260 180.605 20.160 180.775 ;
        RECT 18.260 180.545 18.590 180.605 ;
        RECT 18.740 180.375 19.070 180.435 ;
        RECT 18.410 180.105 19.070 180.375 ;
        RECT 17.900 179.720 18.220 180.050 ;
        RECT 18.400 179.455 19.060 179.935 ;
        RECT 19.260 179.845 19.430 180.605 ;
        RECT 20.330 180.435 20.510 180.845 ;
        RECT 19.600 180.265 19.930 180.385 ;
        RECT 20.680 180.265 20.850 181.025 ;
        RECT 19.600 180.095 20.850 180.265 ;
        RECT 21.020 181.205 22.390 181.455 ;
        RECT 21.020 180.435 21.210 181.205 ;
        RECT 22.140 180.945 22.390 181.205 ;
        RECT 21.380 180.775 21.630 180.935 ;
        RECT 22.560 180.775 22.730 181.620 ;
        RECT 23.625 181.335 23.795 181.835 ;
        RECT 23.965 181.505 24.295 182.005 ;
        RECT 22.900 180.945 23.400 181.325 ;
        RECT 23.625 181.165 24.320 181.335 ;
        RECT 21.380 180.605 22.730 180.775 ;
        RECT 22.310 180.565 22.730 180.605 ;
        RECT 21.020 180.095 21.440 180.435 ;
        RECT 21.730 180.105 22.140 180.435 ;
        RECT 19.260 179.675 20.110 179.845 ;
        RECT 20.670 179.455 20.990 179.915 ;
        RECT 21.190 179.665 21.440 180.095 ;
        RECT 21.730 179.455 22.140 179.895 ;
        RECT 22.310 179.835 22.480 180.565 ;
        RECT 22.650 180.015 23.000 180.385 ;
        RECT 23.180 180.075 23.400 180.945 ;
        RECT 23.570 180.375 23.980 180.995 ;
        RECT 24.150 180.195 24.320 181.165 ;
        RECT 23.625 180.005 24.320 180.195 ;
        RECT 22.310 179.635 23.325 179.835 ;
        RECT 23.625 179.675 23.795 180.005 ;
        RECT 23.965 179.455 24.295 179.835 ;
        RECT 24.510 179.715 24.735 181.835 ;
        RECT 24.905 181.505 25.235 182.005 ;
        RECT 25.405 181.335 25.575 181.835 ;
        RECT 24.910 181.165 25.575 181.335 ;
        RECT 24.910 180.175 25.140 181.165 ;
        RECT 25.310 180.345 25.660 180.995 ;
        RECT 25.835 180.930 26.105 181.835 ;
        RECT 26.275 181.245 26.605 182.005 ;
        RECT 26.785 181.075 26.955 181.835 ;
        RECT 27.680 181.335 27.935 181.835 ;
        RECT 28.105 181.505 28.435 182.005 ;
        RECT 27.680 181.165 28.430 181.335 ;
        RECT 24.910 180.005 25.575 180.175 ;
        RECT 24.905 179.455 25.235 179.835 ;
        RECT 25.405 179.715 25.575 180.005 ;
        RECT 25.835 180.130 26.005 180.930 ;
        RECT 26.290 180.905 26.955 181.075 ;
        RECT 26.290 180.760 26.460 180.905 ;
        RECT 26.175 180.430 26.460 180.760 ;
        RECT 26.290 180.175 26.460 180.430 ;
        RECT 26.695 180.355 27.025 180.725 ;
        RECT 27.680 180.345 28.030 180.995 ;
        RECT 28.200 180.175 28.430 181.165 ;
        RECT 25.835 179.625 26.095 180.130 ;
        RECT 26.290 180.005 26.955 180.175 ;
        RECT 26.275 179.455 26.605 179.835 ;
        RECT 26.785 179.625 26.955 180.005 ;
        RECT 27.680 180.005 28.430 180.175 ;
        RECT 27.680 179.715 27.935 180.005 ;
        RECT 28.105 179.455 28.435 179.835 ;
        RECT 28.605 179.715 28.775 181.835 ;
        RECT 28.945 181.035 29.270 181.820 ;
        RECT 29.440 181.545 29.690 182.005 ;
        RECT 29.860 181.505 30.110 181.835 ;
        RECT 30.325 181.505 31.005 181.835 ;
        RECT 29.860 181.375 30.030 181.505 ;
        RECT 29.635 181.205 30.030 181.375 ;
        RECT 29.005 179.985 29.465 181.035 ;
        RECT 29.635 179.845 29.805 181.205 ;
        RECT 30.200 180.945 30.665 181.335 ;
        RECT 29.975 180.135 30.325 180.755 ;
        RECT 30.495 180.355 30.665 180.945 ;
        RECT 30.835 180.725 31.005 181.505 ;
        RECT 31.175 181.405 31.345 181.745 ;
        RECT 31.580 181.575 31.910 182.005 ;
        RECT 32.080 181.405 32.250 181.745 ;
        RECT 32.545 181.545 32.915 182.005 ;
        RECT 31.175 181.235 32.250 181.405 ;
        RECT 33.085 181.375 33.255 181.835 ;
        RECT 33.490 181.495 34.360 181.835 ;
        RECT 34.530 181.545 34.780 182.005 ;
        RECT 32.695 181.205 33.255 181.375 ;
        RECT 32.695 181.065 32.865 181.205 ;
        RECT 31.365 180.895 32.865 181.065 ;
        RECT 33.560 181.035 34.020 181.325 ;
        RECT 30.835 180.555 32.525 180.725 ;
        RECT 30.495 180.135 30.850 180.355 ;
        RECT 31.020 179.845 31.190 180.555 ;
        RECT 31.395 180.135 32.185 180.385 ;
        RECT 32.355 180.375 32.525 180.555 ;
        RECT 32.695 180.205 32.865 180.895 ;
        RECT 29.135 179.455 29.465 179.815 ;
        RECT 29.635 179.675 30.130 179.845 ;
        RECT 30.335 179.675 31.190 179.845 ;
        RECT 32.065 179.455 32.395 179.915 ;
        RECT 32.605 179.815 32.865 180.205 ;
        RECT 33.055 181.025 34.020 181.035 ;
        RECT 34.190 181.115 34.360 181.495 ;
        RECT 34.950 181.455 35.120 181.745 ;
        RECT 35.300 181.625 35.630 182.005 ;
        RECT 34.950 181.285 35.750 181.455 ;
        RECT 33.055 180.865 33.730 181.025 ;
        RECT 34.190 180.945 35.410 181.115 ;
        RECT 33.055 180.075 33.265 180.865 ;
        RECT 34.190 180.855 34.360 180.945 ;
        RECT 33.435 180.075 33.785 180.695 ;
        RECT 33.955 180.685 34.360 180.855 ;
        RECT 33.955 179.905 34.125 180.685 ;
        RECT 34.295 180.235 34.515 180.515 ;
        RECT 34.695 180.405 35.235 180.775 ;
        RECT 35.580 180.695 35.750 181.285 ;
        RECT 35.970 180.865 36.275 182.005 ;
        RECT 36.445 180.815 36.700 181.695 ;
        RECT 35.580 180.665 36.320 180.695 ;
        RECT 34.295 180.065 34.825 180.235 ;
        RECT 32.605 179.645 32.955 179.815 ;
        RECT 33.175 179.625 34.125 179.905 ;
        RECT 34.295 179.455 34.485 179.895 ;
        RECT 34.655 179.835 34.825 180.065 ;
        RECT 34.995 180.005 35.235 180.405 ;
        RECT 35.405 180.365 36.320 180.665 ;
        RECT 35.405 180.190 35.730 180.365 ;
        RECT 35.405 179.835 35.725 180.190 ;
        RECT 36.490 180.165 36.700 180.815 ;
        RECT 34.655 179.665 35.725 179.835 ;
        RECT 35.970 179.455 36.275 179.915 ;
        RECT 36.445 179.635 36.700 180.165 ;
        RECT 36.880 180.865 37.215 181.835 ;
        RECT 37.385 180.865 37.555 182.005 ;
        RECT 37.725 181.665 39.755 181.835 ;
        RECT 36.880 180.195 37.050 180.865 ;
        RECT 37.725 180.695 37.895 181.665 ;
        RECT 37.220 180.365 37.475 180.695 ;
        RECT 37.700 180.365 37.895 180.695 ;
        RECT 38.065 181.325 39.190 181.495 ;
        RECT 37.305 180.195 37.475 180.365 ;
        RECT 38.065 180.195 38.235 181.325 ;
        RECT 36.880 179.625 37.135 180.195 ;
        RECT 37.305 180.025 38.235 180.195 ;
        RECT 38.405 180.985 39.415 181.155 ;
        RECT 38.405 180.185 38.575 180.985 ;
        RECT 38.060 179.990 38.235 180.025 ;
        RECT 37.305 179.455 37.635 179.855 ;
        RECT 38.060 179.625 38.590 179.990 ;
        RECT 38.780 179.965 39.055 180.785 ;
        RECT 38.775 179.795 39.055 179.965 ;
        RECT 38.780 179.625 39.055 179.795 ;
        RECT 39.225 179.625 39.415 180.985 ;
        RECT 39.585 181.000 39.755 181.665 ;
        RECT 39.925 181.245 40.095 182.005 ;
        RECT 40.330 181.245 40.845 181.655 ;
        RECT 39.585 180.810 40.335 181.000 ;
        RECT 40.505 180.435 40.845 181.245 ;
        RECT 41.475 180.840 41.765 182.005 ;
        RECT 41.985 180.910 42.235 182.005 ;
        RECT 42.970 181.665 45.035 181.835 ;
        RECT 42.405 180.825 42.760 181.240 ;
        RECT 42.970 180.825 43.215 181.665 ;
        RECT 42.590 180.655 42.760 180.825 ;
        RECT 41.935 180.445 42.420 180.655 ;
        RECT 42.590 180.445 43.215 180.655 ;
        RECT 39.615 180.265 40.845 180.435 ;
        RECT 42.590 180.275 42.760 180.445 ;
        RECT 43.385 180.305 43.635 181.495 ;
        RECT 43.805 180.825 44.075 181.665 ;
        RECT 44.365 180.995 44.615 181.495 ;
        RECT 44.785 181.165 45.035 181.665 ;
        RECT 45.205 180.995 45.455 181.835 ;
        RECT 45.625 181.165 45.875 182.005 ;
        RECT 46.045 180.995 46.360 181.835 ;
        RECT 44.365 180.825 46.360 180.995 ;
        RECT 46.720 181.035 47.110 181.210 ;
        RECT 47.595 181.205 47.925 182.005 ;
        RECT 48.095 181.215 48.630 181.835 ;
        RECT 46.720 180.865 48.145 181.035 ;
        RECT 43.810 180.445 45.315 180.655 ;
        RECT 45.485 180.445 46.340 180.655 ;
        RECT 43.375 180.275 43.635 180.305 ;
        RECT 39.595 179.455 40.105 179.990 ;
        RECT 40.325 179.660 40.570 180.265 ;
        RECT 41.475 179.455 41.765 180.180 ;
        RECT 41.945 179.455 42.235 180.195 ;
        RECT 42.405 179.750 42.760 180.275 ;
        RECT 42.970 179.455 43.175 180.265 ;
        RECT 43.345 180.095 45.915 180.275 ;
        RECT 43.345 179.625 43.675 180.095 ;
        RECT 43.845 179.455 44.575 179.925 ;
        RECT 44.745 179.625 45.075 180.095 ;
        RECT 45.245 179.455 45.415 179.925 ;
        RECT 45.585 179.625 45.915 180.095 ;
        RECT 46.085 179.455 46.360 180.275 ;
        RECT 46.595 180.135 46.950 180.695 ;
        RECT 47.120 179.965 47.290 180.865 ;
        RECT 47.460 180.135 47.725 180.695 ;
        RECT 47.975 180.365 48.145 180.865 ;
        RECT 48.315 180.195 48.630 181.215 ;
        RECT 48.925 180.995 49.095 181.835 ;
        RECT 49.265 181.665 50.435 181.835 ;
        RECT 49.265 181.165 49.595 181.665 ;
        RECT 50.105 181.625 50.435 181.665 ;
        RECT 50.625 181.585 50.980 182.005 ;
        RECT 49.765 181.405 49.995 181.495 ;
        RECT 51.150 181.405 51.400 181.835 ;
        RECT 49.765 181.165 51.400 181.405 ;
        RECT 51.570 181.245 51.900 182.005 ;
        RECT 52.070 181.165 52.325 181.835 ;
        RECT 48.925 180.825 51.985 180.995 ;
        RECT 48.840 180.445 49.190 180.655 ;
        RECT 49.360 180.445 49.805 180.645 ;
        RECT 49.975 180.445 50.450 180.645 ;
        RECT 46.700 179.455 46.940 179.965 ;
        RECT 47.120 179.635 47.400 179.965 ;
        RECT 47.630 179.455 47.845 179.965 ;
        RECT 48.015 179.625 48.630 180.195 ;
        RECT 48.925 180.105 49.990 180.275 ;
        RECT 48.925 179.625 49.095 180.105 ;
        RECT 49.265 179.455 49.595 179.935 ;
        RECT 49.820 179.875 49.990 180.105 ;
        RECT 50.170 180.045 50.450 180.445 ;
        RECT 50.720 180.445 51.050 180.645 ;
        RECT 51.220 180.475 51.595 180.645 ;
        RECT 51.220 180.445 51.585 180.475 ;
        RECT 50.720 180.045 51.005 180.445 ;
        RECT 51.815 180.275 51.985 180.825 ;
        RECT 51.185 180.105 51.985 180.275 ;
        RECT 51.185 179.875 51.355 180.105 ;
        RECT 52.155 180.035 52.325 181.165 ;
        RECT 52.140 179.955 52.325 180.035 ;
        RECT 49.820 179.625 51.355 179.875 ;
        RECT 51.525 179.455 51.855 179.935 ;
        RECT 52.070 179.625 52.325 179.955 ;
        RECT 52.525 179.635 52.785 181.825 ;
        RECT 52.955 181.275 53.295 182.005 ;
        RECT 53.475 181.095 53.745 181.825 ;
        RECT 52.975 180.875 53.745 181.095 ;
        RECT 53.925 181.115 54.155 181.825 ;
        RECT 54.325 181.295 54.655 182.005 ;
        RECT 54.825 181.115 55.085 181.825 ;
        RECT 56.200 181.335 56.455 181.835 ;
        RECT 56.625 181.505 56.955 182.005 ;
        RECT 56.200 181.165 56.950 181.335 ;
        RECT 53.925 180.875 55.085 181.115 ;
        RECT 52.975 180.205 53.265 180.875 ;
        RECT 53.445 180.385 53.910 180.695 ;
        RECT 54.090 180.385 54.615 180.695 ;
        RECT 52.975 180.005 54.205 180.205 ;
        RECT 53.045 179.455 53.715 179.825 ;
        RECT 53.895 179.635 54.205 180.005 ;
        RECT 54.385 179.745 54.615 180.385 ;
        RECT 54.795 180.365 55.095 180.695 ;
        RECT 56.200 180.345 56.550 180.995 ;
        RECT 54.795 179.455 55.085 180.185 ;
        RECT 56.720 180.175 56.950 181.165 ;
        RECT 56.200 180.005 56.950 180.175 ;
        RECT 56.200 179.715 56.455 180.005 ;
        RECT 56.625 179.455 56.955 179.835 ;
        RECT 57.125 179.715 57.295 181.835 ;
        RECT 57.465 181.035 57.790 181.820 ;
        RECT 57.960 181.545 58.210 182.005 ;
        RECT 58.380 181.505 58.630 181.835 ;
        RECT 58.845 181.505 59.525 181.835 ;
        RECT 58.380 181.375 58.550 181.505 ;
        RECT 58.155 181.205 58.550 181.375 ;
        RECT 57.525 179.985 57.985 181.035 ;
        RECT 58.155 179.845 58.325 181.205 ;
        RECT 58.720 180.945 59.185 181.335 ;
        RECT 58.495 180.135 58.845 180.755 ;
        RECT 59.015 180.355 59.185 180.945 ;
        RECT 59.355 180.725 59.525 181.505 ;
        RECT 59.695 181.405 59.865 181.745 ;
        RECT 60.100 181.575 60.430 182.005 ;
        RECT 60.600 181.405 60.770 181.745 ;
        RECT 61.065 181.545 61.435 182.005 ;
        RECT 59.695 181.235 60.770 181.405 ;
        RECT 61.605 181.375 61.775 181.835 ;
        RECT 62.010 181.495 62.880 181.835 ;
        RECT 63.050 181.545 63.300 182.005 ;
        RECT 61.215 181.205 61.775 181.375 ;
        RECT 61.215 181.065 61.385 181.205 ;
        RECT 59.885 180.895 61.385 181.065 ;
        RECT 62.080 181.035 62.540 181.325 ;
        RECT 59.355 180.555 61.045 180.725 ;
        RECT 59.015 180.135 59.370 180.355 ;
        RECT 59.540 179.845 59.710 180.555 ;
        RECT 59.915 180.135 60.705 180.385 ;
        RECT 60.875 180.375 61.045 180.555 ;
        RECT 61.215 180.205 61.385 180.895 ;
        RECT 57.655 179.455 57.985 179.815 ;
        RECT 58.155 179.675 58.650 179.845 ;
        RECT 58.855 179.675 59.710 179.845 ;
        RECT 60.585 179.455 60.915 179.915 ;
        RECT 61.125 179.815 61.385 180.205 ;
        RECT 61.575 181.025 62.540 181.035 ;
        RECT 62.710 181.115 62.880 181.495 ;
        RECT 63.470 181.455 63.640 181.745 ;
        RECT 63.820 181.625 64.150 182.005 ;
        RECT 63.470 181.285 64.270 181.455 ;
        RECT 61.575 180.865 62.250 181.025 ;
        RECT 62.710 180.945 63.930 181.115 ;
        RECT 61.575 180.075 61.785 180.865 ;
        RECT 62.710 180.855 62.880 180.945 ;
        RECT 61.955 180.075 62.305 180.695 ;
        RECT 62.475 180.685 62.880 180.855 ;
        RECT 62.475 179.905 62.645 180.685 ;
        RECT 62.815 180.235 63.035 180.515 ;
        RECT 63.215 180.405 63.755 180.775 ;
        RECT 64.100 180.665 64.270 181.285 ;
        RECT 64.445 180.945 64.615 182.005 ;
        RECT 64.825 180.995 65.115 181.835 ;
        RECT 65.285 181.165 65.455 182.005 ;
        RECT 65.665 180.995 65.915 181.835 ;
        RECT 66.125 181.165 66.295 182.005 ;
        RECT 64.825 180.825 66.550 180.995 ;
        RECT 67.235 180.840 67.525 182.005 ;
        RECT 67.700 181.495 69.355 181.785 ;
        RECT 67.700 181.155 69.290 181.325 ;
        RECT 69.525 181.205 69.805 182.005 ;
        RECT 67.700 180.865 68.020 181.155 ;
        RECT 69.120 181.035 69.290 181.155 ;
        RECT 62.815 180.065 63.345 180.235 ;
        RECT 61.125 179.645 61.475 179.815 ;
        RECT 61.695 179.625 62.645 179.905 ;
        RECT 62.815 179.455 63.005 179.895 ;
        RECT 63.175 179.835 63.345 180.065 ;
        RECT 63.515 180.005 63.755 180.405 ;
        RECT 63.925 180.655 64.270 180.665 ;
        RECT 63.925 180.445 65.955 180.655 ;
        RECT 63.925 180.190 64.250 180.445 ;
        RECT 66.140 180.275 66.550 180.825 ;
        RECT 63.925 179.835 64.245 180.190 ;
        RECT 63.175 179.665 64.245 179.835 ;
        RECT 64.445 179.455 64.615 180.265 ;
        RECT 64.785 180.105 66.550 180.275 ;
        RECT 64.785 179.625 65.115 180.105 ;
        RECT 65.285 179.455 65.455 179.925 ;
        RECT 65.625 179.625 65.955 180.105 ;
        RECT 66.125 179.455 66.295 179.925 ;
        RECT 67.235 179.455 67.525 180.180 ;
        RECT 67.700 180.125 68.050 180.695 ;
        RECT 68.220 180.365 68.930 180.985 ;
        RECT 69.120 180.865 69.845 181.035 ;
        RECT 70.015 180.865 70.285 181.835 ;
        RECT 69.675 180.695 69.845 180.865 ;
        RECT 69.100 180.365 69.505 180.695 ;
        RECT 69.675 180.365 69.945 180.695 ;
        RECT 69.675 180.195 69.845 180.365 ;
        RECT 68.235 180.025 69.845 180.195 ;
        RECT 70.115 180.130 70.285 180.865 ;
        RECT 70.480 180.780 70.735 182.005 ;
        RECT 70.905 181.165 71.160 181.835 ;
        RECT 71.330 181.605 71.660 182.005 ;
        RECT 72.530 181.605 72.935 182.005 ;
        RECT 73.205 181.425 73.555 181.795 ;
        RECT 71.470 181.255 73.555 181.425 ;
        RECT 67.705 179.455 68.035 179.955 ;
        RECT 68.235 179.675 68.405 180.025 ;
        RECT 68.605 179.455 68.935 179.855 ;
        RECT 69.105 179.675 69.275 180.025 ;
        RECT 69.445 179.455 69.825 179.855 ;
        RECT 70.015 179.785 70.285 180.130 ;
        RECT 70.480 179.455 70.735 180.280 ;
        RECT 70.905 180.195 71.075 181.165 ;
        RECT 71.470 180.985 71.640 181.255 ;
        RECT 71.245 180.815 71.640 180.985 ;
        RECT 71.810 180.865 72.830 181.085 ;
        RECT 71.245 180.365 71.415 180.815 ;
        RECT 72.565 180.725 72.830 180.865 ;
        RECT 73.000 180.865 73.555 181.255 ;
        RECT 73.725 181.665 73.895 181.795 ;
        RECT 73.725 181.495 73.905 181.665 ;
        RECT 71.585 180.445 72.055 180.645 ;
        RECT 72.225 180.275 72.395 180.470 ;
        RECT 70.905 179.625 71.240 180.195 ;
        RECT 71.885 180.140 72.395 180.275 ;
        RECT 71.435 179.455 71.605 180.120 ;
        RECT 71.885 180.105 72.390 180.140 ;
        RECT 71.885 179.750 72.105 180.105 ;
        RECT 72.565 179.935 72.735 180.725 ;
        RECT 73.000 180.615 73.170 180.865 ;
        RECT 73.725 180.695 73.895 181.495 ;
        RECT 74.100 181.185 74.415 182.005 ;
        RECT 72.980 180.445 73.170 180.615 ;
        RECT 73.340 180.445 73.895 180.695 ;
        RECT 74.070 180.445 74.415 181.015 ;
        RECT 74.595 180.915 75.805 182.005 ;
        RECT 76.065 181.260 76.335 182.005 ;
        RECT 76.965 182.000 83.240 182.005 ;
        RECT 76.505 181.090 76.795 181.830 ;
        RECT 76.965 181.275 77.220 182.000 ;
        RECT 77.405 181.105 77.665 181.830 ;
        RECT 77.835 181.275 78.080 182.000 ;
        RECT 78.265 181.105 78.525 181.830 ;
        RECT 78.695 181.275 78.940 182.000 ;
        RECT 79.125 181.105 79.385 181.830 ;
        RECT 79.555 181.275 79.800 182.000 ;
        RECT 79.970 181.105 80.230 181.830 ;
        RECT 80.400 181.275 80.660 182.000 ;
        RECT 80.830 181.105 81.090 181.830 ;
        RECT 81.260 181.275 81.520 182.000 ;
        RECT 81.690 181.105 81.950 181.830 ;
        RECT 82.120 181.275 82.380 182.000 ;
        RECT 82.550 181.105 82.810 181.830 ;
        RECT 82.980 181.205 83.240 182.000 ;
        RECT 77.405 181.090 82.810 181.105 ;
        RECT 72.980 180.060 73.150 180.445 ;
        RECT 72.275 179.765 72.735 179.935 ;
        RECT 72.905 179.690 73.150 180.060 ;
        RECT 73.325 180.095 74.415 180.275 ;
        RECT 73.325 179.690 73.555 180.095 ;
        RECT 73.745 179.455 73.915 179.925 ;
        RECT 74.085 179.690 74.415 180.095 ;
        RECT 74.595 180.205 75.115 180.745 ;
        RECT 75.285 180.375 75.805 180.915 ;
        RECT 76.065 180.865 82.810 181.090 ;
        RECT 76.065 180.275 77.230 180.865 ;
        RECT 83.410 180.695 83.660 181.830 ;
        RECT 83.840 181.195 84.100 182.005 ;
        RECT 84.275 180.695 84.520 181.835 ;
        RECT 84.700 181.195 84.995 182.005 ;
        RECT 85.180 181.035 85.455 181.835 ;
        RECT 85.625 181.205 85.955 182.005 ;
        RECT 86.125 181.035 86.295 181.835 ;
        RECT 86.465 181.205 86.715 182.005 ;
        RECT 86.885 181.665 88.980 181.835 ;
        RECT 86.885 181.035 87.215 181.665 ;
        RECT 85.180 180.825 87.215 181.035 ;
        RECT 87.385 181.115 87.555 181.495 ;
        RECT 87.725 181.305 88.055 181.665 ;
        RECT 88.225 181.115 88.395 181.495 ;
        RECT 88.565 181.285 88.980 181.665 ;
        RECT 89.370 181.135 89.655 182.005 ;
        RECT 89.825 181.375 90.085 181.835 ;
        RECT 90.260 181.545 90.515 182.005 ;
        RECT 90.685 181.375 90.945 181.835 ;
        RECT 89.825 181.205 90.945 181.375 ;
        RECT 91.115 181.205 91.425 182.005 ;
        RECT 87.385 180.815 89.145 181.115 ;
        RECT 89.825 180.955 90.085 181.205 ;
        RECT 91.595 181.035 91.905 181.835 ;
        RECT 77.400 180.445 84.520 180.695 ;
        RECT 74.595 179.455 75.805 180.205 ;
        RECT 76.065 180.105 82.810 180.275 ;
        RECT 76.065 179.455 76.365 179.935 ;
        RECT 76.535 179.650 76.795 180.105 ;
        RECT 76.965 179.455 77.225 179.935 ;
        RECT 77.405 179.650 77.665 180.105 ;
        RECT 77.835 179.455 78.085 179.935 ;
        RECT 78.265 179.650 78.525 180.105 ;
        RECT 78.695 179.455 78.945 179.935 ;
        RECT 79.125 179.650 79.385 180.105 ;
        RECT 79.555 179.455 79.800 179.935 ;
        RECT 79.970 179.650 80.245 180.105 ;
        RECT 80.415 179.455 80.660 179.935 ;
        RECT 80.830 179.650 81.090 180.105 ;
        RECT 81.260 179.455 81.520 179.935 ;
        RECT 81.690 179.650 81.950 180.105 ;
        RECT 82.120 179.455 82.380 179.935 ;
        RECT 82.550 179.650 82.810 180.105 ;
        RECT 82.980 179.455 83.240 180.015 ;
        RECT 83.410 179.635 83.660 180.445 ;
        RECT 83.840 179.455 84.100 179.980 ;
        RECT 84.270 179.635 84.520 180.445 ;
        RECT 84.690 180.135 85.005 180.695 ;
        RECT 85.230 180.445 86.890 180.645 ;
        RECT 87.210 180.445 88.575 180.645 ;
        RECT 88.745 180.275 89.145 180.815 ;
        RECT 84.700 179.455 85.005 179.965 ;
        RECT 85.180 179.455 85.455 180.275 ;
        RECT 85.625 180.095 89.145 180.275 ;
        RECT 89.330 180.785 90.085 180.955 ;
        RECT 90.875 180.865 91.905 181.035 ;
        RECT 89.330 180.275 89.735 180.785 ;
        RECT 90.875 180.615 91.045 180.865 ;
        RECT 89.905 180.445 91.045 180.615 ;
        RECT 89.330 180.105 90.980 180.275 ;
        RECT 91.215 180.125 91.565 180.695 ;
        RECT 85.625 179.625 85.955 180.095 ;
        RECT 86.125 179.455 86.295 179.925 ;
        RECT 86.465 179.625 86.795 180.095 ;
        RECT 86.965 179.455 87.135 179.925 ;
        RECT 87.305 179.625 87.635 180.095 ;
        RECT 87.805 179.455 87.975 179.925 ;
        RECT 88.145 179.625 88.475 180.095 ;
        RECT 88.645 179.455 88.930 179.925 ;
        RECT 89.375 179.455 89.655 179.935 ;
        RECT 89.825 179.715 90.085 180.105 ;
        RECT 90.260 179.455 90.515 179.935 ;
        RECT 90.685 179.715 90.980 180.105 ;
        RECT 91.735 179.955 91.905 180.865 ;
        RECT 92.995 180.840 93.285 182.005 ;
        RECT 93.455 180.865 93.840 181.835 ;
        RECT 94.010 181.545 94.335 182.005 ;
        RECT 94.855 181.375 95.135 181.835 ;
        RECT 94.010 181.155 95.135 181.375 ;
        RECT 93.455 180.195 93.735 180.865 ;
        RECT 94.010 180.695 94.460 181.155 ;
        RECT 95.325 180.985 95.725 181.835 ;
        RECT 96.125 181.545 96.395 182.005 ;
        RECT 96.565 181.375 96.850 181.835 ;
        RECT 93.905 180.365 94.460 180.695 ;
        RECT 94.630 180.425 95.725 180.985 ;
        RECT 94.010 180.255 94.460 180.365 ;
        RECT 91.160 179.455 91.435 179.935 ;
        RECT 91.605 179.625 91.905 179.955 ;
        RECT 92.995 179.455 93.285 180.180 ;
        RECT 93.455 179.625 93.840 180.195 ;
        RECT 94.010 180.085 95.135 180.255 ;
        RECT 94.010 179.455 94.335 179.915 ;
        RECT 94.855 179.625 95.135 180.085 ;
        RECT 95.325 179.625 95.725 180.425 ;
        RECT 95.895 181.155 96.850 181.375 ;
        RECT 95.895 180.255 96.105 181.155 ;
        RECT 97.135 181.035 97.445 181.835 ;
        RECT 97.615 181.205 97.925 182.005 ;
        RECT 98.095 181.375 98.355 181.835 ;
        RECT 98.525 181.545 98.780 182.005 ;
        RECT 98.955 181.375 99.215 181.835 ;
        RECT 98.095 181.205 99.215 181.375 ;
        RECT 96.275 180.425 96.965 180.985 ;
        RECT 97.135 180.865 98.165 181.035 ;
        RECT 95.895 180.085 96.850 180.255 ;
        RECT 96.125 179.455 96.395 179.915 ;
        RECT 96.565 179.625 96.850 180.085 ;
        RECT 97.135 179.955 97.305 180.865 ;
        RECT 97.475 180.125 97.825 180.695 ;
        RECT 97.995 180.615 98.165 180.865 ;
        RECT 98.955 180.955 99.215 181.205 ;
        RECT 99.385 181.135 99.670 182.005 ;
        RECT 100.355 181.035 100.665 181.835 ;
        RECT 100.835 181.205 101.145 182.005 ;
        RECT 101.315 181.375 101.575 181.835 ;
        RECT 101.745 181.545 102.000 182.005 ;
        RECT 102.175 181.375 102.435 181.835 ;
        RECT 101.315 181.205 102.435 181.375 ;
        RECT 98.955 180.785 99.710 180.955 ;
        RECT 97.995 180.445 99.135 180.615 ;
        RECT 99.305 180.275 99.710 180.785 ;
        RECT 98.060 180.105 99.710 180.275 ;
        RECT 100.355 180.865 101.385 181.035 ;
        RECT 97.135 179.625 97.435 179.955 ;
        RECT 97.605 179.455 97.880 179.935 ;
        RECT 98.060 179.715 98.355 180.105 ;
        RECT 98.525 179.455 98.780 179.935 ;
        RECT 98.955 179.715 99.215 180.105 ;
        RECT 100.355 179.955 100.525 180.865 ;
        RECT 100.695 180.125 101.045 180.695 ;
        RECT 101.215 180.615 101.385 180.865 ;
        RECT 102.175 180.955 102.435 181.205 ;
        RECT 102.605 181.135 102.890 182.005 ;
        RECT 103.115 181.135 103.390 181.835 ;
        RECT 103.560 181.460 103.815 182.005 ;
        RECT 103.985 181.495 104.465 181.835 ;
        RECT 104.640 181.450 105.245 182.005 ;
        RECT 104.630 181.350 105.245 181.450 ;
        RECT 104.630 181.325 104.815 181.350 ;
        RECT 102.175 180.785 102.930 180.955 ;
        RECT 101.215 180.445 102.355 180.615 ;
        RECT 102.525 180.275 102.930 180.785 ;
        RECT 101.280 180.105 102.930 180.275 ;
        RECT 103.115 180.105 103.285 181.135 ;
        RECT 103.560 181.005 104.315 181.255 ;
        RECT 104.485 181.080 104.815 181.325 ;
        RECT 103.560 180.970 104.330 181.005 ;
        RECT 103.560 180.960 104.345 180.970 ;
        RECT 103.455 180.945 104.350 180.960 ;
        RECT 103.455 180.930 104.370 180.945 ;
        RECT 103.455 180.920 104.390 180.930 ;
        RECT 103.455 180.910 104.415 180.920 ;
        RECT 103.455 180.880 104.485 180.910 ;
        RECT 103.455 180.850 104.505 180.880 ;
        RECT 103.455 180.820 104.525 180.850 ;
        RECT 103.455 180.795 104.555 180.820 ;
        RECT 103.455 180.760 104.590 180.795 ;
        RECT 103.455 180.755 104.620 180.760 ;
        RECT 103.455 180.360 103.685 180.755 ;
        RECT 104.230 180.750 104.620 180.755 ;
        RECT 104.255 180.740 104.620 180.750 ;
        RECT 104.270 180.735 104.620 180.740 ;
        RECT 104.285 180.730 104.620 180.735 ;
        RECT 104.985 180.730 105.245 181.180 ;
        RECT 105.415 180.915 108.925 182.005 ;
        RECT 109.095 180.915 110.305 182.005 ;
        RECT 104.285 180.725 105.245 180.730 ;
        RECT 104.295 180.715 105.245 180.725 ;
        RECT 104.305 180.710 105.245 180.715 ;
        RECT 104.315 180.700 105.245 180.710 ;
        RECT 104.320 180.690 105.245 180.700 ;
        RECT 104.325 180.685 105.245 180.690 ;
        RECT 104.335 180.670 105.245 180.685 ;
        RECT 104.340 180.655 105.245 180.670 ;
        RECT 104.350 180.630 105.245 180.655 ;
        RECT 103.855 180.160 104.185 180.585 ;
        RECT 99.385 179.455 99.665 179.935 ;
        RECT 100.355 179.625 100.655 179.955 ;
        RECT 100.825 179.455 101.100 179.935 ;
        RECT 101.280 179.715 101.575 180.105 ;
        RECT 101.745 179.455 102.000 179.935 ;
        RECT 102.175 179.715 102.435 180.105 ;
        RECT 102.605 179.455 102.885 179.935 ;
        RECT 103.115 179.625 103.375 180.105 ;
        RECT 103.545 179.455 103.795 179.995 ;
        RECT 103.965 179.675 104.185 180.160 ;
        RECT 104.355 180.560 105.245 180.630 ;
        RECT 104.355 179.835 104.525 180.560 ;
        RECT 104.695 180.005 105.245 180.390 ;
        RECT 105.415 180.225 107.065 180.745 ;
        RECT 107.235 180.395 108.925 180.915 ;
        RECT 104.355 179.665 105.245 179.835 ;
        RECT 105.415 179.455 108.925 180.225 ;
        RECT 109.095 180.205 109.615 180.745 ;
        RECT 109.785 180.375 110.305 180.915 ;
        RECT 110.485 181.665 111.655 181.835 ;
        RECT 110.485 180.995 110.815 181.665 ;
        RECT 111.325 181.625 111.655 181.665 ;
        RECT 111.845 181.585 112.200 182.005 ;
        RECT 110.985 181.405 111.215 181.495 ;
        RECT 112.370 181.405 112.620 181.835 ;
        RECT 110.985 181.165 112.620 181.405 ;
        RECT 112.790 181.245 113.120 182.005 ;
        RECT 113.290 181.155 113.550 181.835 ;
        RECT 110.485 180.825 113.205 180.995 ;
        RECT 110.480 180.445 110.965 180.645 ;
        RECT 111.155 180.445 111.630 180.655 ;
        RECT 109.095 179.455 110.305 180.205 ;
        RECT 110.485 179.455 110.935 180.220 ;
        RECT 111.410 180.045 111.630 180.445 ;
        RECT 111.900 180.445 112.230 180.655 ;
        RECT 112.400 180.445 112.805 180.645 ;
        RECT 111.900 180.045 112.110 180.445 ;
        RECT 113.035 180.275 113.205 180.825 ;
        RECT 112.365 180.105 113.205 180.275 ;
        RECT 112.365 179.875 112.535 180.105 ;
        RECT 113.380 179.955 113.550 181.155 ;
        RECT 113.720 180.815 113.890 182.005 ;
        RECT 114.155 180.995 114.415 182.005 ;
        RECT 114.585 181.165 114.860 181.835 ;
        RECT 114.585 180.815 114.755 181.165 ;
        RECT 115.060 181.160 115.275 182.005 ;
        RECT 115.460 181.495 115.935 181.835 ;
        RECT 116.115 181.500 116.745 182.005 ;
        RECT 116.115 181.325 116.305 181.500 ;
        RECT 115.500 180.965 115.750 181.260 ;
        RECT 115.975 181.135 116.305 181.325 ;
        RECT 116.475 180.965 116.730 181.330 ;
        RECT 111.210 179.625 112.535 179.875 ;
        RECT 112.745 179.455 113.075 179.935 ;
        RECT 113.290 179.625 113.550 179.955 ;
        RECT 113.720 179.455 113.890 180.355 ;
        RECT 114.155 180.295 114.770 180.815 ;
        RECT 114.940 180.795 116.730 180.965 ;
        RECT 116.915 180.915 118.585 182.005 ;
        RECT 114.940 180.365 115.170 180.795 ;
        RECT 114.155 179.455 114.430 180.115 ;
        RECT 114.600 180.085 114.770 180.295 ;
        RECT 115.355 180.120 115.765 180.615 ;
        RECT 114.600 179.625 114.850 180.085 ;
        RECT 115.025 179.455 115.355 179.950 ;
        RECT 115.535 179.675 115.765 180.120 ;
        RECT 115.935 179.940 116.190 180.795 ;
        RECT 116.360 180.135 116.745 180.615 ;
        RECT 116.915 180.225 117.665 180.745 ;
        RECT 117.835 180.395 118.585 180.915 ;
        RECT 118.755 180.840 119.045 182.005 ;
        RECT 119.220 181.625 119.555 182.005 ;
        RECT 115.935 179.675 116.725 179.940 ;
        RECT 116.915 179.455 118.585 180.225 ;
        RECT 118.755 179.455 119.045 180.180 ;
        RECT 119.215 180.135 119.455 181.445 ;
        RECT 119.725 181.035 119.975 181.835 ;
        RECT 120.195 181.285 120.525 182.005 ;
        RECT 120.710 181.035 120.960 181.835 ;
        RECT 121.425 181.205 121.755 182.005 ;
        RECT 121.925 181.575 122.265 181.835 ;
        RECT 119.625 180.865 121.815 181.035 ;
        RECT 119.625 179.955 119.795 180.865 ;
        RECT 121.500 180.695 121.815 180.865 ;
        RECT 119.300 179.625 119.795 179.955 ;
        RECT 120.015 179.730 120.365 180.695 ;
        RECT 120.545 179.725 120.845 180.695 ;
        RECT 121.025 179.725 121.305 180.695 ;
        RECT 121.500 180.445 121.830 180.695 ;
        RECT 121.485 179.455 121.755 180.255 ;
        RECT 122.005 180.175 122.265 181.575 ;
        RECT 122.955 181.305 123.175 181.835 ;
        RECT 123.345 181.495 123.675 182.005 ;
        RECT 123.845 181.305 124.070 181.835 ;
        RECT 122.955 181.040 124.070 181.305 ;
        RECT 124.240 181.290 124.555 181.835 ;
        RECT 124.745 181.590 125.075 182.005 ;
        RECT 124.240 181.060 125.075 181.290 ;
        RECT 121.925 179.665 122.265 180.175 ;
        RECT 122.905 180.120 123.220 180.695 ;
        RECT 122.895 179.455 123.225 179.935 ;
        RECT 123.410 179.735 123.790 180.695 ;
        RECT 124.240 180.365 124.565 180.780 ;
        RECT 124.735 180.365 125.075 181.060 ;
        RECT 124.735 180.195 124.905 180.365 ;
        RECT 125.245 180.195 125.475 181.835 ;
        RECT 125.645 181.035 125.935 182.005 ;
        RECT 127.035 180.865 127.295 182.005 ;
        RECT 127.465 181.035 127.795 181.835 ;
        RECT 127.965 181.205 128.135 182.005 ;
        RECT 128.305 181.035 128.635 181.835 ;
        RECT 128.805 181.205 129.060 182.005 ;
        RECT 129.335 181.570 134.680 182.005 ;
        RECT 127.465 180.865 129.165 181.035 ;
        RECT 127.035 180.445 127.795 180.695 ;
        RECT 127.965 180.445 128.715 180.695 ;
        RECT 128.885 180.275 129.165 180.865 ;
        RECT 124.165 180.025 124.905 180.195 ;
        RECT 124.165 179.625 124.355 180.025 ;
        RECT 125.075 180.005 125.475 180.195 ;
        RECT 127.035 180.085 128.135 180.255 ;
        RECT 124.575 179.455 124.905 179.815 ;
        RECT 125.075 179.625 125.265 180.005 ;
        RECT 125.435 179.455 125.765 179.835 ;
        RECT 127.035 179.625 127.375 180.085 ;
        RECT 127.545 179.455 127.715 179.915 ;
        RECT 127.885 179.835 128.135 180.085 ;
        RECT 128.305 180.025 129.165 180.275 ;
        RECT 130.920 180.000 131.260 180.830 ;
        RECT 132.740 180.320 133.090 181.570 ;
        RECT 134.855 180.915 136.525 182.005 ;
        RECT 134.855 180.225 135.605 180.745 ;
        RECT 135.775 180.395 136.525 180.915 ;
        RECT 137.160 180.865 137.495 181.835 ;
        RECT 137.665 180.865 137.835 182.005 ;
        RECT 138.005 181.665 140.035 181.835 ;
        RECT 128.725 179.835 129.055 179.855 ;
        RECT 127.885 179.625 129.055 179.835 ;
        RECT 129.335 179.455 134.680 180.000 ;
        RECT 134.855 179.455 136.525 180.225 ;
        RECT 137.160 180.195 137.330 180.865 ;
        RECT 138.005 180.695 138.175 181.665 ;
        RECT 137.500 180.365 137.755 180.695 ;
        RECT 137.980 180.365 138.175 180.695 ;
        RECT 138.345 181.325 139.470 181.495 ;
        RECT 137.585 180.195 137.755 180.365 ;
        RECT 138.345 180.195 138.515 181.325 ;
        RECT 137.160 179.625 137.415 180.195 ;
        RECT 137.585 180.025 138.515 180.195 ;
        RECT 138.685 180.985 139.695 181.155 ;
        RECT 138.685 180.185 138.855 180.985 ;
        RECT 139.060 180.305 139.335 180.785 ;
        RECT 139.055 180.135 139.335 180.305 ;
        RECT 138.340 179.990 138.515 180.025 ;
        RECT 137.585 179.455 137.915 179.855 ;
        RECT 138.340 179.625 138.870 179.990 ;
        RECT 139.060 179.625 139.335 180.135 ;
        RECT 139.505 179.625 139.695 180.985 ;
        RECT 139.865 181.000 140.035 181.665 ;
        RECT 140.205 181.245 140.375 182.005 ;
        RECT 140.610 181.245 141.125 181.655 ;
        RECT 139.865 180.810 140.615 181.000 ;
        RECT 140.785 180.435 141.125 181.245 ;
        RECT 141.295 180.915 143.885 182.005 ;
        RECT 139.895 180.265 141.125 180.435 ;
        RECT 139.875 179.455 140.385 179.990 ;
        RECT 140.605 179.660 140.850 180.265 ;
        RECT 141.295 180.225 142.505 180.745 ;
        RECT 142.675 180.395 143.885 180.915 ;
        RECT 144.515 180.840 144.805 182.005 ;
        RECT 144.975 181.570 150.320 182.005 ;
        RECT 141.295 179.455 143.885 180.225 ;
        RECT 144.515 179.455 144.805 180.180 ;
        RECT 146.560 180.000 146.900 180.830 ;
        RECT 148.380 180.320 148.730 181.570 ;
        RECT 150.965 181.025 151.295 181.835 ;
        RECT 151.465 181.205 151.705 182.005 ;
        RECT 150.965 180.855 151.680 181.025 ;
        RECT 150.960 180.445 151.340 180.685 ;
        RECT 151.510 180.615 151.680 180.855 ;
        RECT 151.885 180.985 152.055 181.835 ;
        RECT 152.225 181.205 152.555 182.005 ;
        RECT 152.725 180.985 152.895 181.835 ;
        RECT 151.885 180.815 152.895 180.985 ;
        RECT 153.065 180.855 153.395 182.005 ;
        RECT 153.715 180.915 156.305 182.005 ;
        RECT 152.400 180.645 152.895 180.815 ;
        RECT 151.510 180.445 152.010 180.615 ;
        RECT 152.395 180.475 152.895 180.645 ;
        RECT 151.510 180.275 151.680 180.445 ;
        RECT 152.400 180.275 152.895 180.475 ;
        RECT 151.045 180.105 151.680 180.275 ;
        RECT 151.885 180.105 152.895 180.275 ;
        RECT 144.975 179.455 150.320 180.000 ;
        RECT 151.045 179.625 151.215 180.105 ;
        RECT 151.395 179.455 151.635 179.935 ;
        RECT 151.885 179.625 152.055 180.105 ;
        RECT 152.225 179.455 152.555 179.935 ;
        RECT 152.725 179.625 152.895 180.105 ;
        RECT 153.065 179.455 153.395 180.255 ;
        RECT 153.715 180.225 154.925 180.745 ;
        RECT 155.095 180.395 156.305 180.915 ;
        RECT 156.935 180.915 158.145 182.005 ;
        RECT 156.935 180.375 157.455 180.915 ;
        RECT 153.715 179.455 156.305 180.225 ;
        RECT 157.625 180.205 158.145 180.745 ;
        RECT 156.935 179.455 158.145 180.205 ;
        RECT 2.750 179.285 158.230 179.455 ;
        RECT 2.835 178.535 4.045 179.285 ;
        RECT 2.835 177.995 3.355 178.535 ;
        RECT 4.215 178.515 5.885 179.285 ;
        RECT 6.055 178.610 6.315 179.115 ;
        RECT 6.495 178.905 6.825 179.285 ;
        RECT 7.005 178.735 7.175 179.115 ;
        RECT 3.525 177.825 4.045 178.365 ;
        RECT 4.215 177.995 4.965 178.515 ;
        RECT 5.135 177.825 5.885 178.345 ;
        RECT 2.835 176.735 4.045 177.825 ;
        RECT 4.215 176.735 5.885 177.825 ;
        RECT 6.055 177.810 6.225 178.610 ;
        RECT 6.510 178.565 7.175 178.735 ;
        RECT 6.510 178.310 6.680 178.565 ;
        RECT 7.435 178.515 9.105 179.285 ;
        RECT 9.280 178.545 9.535 179.115 ;
        RECT 9.705 178.885 10.035 179.285 ;
        RECT 10.460 178.750 10.990 179.115 ;
        RECT 11.180 178.945 11.455 179.115 ;
        RECT 11.175 178.775 11.455 178.945 ;
        RECT 10.460 178.715 10.635 178.750 ;
        RECT 9.705 178.545 10.635 178.715 ;
        RECT 6.395 177.980 6.680 178.310 ;
        RECT 6.915 178.015 7.245 178.385 ;
        RECT 7.435 177.995 8.185 178.515 ;
        RECT 6.510 177.835 6.680 177.980 ;
        RECT 6.055 176.905 6.325 177.810 ;
        RECT 6.510 177.665 7.175 177.835 ;
        RECT 8.355 177.825 9.105 178.345 ;
        RECT 6.495 176.735 6.825 177.495 ;
        RECT 7.005 176.905 7.175 177.665 ;
        RECT 7.435 176.735 9.105 177.825 ;
        RECT 9.280 177.875 9.450 178.545 ;
        RECT 9.705 178.375 9.875 178.545 ;
        RECT 9.620 178.045 9.875 178.375 ;
        RECT 10.100 178.045 10.295 178.375 ;
        RECT 9.280 176.905 9.615 177.875 ;
        RECT 9.785 176.735 9.955 177.875 ;
        RECT 10.125 177.075 10.295 178.045 ;
        RECT 10.465 177.415 10.635 178.545 ;
        RECT 10.805 177.755 10.975 178.555 ;
        RECT 11.180 177.955 11.455 178.775 ;
        RECT 11.625 177.755 11.815 179.115 ;
        RECT 11.995 178.750 12.505 179.285 ;
        RECT 12.725 178.475 12.970 179.080 ;
        RECT 13.415 178.515 15.085 179.285 ;
        RECT 15.260 178.545 15.515 179.115 ;
        RECT 15.685 178.885 16.015 179.285 ;
        RECT 16.440 178.750 16.970 179.115 ;
        RECT 17.160 178.945 17.435 179.115 ;
        RECT 17.155 178.775 17.435 178.945 ;
        RECT 16.440 178.715 16.615 178.750 ;
        RECT 15.685 178.545 16.615 178.715 ;
        RECT 12.015 178.305 13.245 178.475 ;
        RECT 10.805 177.585 11.815 177.755 ;
        RECT 11.985 177.740 12.735 177.930 ;
        RECT 10.465 177.245 11.590 177.415 ;
        RECT 11.985 177.075 12.155 177.740 ;
        RECT 12.905 177.495 13.245 178.305 ;
        RECT 13.415 177.995 14.165 178.515 ;
        RECT 14.335 177.825 15.085 178.345 ;
        RECT 10.125 176.905 12.155 177.075 ;
        RECT 12.325 176.735 12.495 177.495 ;
        RECT 12.730 177.085 13.245 177.495 ;
        RECT 13.415 176.735 15.085 177.825 ;
        RECT 15.260 177.875 15.430 178.545 ;
        RECT 15.685 178.375 15.855 178.545 ;
        RECT 15.600 178.045 15.855 178.375 ;
        RECT 16.080 178.045 16.275 178.375 ;
        RECT 15.260 176.905 15.595 177.875 ;
        RECT 15.765 176.735 15.935 177.875 ;
        RECT 16.105 177.075 16.275 178.045 ;
        RECT 16.445 177.415 16.615 178.545 ;
        RECT 16.785 177.755 16.955 178.555 ;
        RECT 17.160 177.955 17.435 178.775 ;
        RECT 17.605 177.755 17.795 179.115 ;
        RECT 17.975 178.750 18.485 179.285 ;
        RECT 18.705 178.475 18.950 179.080 ;
        RECT 19.400 178.735 19.655 179.025 ;
        RECT 19.825 178.905 20.155 179.285 ;
        RECT 19.400 178.565 20.150 178.735 ;
        RECT 17.995 178.305 19.225 178.475 ;
        RECT 16.785 177.585 17.795 177.755 ;
        RECT 17.965 177.740 18.715 177.930 ;
        RECT 16.445 177.245 17.570 177.415 ;
        RECT 17.965 177.075 18.135 177.740 ;
        RECT 18.885 177.495 19.225 178.305 ;
        RECT 19.400 177.745 19.750 178.395 ;
        RECT 19.920 177.575 20.150 178.565 ;
        RECT 16.105 176.905 18.135 177.075 ;
        RECT 18.305 176.735 18.475 177.495 ;
        RECT 18.710 177.085 19.225 177.495 ;
        RECT 19.400 177.405 20.150 177.575 ;
        RECT 19.400 176.905 19.655 177.405 ;
        RECT 19.825 176.735 20.155 177.235 ;
        RECT 20.325 176.905 20.495 179.025 ;
        RECT 20.855 178.925 21.185 179.285 ;
        RECT 21.355 178.895 21.850 179.065 ;
        RECT 22.055 178.895 22.910 179.065 ;
        RECT 20.725 177.705 21.185 178.755 ;
        RECT 20.665 176.920 20.990 177.705 ;
        RECT 21.355 177.535 21.525 178.895 ;
        RECT 21.695 177.985 22.045 178.605 ;
        RECT 22.215 178.385 22.570 178.605 ;
        RECT 22.215 177.795 22.385 178.385 ;
        RECT 22.740 178.185 22.910 178.895 ;
        RECT 23.785 178.825 24.115 179.285 ;
        RECT 24.325 178.925 24.675 179.095 ;
        RECT 23.115 178.355 23.905 178.605 ;
        RECT 24.325 178.535 24.585 178.925 ;
        RECT 24.895 178.835 25.845 179.115 ;
        RECT 26.015 178.845 26.205 179.285 ;
        RECT 26.375 178.905 27.445 179.075 ;
        RECT 24.075 178.185 24.245 178.365 ;
        RECT 21.355 177.365 21.750 177.535 ;
        RECT 21.920 177.405 22.385 177.795 ;
        RECT 22.555 178.015 24.245 178.185 ;
        RECT 21.580 177.235 21.750 177.365 ;
        RECT 22.555 177.235 22.725 178.015 ;
        RECT 24.415 177.845 24.585 178.535 ;
        RECT 23.085 177.675 24.585 177.845 ;
        RECT 24.775 177.875 24.985 178.665 ;
        RECT 25.155 178.045 25.505 178.665 ;
        RECT 25.675 178.055 25.845 178.835 ;
        RECT 26.375 178.675 26.545 178.905 ;
        RECT 26.015 178.505 26.545 178.675 ;
        RECT 26.015 178.225 26.235 178.505 ;
        RECT 26.715 178.335 26.955 178.735 ;
        RECT 25.675 177.885 26.080 178.055 ;
        RECT 26.415 177.965 26.955 178.335 ;
        RECT 27.125 178.550 27.445 178.905 ;
        RECT 27.690 178.825 27.995 179.285 ;
        RECT 28.165 178.575 28.420 179.105 ;
        RECT 27.125 178.375 27.450 178.550 ;
        RECT 27.125 178.075 28.040 178.375 ;
        RECT 27.300 178.045 28.040 178.075 ;
        RECT 24.775 177.715 25.450 177.875 ;
        RECT 25.910 177.795 26.080 177.885 ;
        RECT 24.775 177.705 25.740 177.715 ;
        RECT 24.415 177.535 24.585 177.675 ;
        RECT 21.160 176.735 21.410 177.195 ;
        RECT 21.580 176.905 21.830 177.235 ;
        RECT 22.045 176.905 22.725 177.235 ;
        RECT 22.895 177.335 23.970 177.505 ;
        RECT 24.415 177.365 24.975 177.535 ;
        RECT 25.280 177.415 25.740 177.705 ;
        RECT 25.910 177.625 27.130 177.795 ;
        RECT 22.895 176.995 23.065 177.335 ;
        RECT 23.300 176.735 23.630 177.165 ;
        RECT 23.800 176.995 23.970 177.335 ;
        RECT 24.265 176.735 24.635 177.195 ;
        RECT 24.805 176.905 24.975 177.365 ;
        RECT 25.910 177.245 26.080 177.625 ;
        RECT 27.300 177.455 27.470 178.045 ;
        RECT 28.210 177.925 28.420 178.575 ;
        RECT 28.595 178.560 28.885 179.285 ;
        RECT 29.975 178.610 30.235 179.115 ;
        RECT 30.415 178.905 30.745 179.285 ;
        RECT 30.925 178.735 31.095 179.115 ;
        RECT 25.210 176.905 26.080 177.245 ;
        RECT 26.670 177.285 27.470 177.455 ;
        RECT 26.250 176.735 26.500 177.195 ;
        RECT 26.670 176.995 26.840 177.285 ;
        RECT 27.020 176.735 27.350 177.115 ;
        RECT 27.690 176.735 27.995 177.875 ;
        RECT 28.165 177.045 28.420 177.925 ;
        RECT 28.595 176.735 28.885 177.900 ;
        RECT 29.975 177.810 30.145 178.610 ;
        RECT 30.430 178.565 31.095 178.735 ;
        RECT 31.445 178.735 31.615 179.115 ;
        RECT 31.795 178.905 32.125 179.285 ;
        RECT 31.445 178.565 32.110 178.735 ;
        RECT 32.305 178.610 32.565 179.115 ;
        RECT 30.430 178.310 30.600 178.565 ;
        RECT 30.315 177.980 30.600 178.310 ;
        RECT 30.835 178.015 31.165 178.385 ;
        RECT 31.375 178.015 31.705 178.385 ;
        RECT 31.940 178.310 32.110 178.565 ;
        RECT 30.430 177.835 30.600 177.980 ;
        RECT 31.940 177.980 32.225 178.310 ;
        RECT 31.940 177.835 32.110 177.980 ;
        RECT 29.975 176.905 30.245 177.810 ;
        RECT 30.430 177.665 31.095 177.835 ;
        RECT 30.415 176.735 30.745 177.495 ;
        RECT 30.925 176.905 31.095 177.665 ;
        RECT 31.445 177.665 32.110 177.835 ;
        RECT 32.395 177.810 32.565 178.610 ;
        RECT 32.740 178.735 32.995 179.025 ;
        RECT 33.165 178.905 33.495 179.285 ;
        RECT 32.740 178.565 33.490 178.735 ;
        RECT 31.445 176.905 31.615 177.665 ;
        RECT 31.795 176.735 32.125 177.495 ;
        RECT 32.295 176.905 32.565 177.810 ;
        RECT 32.740 177.745 33.090 178.395 ;
        RECT 33.260 177.575 33.490 178.565 ;
        RECT 32.740 177.405 33.490 177.575 ;
        RECT 32.740 176.905 32.995 177.405 ;
        RECT 33.165 176.735 33.495 177.235 ;
        RECT 33.665 176.905 33.835 179.025 ;
        RECT 34.195 178.925 34.525 179.285 ;
        RECT 34.695 178.895 35.190 179.065 ;
        RECT 35.395 178.895 36.250 179.065 ;
        RECT 34.065 177.705 34.525 178.755 ;
        RECT 34.005 176.920 34.330 177.705 ;
        RECT 34.695 177.535 34.865 178.895 ;
        RECT 35.035 177.985 35.385 178.605 ;
        RECT 35.555 178.385 35.910 178.605 ;
        RECT 35.555 177.795 35.725 178.385 ;
        RECT 36.080 178.185 36.250 178.895 ;
        RECT 37.125 178.825 37.455 179.285 ;
        RECT 37.665 178.925 38.015 179.095 ;
        RECT 36.455 178.355 37.245 178.605 ;
        RECT 37.665 178.535 37.925 178.925 ;
        RECT 38.235 178.835 39.185 179.115 ;
        RECT 39.355 178.845 39.545 179.285 ;
        RECT 39.715 178.905 40.785 179.075 ;
        RECT 37.415 178.185 37.585 178.365 ;
        RECT 34.695 177.365 35.090 177.535 ;
        RECT 35.260 177.405 35.725 177.795 ;
        RECT 35.895 178.015 37.585 178.185 ;
        RECT 34.920 177.235 35.090 177.365 ;
        RECT 35.895 177.235 36.065 178.015 ;
        RECT 37.755 177.845 37.925 178.535 ;
        RECT 36.425 177.675 37.925 177.845 ;
        RECT 38.115 177.875 38.325 178.665 ;
        RECT 38.495 178.045 38.845 178.665 ;
        RECT 39.015 178.055 39.185 178.835 ;
        RECT 39.715 178.675 39.885 178.905 ;
        RECT 39.355 178.505 39.885 178.675 ;
        RECT 39.355 178.225 39.575 178.505 ;
        RECT 40.055 178.335 40.295 178.735 ;
        RECT 39.015 177.885 39.420 178.055 ;
        RECT 39.755 177.965 40.295 178.335 ;
        RECT 40.465 178.550 40.785 178.905 ;
        RECT 41.030 178.825 41.335 179.285 ;
        RECT 41.505 178.575 41.760 179.105 ;
        RECT 40.465 178.375 40.790 178.550 ;
        RECT 40.465 178.075 41.380 178.375 ;
        RECT 40.640 178.045 41.380 178.075 ;
        RECT 38.115 177.715 38.790 177.875 ;
        RECT 39.250 177.795 39.420 177.885 ;
        RECT 38.115 177.705 39.080 177.715 ;
        RECT 37.755 177.535 37.925 177.675 ;
        RECT 34.500 176.735 34.750 177.195 ;
        RECT 34.920 176.905 35.170 177.235 ;
        RECT 35.385 176.905 36.065 177.235 ;
        RECT 36.235 177.335 37.310 177.505 ;
        RECT 37.755 177.365 38.315 177.535 ;
        RECT 38.620 177.415 39.080 177.705 ;
        RECT 39.250 177.625 40.470 177.795 ;
        RECT 36.235 176.995 36.405 177.335 ;
        RECT 36.640 176.735 36.970 177.165 ;
        RECT 37.140 176.995 37.310 177.335 ;
        RECT 37.605 176.735 37.975 177.195 ;
        RECT 38.145 176.905 38.315 177.365 ;
        RECT 39.250 177.245 39.420 177.625 ;
        RECT 40.640 177.455 40.810 178.045 ;
        RECT 41.550 177.925 41.760 178.575 ;
        RECT 41.945 178.475 42.215 179.285 ;
        RECT 42.385 178.475 42.715 179.115 ;
        RECT 42.885 178.475 43.125 179.285 ;
        RECT 43.480 178.775 43.720 179.285 ;
        RECT 43.900 178.775 44.180 179.105 ;
        RECT 44.410 178.775 44.625 179.285 ;
        RECT 41.935 178.045 42.285 178.295 ;
        RECT 38.550 176.905 39.420 177.245 ;
        RECT 40.010 177.285 40.810 177.455 ;
        RECT 39.590 176.735 39.840 177.195 ;
        RECT 40.010 176.995 40.180 177.285 ;
        RECT 40.360 176.735 40.690 177.115 ;
        RECT 41.030 176.735 41.335 177.875 ;
        RECT 41.505 177.045 41.760 177.925 ;
        RECT 42.455 177.875 42.625 178.475 ;
        RECT 42.795 178.045 43.145 178.295 ;
        RECT 43.375 178.045 43.730 178.605 ;
        RECT 43.900 177.875 44.070 178.775 ;
        RECT 44.240 178.045 44.505 178.605 ;
        RECT 44.795 178.545 45.410 179.115 ;
        RECT 44.755 177.875 44.925 178.375 ;
        RECT 41.945 176.735 42.275 177.875 ;
        RECT 42.455 177.705 43.135 177.875 ;
        RECT 42.805 176.920 43.135 177.705 ;
        RECT 43.500 177.705 44.925 177.875 ;
        RECT 43.500 177.530 43.890 177.705 ;
        RECT 44.375 176.735 44.705 177.535 ;
        RECT 45.095 177.525 45.410 178.545 ;
        RECT 44.875 176.905 45.410 177.525 ;
        RECT 45.615 178.635 45.875 179.115 ;
        RECT 46.045 178.745 46.295 179.285 ;
        RECT 45.615 177.605 45.785 178.635 ;
        RECT 46.465 178.580 46.685 179.065 ;
        RECT 45.955 177.985 46.185 178.380 ;
        RECT 46.355 178.155 46.685 178.580 ;
        RECT 46.855 178.905 47.745 179.075 ;
        RECT 46.855 178.180 47.025 178.905 ;
        RECT 47.195 178.350 47.745 178.735 ;
        RECT 48.005 178.635 48.175 179.115 ;
        RECT 48.345 178.805 48.675 179.285 ;
        RECT 48.900 178.865 50.435 179.115 ;
        RECT 48.900 178.635 49.070 178.865 ;
        RECT 48.005 178.465 49.070 178.635 ;
        RECT 49.250 178.295 49.530 178.695 ;
        RECT 46.855 178.110 47.745 178.180 ;
        RECT 46.850 178.085 47.745 178.110 ;
        RECT 47.920 178.085 48.270 178.295 ;
        RECT 48.440 178.095 48.885 178.295 ;
        RECT 49.055 178.095 49.530 178.295 ;
        RECT 49.800 178.295 50.085 178.695 ;
        RECT 50.265 178.635 50.435 178.865 ;
        RECT 50.605 178.805 50.935 179.285 ;
        RECT 51.150 178.785 51.405 179.115 ;
        RECT 51.220 178.705 51.405 178.785 ;
        RECT 50.265 178.465 51.065 178.635 ;
        RECT 49.800 178.095 50.130 178.295 ;
        RECT 50.300 178.095 50.665 178.295 ;
        RECT 46.840 178.070 47.745 178.085 ;
        RECT 46.835 178.055 47.745 178.070 ;
        RECT 46.825 178.050 47.745 178.055 ;
        RECT 46.820 178.040 47.745 178.050 ;
        RECT 46.815 178.030 47.745 178.040 ;
        RECT 46.805 178.025 47.745 178.030 ;
        RECT 46.795 178.015 47.745 178.025 ;
        RECT 46.785 178.010 47.745 178.015 ;
        RECT 46.785 178.005 47.120 178.010 ;
        RECT 46.770 178.000 47.120 178.005 ;
        RECT 46.755 177.990 47.120 178.000 ;
        RECT 46.730 177.985 47.120 177.990 ;
        RECT 45.955 177.980 47.120 177.985 ;
        RECT 45.955 177.945 47.090 177.980 ;
        RECT 45.955 177.920 47.055 177.945 ;
        RECT 45.955 177.890 47.025 177.920 ;
        RECT 45.955 177.860 47.005 177.890 ;
        RECT 45.955 177.830 46.985 177.860 ;
        RECT 45.955 177.820 46.915 177.830 ;
        RECT 45.955 177.810 46.890 177.820 ;
        RECT 45.955 177.795 46.870 177.810 ;
        RECT 45.955 177.780 46.850 177.795 ;
        RECT 46.060 177.770 46.845 177.780 ;
        RECT 46.060 177.735 46.830 177.770 ;
        RECT 45.615 176.905 45.890 177.605 ;
        RECT 46.060 177.485 46.815 177.735 ;
        RECT 46.985 177.415 47.315 177.660 ;
        RECT 47.485 177.560 47.745 178.010 ;
        RECT 50.895 177.915 51.065 178.465 ;
        RECT 48.005 177.745 51.065 177.915 ;
        RECT 47.130 177.390 47.315 177.415 ;
        RECT 47.130 177.290 47.745 177.390 ;
        RECT 46.060 176.735 46.315 177.280 ;
        RECT 46.485 176.905 46.965 177.245 ;
        RECT 47.140 176.735 47.745 177.290 ;
        RECT 48.005 176.905 48.175 177.745 ;
        RECT 51.235 177.575 51.405 178.705 ;
        RECT 48.345 177.075 48.675 177.575 ;
        RECT 48.845 177.335 50.480 177.575 ;
        RECT 48.845 177.245 49.075 177.335 ;
        RECT 49.185 177.075 49.515 177.115 ;
        RECT 48.345 176.905 49.515 177.075 ;
        RECT 49.705 176.735 50.060 177.155 ;
        RECT 50.230 176.905 50.480 177.335 ;
        RECT 50.650 176.735 50.980 177.495 ;
        RECT 51.150 176.905 51.405 177.575 ;
        RECT 51.595 178.785 51.895 179.115 ;
        RECT 52.065 178.805 52.340 179.285 ;
        RECT 51.595 177.875 51.765 178.785 ;
        RECT 52.520 178.635 52.815 179.025 ;
        RECT 52.985 178.805 53.240 179.285 ;
        RECT 53.415 178.635 53.675 179.025 ;
        RECT 53.845 178.805 54.125 179.285 ;
        RECT 51.935 178.045 52.285 178.615 ;
        RECT 52.520 178.465 54.170 178.635 ;
        RECT 54.355 178.560 54.645 179.285 ;
        RECT 55.280 178.785 55.615 179.285 ;
        RECT 55.815 178.715 55.985 179.065 ;
        RECT 56.185 178.885 56.515 179.285 ;
        RECT 56.685 178.715 56.855 179.065 ;
        RECT 57.025 178.885 57.405 179.285 ;
        RECT 52.455 178.125 53.595 178.295 ;
        RECT 52.455 177.875 52.625 178.125 ;
        RECT 53.765 177.955 54.170 178.465 ;
        RECT 55.275 178.045 55.630 178.615 ;
        RECT 55.815 178.545 57.425 178.715 ;
        RECT 57.595 178.610 57.870 178.955 ;
        RECT 57.255 178.375 57.425 178.545 ;
        RECT 51.595 177.705 52.625 177.875 ;
        RECT 53.415 177.785 54.170 177.955 ;
        RECT 51.595 176.905 51.905 177.705 ;
        RECT 53.415 177.535 53.675 177.785 ;
        RECT 52.075 176.735 52.385 177.535 ;
        RECT 52.555 177.365 53.675 177.535 ;
        RECT 52.555 176.905 52.815 177.365 ;
        RECT 52.985 176.735 53.240 177.195 ;
        RECT 53.415 176.905 53.675 177.365 ;
        RECT 53.845 176.735 54.130 177.605 ;
        RECT 54.355 176.735 54.645 177.900 ;
        RECT 55.275 177.585 55.600 177.875 ;
        RECT 55.800 177.755 56.510 178.375 ;
        RECT 56.680 178.045 57.085 178.375 ;
        RECT 57.255 178.045 57.530 178.375 ;
        RECT 57.255 177.875 57.425 178.045 ;
        RECT 57.700 177.875 57.870 178.610 ;
        RECT 58.040 178.370 58.210 179.285 ;
        RECT 58.500 178.735 58.755 179.025 ;
        RECT 58.925 178.905 59.255 179.285 ;
        RECT 58.500 178.565 59.250 178.735 ;
        RECT 56.700 177.705 57.425 177.875 ;
        RECT 56.700 177.585 56.870 177.705 ;
        RECT 55.275 177.415 56.870 177.585 ;
        RECT 55.275 176.955 56.935 177.245 ;
        RECT 57.105 176.735 57.385 177.535 ;
        RECT 57.595 176.905 57.870 177.875 ;
        RECT 58.040 176.735 58.210 177.915 ;
        RECT 58.500 177.745 58.850 178.395 ;
        RECT 59.020 177.575 59.250 178.565 ;
        RECT 58.500 177.405 59.250 177.575 ;
        RECT 58.500 176.905 58.755 177.405 ;
        RECT 58.925 176.735 59.255 177.235 ;
        RECT 59.425 176.905 59.595 179.025 ;
        RECT 59.955 178.925 60.285 179.285 ;
        RECT 60.455 178.895 60.950 179.065 ;
        RECT 61.155 178.895 62.010 179.065 ;
        RECT 59.825 177.705 60.285 178.755 ;
        RECT 59.765 176.920 60.090 177.705 ;
        RECT 60.455 177.535 60.625 178.895 ;
        RECT 60.795 177.985 61.145 178.605 ;
        RECT 61.315 178.385 61.670 178.605 ;
        RECT 61.315 177.795 61.485 178.385 ;
        RECT 61.840 178.185 62.010 178.895 ;
        RECT 62.885 178.825 63.215 179.285 ;
        RECT 63.425 178.925 63.775 179.095 ;
        RECT 62.215 178.355 63.005 178.605 ;
        RECT 63.425 178.535 63.685 178.925 ;
        RECT 63.995 178.835 64.945 179.115 ;
        RECT 65.115 178.845 65.305 179.285 ;
        RECT 65.475 178.905 66.545 179.075 ;
        RECT 63.175 178.185 63.345 178.365 ;
        RECT 60.455 177.365 60.850 177.535 ;
        RECT 61.020 177.405 61.485 177.795 ;
        RECT 61.655 178.015 63.345 178.185 ;
        RECT 60.680 177.235 60.850 177.365 ;
        RECT 61.655 177.235 61.825 178.015 ;
        RECT 63.515 177.845 63.685 178.535 ;
        RECT 62.185 177.675 63.685 177.845 ;
        RECT 63.875 177.875 64.085 178.665 ;
        RECT 64.255 178.045 64.605 178.665 ;
        RECT 64.775 178.055 64.945 178.835 ;
        RECT 65.475 178.675 65.645 178.905 ;
        RECT 65.115 178.505 65.645 178.675 ;
        RECT 65.115 178.225 65.335 178.505 ;
        RECT 65.815 178.335 66.055 178.735 ;
        RECT 64.775 177.885 65.180 178.055 ;
        RECT 65.515 177.965 66.055 178.335 ;
        RECT 66.225 178.550 66.545 178.905 ;
        RECT 66.225 178.295 66.550 178.550 ;
        RECT 66.745 178.475 66.915 179.285 ;
        RECT 67.085 178.635 67.415 179.115 ;
        RECT 67.585 178.815 67.755 179.285 ;
        RECT 67.925 178.635 68.255 179.115 ;
        RECT 68.425 178.815 68.595 179.285 ;
        RECT 67.085 178.465 68.850 178.635 ;
        RECT 66.225 178.085 68.255 178.295 ;
        RECT 66.225 178.075 66.570 178.085 ;
        RECT 63.875 177.715 64.550 177.875 ;
        RECT 65.010 177.795 65.180 177.885 ;
        RECT 63.875 177.705 64.840 177.715 ;
        RECT 63.515 177.535 63.685 177.675 ;
        RECT 60.260 176.735 60.510 177.195 ;
        RECT 60.680 176.905 60.930 177.235 ;
        RECT 61.145 176.905 61.825 177.235 ;
        RECT 61.995 177.335 63.070 177.505 ;
        RECT 63.515 177.365 64.075 177.535 ;
        RECT 64.380 177.415 64.840 177.705 ;
        RECT 65.010 177.625 66.230 177.795 ;
        RECT 61.995 176.995 62.165 177.335 ;
        RECT 62.400 176.735 62.730 177.165 ;
        RECT 62.900 176.995 63.070 177.335 ;
        RECT 63.365 176.735 63.735 177.195 ;
        RECT 63.905 176.905 64.075 177.365 ;
        RECT 65.010 177.245 65.180 177.625 ;
        RECT 66.400 177.455 66.570 178.075 ;
        RECT 68.440 177.915 68.850 178.465 ;
        RECT 69.075 178.515 71.665 179.285 ;
        RECT 71.890 178.890 72.590 179.060 ;
        RECT 72.835 178.920 74.290 179.100 ;
        RECT 71.890 178.775 72.060 178.890 ;
        RECT 72.835 178.715 73.005 178.920 ;
        RECT 74.650 178.915 75.965 179.115 ;
        RECT 76.135 178.925 76.465 179.285 ;
        RECT 76.995 178.925 77.325 179.285 ;
        RECT 75.735 178.745 75.965 178.915 ;
        RECT 77.935 178.845 78.105 179.285 ;
        RECT 78.330 178.745 78.545 178.945 ;
        RECT 78.715 178.925 79.045 179.285 ;
        RECT 79.215 178.745 79.415 178.835 ;
        RECT 72.220 178.545 73.005 178.715 ;
        RECT 73.400 178.555 75.565 178.735 ;
        RECT 75.735 178.675 77.795 178.745 ;
        RECT 78.330 178.675 79.415 178.745 ;
        RECT 75.735 178.575 79.415 178.675 ;
        RECT 69.075 177.995 70.285 178.515 ;
        RECT 64.310 176.905 65.180 177.245 ;
        RECT 65.770 177.285 66.570 177.455 ;
        RECT 65.350 176.735 65.600 177.195 ;
        RECT 65.770 176.995 65.940 177.285 ;
        RECT 66.120 176.735 66.450 177.115 ;
        RECT 66.745 176.735 66.915 177.795 ;
        RECT 67.125 177.745 68.850 177.915 ;
        RECT 70.455 177.825 71.665 178.345 ;
        RECT 72.220 178.030 72.400 178.545 ;
        RECT 76.440 178.505 79.415 178.575 ;
        RECT 80.115 178.560 80.405 179.285 ;
        RECT 80.575 178.560 80.835 179.115 ;
        RECT 81.005 178.840 81.435 179.285 ;
        RECT 81.670 178.715 81.840 179.115 ;
        RECT 82.010 178.885 82.730 179.285 ;
        RECT 77.775 178.465 79.415 178.505 ;
        RECT 67.125 176.905 67.415 177.745 ;
        RECT 67.585 176.735 67.755 177.575 ;
        RECT 67.965 176.905 68.215 177.745 ;
        RECT 68.425 176.735 68.595 177.575 ;
        RECT 69.075 176.735 71.665 177.825 ;
        RECT 71.890 177.515 72.400 178.030 ;
        RECT 72.570 177.855 72.740 178.375 ;
        RECT 73.130 178.025 74.200 178.295 ;
        RECT 74.595 177.960 75.770 178.375 ;
        RECT 74.595 177.855 75.310 177.960 ;
        RECT 72.570 177.685 75.310 177.855 ;
        RECT 75.940 177.855 76.220 178.375 ;
        RECT 76.390 178.025 77.865 178.295 ;
        RECT 78.160 178.040 79.170 178.295 ;
        RECT 78.160 177.855 78.605 178.040 ;
        RECT 75.940 177.685 78.605 177.855 ;
        RECT 75.575 177.515 75.745 177.585 ;
        RECT 71.890 177.345 77.765 177.515 ;
        RECT 78.795 177.435 79.015 177.510 ;
        RECT 71.890 177.265 75.525 177.345 ;
        RECT 76.100 177.265 77.765 177.345 ;
        RECT 77.935 177.265 79.015 177.435 ;
        RECT 71.885 176.735 72.215 177.095 ;
        RECT 73.115 176.735 73.450 177.095 ;
        RECT 73.960 176.735 74.290 177.095 ;
        RECT 74.805 176.735 75.135 177.095 ;
        RECT 75.685 176.735 75.955 177.175 ;
        RECT 77.935 177.095 78.115 177.265 ;
        RECT 78.795 177.180 79.015 177.265 ;
        RECT 76.135 176.905 78.115 177.095 ;
        RECT 78.285 176.735 78.615 177.095 ;
        RECT 79.185 176.735 79.480 177.705 ;
        RECT 80.115 176.735 80.405 177.900 ;
        RECT 80.575 177.845 80.750 178.560 ;
        RECT 81.670 178.545 82.550 178.715 ;
        RECT 82.900 178.670 83.070 179.115 ;
        RECT 83.645 178.775 84.045 179.285 ;
        RECT 80.920 178.045 81.175 178.375 ;
        RECT 80.575 176.905 80.835 177.845 ;
        RECT 81.005 177.565 81.175 178.045 ;
        RECT 81.400 177.755 81.730 178.375 ;
        RECT 81.900 177.995 82.190 178.375 ;
        RECT 82.380 177.825 82.550 178.545 ;
        RECT 82.030 177.655 82.550 177.825 ;
        RECT 82.720 178.500 83.070 178.670 ;
        RECT 81.005 177.395 81.765 177.565 ;
        RECT 82.030 177.465 82.200 177.655 ;
        RECT 82.720 177.475 82.890 178.500 ;
        RECT 83.310 178.015 83.570 178.605 ;
        RECT 83.090 177.715 83.570 178.015 ;
        RECT 83.770 177.715 84.030 178.605 ;
        RECT 84.725 178.565 85.055 179.285 ;
        RECT 85.600 178.885 87.215 179.055 ;
        RECT 87.385 178.885 87.715 179.285 ;
        RECT 87.045 178.715 87.215 178.885 ;
        RECT 87.885 178.810 88.220 179.070 ;
        RECT 88.575 178.905 88.905 179.285 ;
        RECT 84.780 178.265 85.130 178.375 ;
        RECT 84.775 178.095 85.130 178.265 ;
        RECT 84.780 178.045 85.130 178.095 ;
        RECT 85.440 178.045 85.860 178.710 ;
        RECT 86.030 178.265 86.320 178.705 ;
        RECT 86.510 178.265 86.780 178.705 ;
        RECT 87.045 178.545 87.605 178.715 ;
        RECT 87.435 178.375 87.605 178.545 ;
        RECT 86.990 178.265 87.240 178.375 ;
        RECT 86.030 178.095 86.325 178.265 ;
        RECT 86.510 178.095 86.785 178.265 ;
        RECT 86.990 178.095 87.245 178.265 ;
        RECT 86.030 178.045 86.320 178.095 ;
        RECT 86.510 178.045 86.780 178.095 ;
        RECT 86.990 178.045 87.240 178.095 ;
        RECT 87.435 178.045 87.740 178.375 ;
        RECT 84.780 177.755 84.985 178.045 ;
        RECT 87.435 177.875 87.605 178.045 ;
        RECT 85.235 177.705 87.605 177.875 ;
        RECT 81.595 177.170 81.765 177.395 ;
        RECT 82.480 177.305 82.890 177.475 ;
        RECT 83.065 177.365 84.005 177.535 ;
        RECT 82.480 177.170 82.735 177.305 ;
        RECT 81.005 176.735 81.335 177.135 ;
        RECT 81.595 177.000 82.735 177.170 ;
        RECT 83.065 177.115 83.235 177.365 ;
        RECT 82.480 176.905 82.735 177.000 ;
        RECT 82.905 176.945 83.235 177.115 ;
        RECT 83.405 176.735 83.655 177.195 ;
        RECT 83.825 176.905 84.005 177.365 ;
        RECT 84.805 177.075 84.975 177.575 ;
        RECT 85.235 177.245 85.405 177.705 ;
        RECT 85.635 177.325 87.060 177.495 ;
        RECT 85.635 177.075 85.965 177.325 ;
        RECT 84.805 176.905 85.965 177.075 ;
        RECT 86.190 176.735 86.520 177.155 ;
        RECT 86.775 176.905 87.060 177.325 ;
        RECT 87.305 176.735 87.635 177.535 ;
        RECT 87.965 177.455 88.220 178.810 ;
        RECT 89.075 178.735 89.265 179.115 ;
        RECT 89.435 178.925 89.765 179.285 ;
        RECT 88.865 178.545 89.265 178.735 ;
        RECT 89.985 178.715 90.175 179.115 ;
        RECT 89.435 178.545 90.175 178.715 ;
        RECT 87.885 176.945 88.220 177.455 ;
        RECT 88.405 176.735 88.695 177.705 ;
        RECT 88.865 176.905 89.095 178.545 ;
        RECT 89.435 178.375 89.605 178.545 ;
        RECT 89.265 177.680 89.605 178.375 ;
        RECT 89.775 177.960 90.100 178.375 ;
        RECT 90.550 178.045 90.930 179.005 ;
        RECT 91.115 178.805 91.445 179.285 ;
        RECT 91.705 178.735 91.875 179.115 ;
        RECT 92.090 178.905 92.420 179.285 ;
        RECT 91.120 178.045 91.435 178.620 ;
        RECT 91.705 178.565 92.420 178.735 ;
        RECT 91.615 178.015 91.970 178.385 ;
        RECT 92.250 178.375 92.420 178.565 ;
        RECT 92.590 178.540 92.845 179.115 ;
        RECT 92.250 178.045 92.505 178.375 ;
        RECT 92.250 177.835 92.420 178.045 ;
        RECT 89.265 177.450 90.100 177.680 ;
        RECT 89.265 176.735 89.595 177.150 ;
        RECT 89.785 176.905 90.100 177.450 ;
        RECT 90.270 177.435 91.385 177.700 ;
        RECT 90.270 176.905 90.495 177.435 ;
        RECT 90.665 176.735 90.995 177.245 ;
        RECT 91.165 176.905 91.385 177.435 ;
        RECT 91.705 177.665 92.420 177.835 ;
        RECT 92.675 177.810 92.845 178.540 ;
        RECT 93.020 178.445 93.280 179.285 ;
        RECT 93.465 178.905 93.795 179.285 ;
        RECT 93.965 178.755 94.135 179.115 ;
        RECT 94.305 178.925 94.635 179.285 ;
        RECT 94.805 178.755 94.975 179.115 ;
        RECT 95.145 178.905 95.510 179.285 ;
        RECT 95.700 178.905 97.870 179.115 ;
        RECT 93.965 178.735 94.975 178.755 ;
        RECT 93.455 178.565 94.975 178.735 ;
        RECT 93.455 177.935 93.735 178.565 ;
        RECT 95.570 178.555 96.890 178.735 ;
        RECT 97.540 178.675 97.870 178.905 ;
        RECT 98.040 178.845 98.355 179.285 ;
        RECT 98.525 178.675 98.855 179.115 ;
        RECT 99.025 178.845 99.215 179.285 ;
        RECT 99.385 178.675 99.715 179.115 ;
        RECT 95.570 178.305 95.740 178.555 ;
        RECT 97.540 178.505 99.715 178.675 ;
        RECT 99.895 178.645 100.235 179.115 ;
        RECT 100.405 178.815 100.575 179.285 ;
        RECT 100.745 178.645 101.075 179.115 ;
        RECT 101.245 178.815 101.945 179.285 ;
        RECT 99.895 178.465 101.900 178.645 ;
        RECT 102.115 178.635 102.445 179.105 ;
        RECT 102.615 178.815 102.785 179.285 ;
        RECT 102.955 178.635 103.285 179.105 ;
        RECT 103.455 178.815 103.625 179.285 ;
        RECT 102.115 178.465 103.865 178.635 ;
        RECT 93.905 178.105 95.740 178.305 ;
        RECT 91.705 176.905 91.875 177.665 ;
        RECT 92.090 176.735 92.420 177.495 ;
        RECT 92.590 176.905 92.845 177.810 ;
        RECT 93.020 176.735 93.280 177.885 ;
        RECT 93.455 177.670 95.400 177.935 ;
        RECT 93.850 176.735 94.180 177.500 ;
        RECT 94.350 176.905 94.530 177.670 ;
        RECT 94.710 176.735 95.040 177.500 ;
        RECT 95.210 176.905 95.400 177.670 ;
        RECT 95.570 177.515 95.740 178.105 ;
        RECT 95.910 177.925 96.200 178.375 ;
        RECT 96.425 178.095 97.110 178.335 ;
        RECT 97.320 177.925 97.650 178.335 ;
        RECT 95.910 177.685 97.650 177.925 ;
        RECT 97.860 177.875 98.215 178.335 ;
        RECT 98.400 178.045 99.075 178.335 ;
        RECT 99.260 178.265 99.660 178.335 ;
        RECT 101.680 178.295 101.900 178.465 ;
        RECT 99.260 178.095 99.665 178.265 ;
        RECT 99.260 177.875 99.660 178.095 ;
        RECT 99.895 178.045 100.235 178.295 ;
        RECT 100.405 178.045 100.865 178.295 ;
        RECT 101.035 178.045 101.510 178.295 ;
        RECT 101.680 178.125 103.405 178.295 ;
        RECT 97.860 177.685 99.660 177.875 ;
        RECT 95.570 177.345 98.855 177.515 ;
        RECT 95.570 176.735 95.900 177.170 ;
        RECT 96.070 176.905 96.430 177.345 ;
        RECT 96.655 176.735 96.985 177.175 ;
        RECT 97.155 176.905 97.490 177.345 ;
        RECT 97.660 176.735 97.925 177.175 ;
        RECT 98.525 176.905 98.855 177.345 ;
        RECT 99.385 176.735 99.715 177.455 ;
        RECT 99.895 177.075 100.235 177.875 ;
        RECT 100.405 177.320 100.640 178.045 ;
        RECT 101.680 177.875 101.900 178.125 ;
        RECT 102.715 177.915 102.885 177.925 ;
        RECT 103.575 177.915 103.865 178.465 ;
        RECT 104.035 178.515 105.705 179.285 ;
        RECT 105.875 178.560 106.165 179.285 ;
        RECT 106.345 178.675 106.675 179.095 ;
        RECT 106.845 178.845 107.120 179.285 ;
        RECT 107.325 178.675 107.655 179.095 ;
        RECT 108.135 178.925 108.985 179.285 ;
        RECT 109.155 178.735 109.375 179.115 ;
        RECT 104.035 177.995 104.785 178.515 ;
        RECT 106.345 178.495 108.930 178.675 ;
        RECT 100.810 177.705 101.900 177.875 ;
        RECT 102.155 177.745 103.865 177.915 ;
        RECT 104.955 177.825 105.705 178.345 ;
        RECT 106.335 178.095 106.670 178.325 ;
        RECT 106.860 178.265 107.310 178.325 ;
        RECT 106.855 178.095 107.310 178.265 ;
        RECT 107.480 178.095 107.950 178.325 ;
        RECT 108.120 178.095 108.450 178.325 ;
        RECT 100.810 177.075 101.075 177.705 ;
        RECT 99.895 176.905 101.075 177.075 ;
        RECT 101.245 176.735 101.945 177.535 ;
        RECT 102.155 176.905 102.405 177.745 ;
        RECT 102.575 176.735 102.825 177.575 ;
        RECT 102.995 176.905 103.245 177.745 ;
        RECT 103.415 176.735 103.665 177.575 ;
        RECT 104.035 176.735 105.705 177.825 ;
        RECT 105.875 176.735 106.165 177.900 ;
        RECT 108.620 177.880 108.930 178.495 ;
        RECT 106.345 177.710 108.930 177.880 ;
        RECT 106.345 177.045 106.675 177.710 ;
        RECT 107.135 177.350 108.475 177.530 ;
        RECT 107.135 176.905 107.465 177.350 ;
        RECT 107.700 176.735 107.975 177.180 ;
        RECT 108.145 176.905 108.475 177.350 ;
        RECT 108.675 176.735 108.930 177.540 ;
        RECT 109.145 177.035 109.375 178.735 ;
        RECT 109.545 178.465 109.840 179.285 ;
        RECT 110.015 178.785 110.315 179.115 ;
        RECT 110.485 178.805 110.760 179.285 ;
        RECT 109.545 176.735 109.840 177.880 ;
        RECT 110.015 177.875 110.185 178.785 ;
        RECT 110.940 178.635 111.235 179.025 ;
        RECT 111.405 178.805 111.660 179.285 ;
        RECT 111.835 178.635 112.095 179.025 ;
        RECT 112.265 178.805 112.545 179.285 ;
        RECT 110.355 178.045 110.705 178.615 ;
        RECT 110.940 178.465 112.590 178.635 ;
        RECT 112.985 178.485 113.265 179.285 ;
        RECT 113.845 178.700 114.125 178.965 ;
        RECT 114.625 178.925 114.955 179.285 ;
        RECT 115.165 178.755 115.335 179.115 ;
        RECT 115.525 178.925 116.300 179.285 ;
        RECT 116.905 178.925 117.235 179.285 ;
        RECT 117.765 178.925 118.105 179.285 ;
        RECT 115.165 178.700 116.175 178.755 ;
        RECT 113.845 178.585 116.175 178.700 ;
        RECT 116.475 178.585 118.065 178.755 ;
        RECT 113.845 178.530 115.335 178.585 ;
        RECT 110.875 178.125 112.015 178.295 ;
        RECT 110.875 177.875 111.045 178.125 ;
        RECT 112.185 177.955 112.590 178.465 ;
        RECT 113.110 178.080 113.525 178.315 ;
        RECT 113.695 178.095 114.220 178.360 ;
        RECT 114.390 178.265 114.785 178.360 ;
        RECT 114.390 178.095 114.845 178.265 ;
        RECT 110.015 177.705 111.045 177.875 ;
        RECT 111.835 177.785 112.590 177.955 ;
        RECT 110.015 176.905 110.325 177.705 ;
        RECT 111.835 177.535 112.095 177.785 ;
        RECT 110.495 176.735 110.805 177.535 ;
        RECT 110.975 177.365 112.095 177.535 ;
        RECT 110.975 176.905 111.235 177.365 ;
        RECT 111.405 176.735 111.660 177.195 ;
        RECT 111.835 176.905 112.095 177.365 ;
        RECT 112.265 176.735 112.550 177.605 ;
        RECT 112.850 177.520 113.105 177.910 ;
        RECT 113.275 177.860 113.525 178.080 ;
        RECT 114.390 177.860 114.565 178.095 ;
        RECT 113.275 177.690 114.565 177.860 ;
        RECT 114.745 177.520 114.925 177.925 ;
        RECT 112.850 177.350 114.925 177.520 ;
        RECT 112.850 176.975 113.180 177.350 ;
        RECT 113.405 176.735 113.735 177.095 ;
        RECT 113.905 176.905 114.075 177.350 ;
        RECT 114.245 176.735 114.575 177.095 ;
        RECT 114.745 177.075 114.925 177.350 ;
        RECT 115.165 177.245 115.335 178.530 ;
        RECT 116.005 178.375 116.175 178.585 ;
        RECT 115.505 177.845 115.815 178.375 ;
        RECT 116.005 178.045 117.410 178.375 ;
        RECT 115.585 177.075 115.755 177.675 ;
        RECT 114.745 176.905 115.755 177.075 ;
        RECT 116.045 176.735 116.295 177.855 ;
        RECT 117.580 177.785 118.065 178.585 ;
        RECT 118.385 178.735 118.555 179.115 ;
        RECT 118.770 178.905 119.100 179.285 ;
        RECT 118.385 178.565 119.100 178.735 ;
        RECT 118.295 178.015 118.650 178.385 ;
        RECT 118.930 178.375 119.100 178.565 ;
        RECT 119.270 178.540 119.525 179.115 ;
        RECT 118.930 178.045 119.185 178.375 ;
        RECT 118.930 177.835 119.100 178.045 ;
        RECT 116.475 177.615 118.065 177.785 ;
        RECT 118.385 177.665 119.100 177.835 ;
        RECT 119.355 177.810 119.525 178.540 ;
        RECT 119.700 178.445 119.960 179.285 ;
        RECT 120.135 178.485 120.445 179.285 ;
        RECT 120.650 178.485 121.345 179.115 ;
        RECT 121.515 178.515 123.185 179.285 ;
        RECT 123.465 178.905 124.635 179.115 ;
        RECT 123.465 178.885 123.795 178.905 ;
        RECT 120.145 178.045 120.480 178.315 ;
        RECT 120.650 177.885 120.820 178.485 ;
        RECT 120.990 178.045 121.325 178.295 ;
        RECT 121.515 177.995 122.265 178.515 ;
        RECT 123.355 178.465 124.215 178.715 ;
        RECT 124.385 178.655 124.635 178.905 ;
        RECT 124.805 178.825 124.975 179.285 ;
        RECT 125.145 178.655 125.485 179.115 ;
        RECT 124.385 178.485 125.485 178.655 ;
        RECT 125.655 178.515 128.245 179.285 ;
        RECT 128.935 178.805 129.215 179.285 ;
        RECT 129.385 178.635 129.645 179.025 ;
        RECT 129.820 178.805 130.075 179.285 ;
        RECT 130.245 178.635 130.540 179.025 ;
        RECT 130.720 178.805 130.995 179.285 ;
        RECT 131.165 178.785 131.465 179.115 ;
        RECT 116.475 177.185 116.725 177.615 ;
        RECT 116.905 176.735 117.235 177.435 ;
        RECT 117.415 177.185 117.585 177.615 ;
        RECT 117.765 176.735 118.095 177.435 ;
        RECT 118.385 176.905 118.555 177.665 ;
        RECT 118.770 176.735 119.100 177.495 ;
        RECT 119.270 176.905 119.525 177.810 ;
        RECT 119.700 176.735 119.960 177.885 ;
        RECT 120.135 176.735 120.415 177.875 ;
        RECT 120.585 176.905 120.915 177.885 ;
        RECT 121.085 176.735 121.345 177.875 ;
        RECT 122.435 177.825 123.185 178.345 ;
        RECT 121.515 176.735 123.185 177.825 ;
        RECT 123.355 177.875 123.635 178.465 ;
        RECT 123.805 178.045 124.555 178.295 ;
        RECT 124.725 178.045 125.485 178.295 ;
        RECT 125.655 177.995 126.865 178.515 ;
        RECT 128.890 178.465 130.540 178.635 ;
        RECT 123.355 177.705 125.055 177.875 ;
        RECT 123.460 176.735 123.715 177.535 ;
        RECT 123.885 176.905 124.215 177.705 ;
        RECT 124.385 176.735 124.555 177.535 ;
        RECT 124.725 176.905 125.055 177.705 ;
        RECT 125.225 176.735 125.485 177.875 ;
        RECT 127.035 177.825 128.245 178.345 ;
        RECT 125.655 176.735 128.245 177.825 ;
        RECT 128.890 177.955 129.295 178.465 ;
        RECT 129.465 178.125 130.605 178.295 ;
        RECT 128.890 177.785 129.645 177.955 ;
        RECT 128.930 176.735 129.215 177.605 ;
        RECT 129.385 177.535 129.645 177.785 ;
        RECT 130.435 177.875 130.605 178.125 ;
        RECT 130.775 178.045 131.125 178.615 ;
        RECT 131.295 177.875 131.465 178.785 ;
        RECT 131.635 178.560 131.925 179.285 ;
        RECT 132.185 178.715 132.355 179.115 ;
        RECT 132.595 178.885 132.925 179.285 ;
        RECT 133.195 178.945 134.600 179.115 ;
        RECT 133.195 178.715 133.365 178.945 ;
        RECT 132.185 178.545 133.365 178.715 ;
        RECT 134.430 178.715 134.600 178.945 ;
        RECT 134.770 178.905 135.100 179.285 ;
        RECT 133.535 178.375 133.725 178.605 ;
        RECT 132.155 178.045 132.340 178.375 ;
        RECT 132.595 178.045 133.070 178.375 ;
        RECT 133.380 178.045 133.725 178.375 ;
        RECT 133.985 178.045 134.180 178.620 ;
        RECT 134.430 178.545 135.125 178.715 ;
        RECT 135.295 178.700 135.605 179.115 ;
        RECT 134.955 178.375 135.125 178.545 ;
        RECT 134.450 178.045 134.785 178.375 ;
        RECT 134.955 178.045 135.265 178.375 ;
        RECT 130.435 177.705 131.465 177.875 ;
        RECT 129.385 177.365 130.505 177.535 ;
        RECT 129.385 176.905 129.645 177.365 ;
        RECT 129.820 176.735 130.075 177.195 ;
        RECT 130.245 176.905 130.505 177.365 ;
        RECT 130.675 176.735 130.985 177.535 ;
        RECT 131.155 176.905 131.465 177.705 ;
        RECT 131.635 176.735 131.925 177.900 ;
        RECT 134.955 177.875 135.125 178.045 ;
        RECT 132.185 177.705 135.125 177.875 ;
        RECT 132.185 176.905 132.355 177.705 ;
        RECT 135.435 177.585 135.605 178.700 ;
        RECT 135.775 178.515 137.445 179.285 ;
        RECT 137.615 178.905 139.000 179.115 ;
        RECT 137.615 178.635 137.905 178.905 ;
        RECT 138.075 178.545 138.500 178.735 ;
        RECT 138.670 178.715 139.000 178.905 ;
        RECT 139.235 178.885 139.565 179.285 ;
        RECT 139.740 178.715 140.070 179.115 ;
        RECT 140.275 178.725 140.445 179.285 ;
        RECT 138.670 178.545 140.070 178.715 ;
        RECT 140.615 178.545 141.125 179.115 ;
        RECT 135.775 177.995 136.525 178.515 ;
        RECT 136.695 177.825 137.445 178.345 ;
        RECT 137.615 178.045 137.890 178.375 ;
        RECT 133.115 177.365 134.675 177.535 ;
        RECT 133.115 176.905 133.365 177.365 ;
        RECT 133.565 176.735 134.235 177.115 ;
        RECT 134.425 176.905 134.675 177.365 ;
        RECT 134.850 176.735 135.095 177.195 ;
        RECT 135.265 176.945 135.605 177.585 ;
        RECT 135.775 176.735 137.445 177.825 ;
        RECT 137.615 176.735 137.905 177.875 ;
        RECT 138.075 177.535 138.245 178.545 ;
        RECT 138.415 177.710 138.770 178.375 ;
        RECT 138.955 177.710 139.230 178.375 ;
        RECT 139.400 178.045 139.745 178.375 ;
        RECT 140.035 178.295 140.205 178.375 ;
        RECT 140.575 178.295 140.765 178.375 ;
        RECT 139.955 178.045 140.205 178.295 ;
        RECT 140.400 178.045 140.765 178.295 ;
        RECT 138.075 177.285 139.030 177.535 ;
        RECT 138.700 177.075 139.030 177.285 ;
        RECT 139.400 177.245 139.725 178.045 ;
        RECT 140.400 177.875 140.570 178.045 ;
        RECT 140.950 177.925 141.125 178.545 ;
        RECT 141.295 178.535 142.505 179.285 ;
        RECT 142.705 178.895 148.175 179.115 ;
        RECT 141.295 177.995 141.815 178.535 ;
        RECT 142.705 178.475 142.955 178.895 ;
        RECT 148.345 178.725 148.675 179.115 ;
        RECT 148.845 178.815 149.015 179.285 ;
        RECT 143.125 178.505 144.715 178.725 ;
        RECT 144.905 178.635 148.675 178.725 ;
        RECT 149.185 178.645 149.515 179.115 ;
        RECT 149.685 178.815 149.855 179.285 ;
        RECT 150.025 178.645 150.355 179.115 ;
        RECT 150.525 178.815 150.695 179.285 ;
        RECT 149.185 178.635 150.355 178.645 ;
        RECT 150.865 178.645 151.195 179.115 ;
        RECT 151.365 178.815 151.535 179.285 ;
        RECT 151.705 178.645 152.035 179.115 ;
        RECT 150.865 178.635 152.035 178.645 ;
        RECT 144.905 178.550 152.035 178.635 ;
        RECT 140.895 177.875 141.125 177.925 ;
        RECT 139.895 177.705 140.570 177.875 ;
        RECT 139.895 177.075 140.065 177.705 ;
        RECT 138.700 176.905 140.065 177.075 ;
        RECT 140.235 176.735 140.525 177.535 ;
        RECT 140.740 176.915 141.125 177.875 ;
        RECT 141.985 177.825 142.505 178.365 ;
        RECT 142.680 178.095 144.340 178.295 ;
        RECT 144.510 177.925 144.715 178.505 ;
        RECT 148.055 178.465 152.035 178.550 ;
        RECT 144.950 178.095 147.095 178.295 ;
        RECT 141.295 176.735 142.505 177.825 ;
        RECT 142.745 176.735 142.995 177.885 ;
        RECT 143.165 177.755 146.755 177.925 ;
        RECT 143.165 176.905 143.415 177.755 ;
        RECT 143.585 176.735 143.835 177.545 ;
        RECT 144.005 177.415 144.715 177.755 ;
        RECT 145.365 177.415 146.415 177.585 ;
        RECT 144.005 176.905 144.255 177.415 ;
        RECT 144.425 176.735 145.195 177.245 ;
        RECT 145.365 176.905 145.615 177.415 ;
        RECT 145.785 176.735 146.035 177.245 ;
        RECT 146.205 177.075 146.415 177.415 ;
        RECT 146.585 177.535 146.755 177.755 ;
        RECT 146.925 177.875 147.095 178.095 ;
        RECT 147.265 178.045 147.875 178.375 ;
        RECT 148.055 177.875 148.385 178.295 ;
        RECT 146.925 177.705 148.385 177.875 ;
        RECT 148.555 177.925 148.885 178.295 ;
        RECT 149.065 178.095 150.475 178.295 ;
        RECT 150.745 178.095 152.165 178.295 ;
        RECT 150.745 177.925 151.010 178.095 ;
        RECT 148.555 177.755 151.010 177.925 ;
        RECT 151.325 177.585 151.575 177.925 ;
        RECT 148.555 177.535 150.315 177.585 ;
        RECT 146.585 177.415 150.315 177.535 ;
        RECT 146.585 177.365 149.475 177.415 ;
        RECT 146.585 177.245 146.875 177.365 ;
        RECT 147.465 177.245 147.675 177.365 ;
        RECT 149.265 177.245 149.475 177.365 ;
        RECT 150.065 177.245 150.315 177.415 ;
        RECT 150.485 177.415 151.575 177.585 ;
        RECT 147.045 177.075 147.295 177.195 ;
        RECT 147.845 177.075 148.175 177.195 ;
        RECT 146.205 176.905 148.175 177.075 ;
        RECT 148.345 176.735 148.595 177.195 ;
        RECT 148.765 177.075 149.095 177.195 ;
        RECT 149.645 177.075 149.895 177.245 ;
        RECT 150.485 177.075 150.735 177.415 ;
        RECT 148.765 176.905 150.735 177.075 ;
        RECT 150.905 176.735 151.155 177.245 ;
        RECT 151.325 176.905 151.575 177.415 ;
        RECT 151.745 176.735 151.995 177.925 ;
        RECT 152.340 177.685 152.675 179.105 ;
        RECT 152.855 178.915 153.600 179.285 ;
        RECT 154.165 178.745 154.420 179.105 ;
        RECT 154.600 178.915 154.930 179.285 ;
        RECT 155.110 178.745 155.335 179.105 ;
        RECT 152.850 178.555 155.335 178.745 ;
        RECT 152.850 177.865 153.075 178.555 ;
        RECT 155.555 178.535 156.765 179.285 ;
        RECT 156.935 178.535 158.145 179.285 ;
        RECT 153.275 178.045 153.555 178.375 ;
        RECT 153.735 178.045 154.310 178.375 ;
        RECT 154.490 178.045 154.925 178.375 ;
        RECT 155.105 178.045 155.375 178.375 ;
        RECT 155.555 177.995 156.075 178.535 ;
        RECT 152.850 177.685 155.345 177.865 ;
        RECT 156.245 177.825 156.765 178.365 ;
        RECT 152.340 176.915 152.605 177.685 ;
        RECT 152.775 176.735 153.105 177.455 ;
        RECT 153.295 177.275 154.485 177.505 ;
        RECT 153.295 176.915 153.555 177.275 ;
        RECT 153.725 176.735 154.055 177.105 ;
        RECT 154.225 176.915 154.485 177.275 ;
        RECT 155.055 176.915 155.345 177.685 ;
        RECT 155.555 176.735 156.765 177.825 ;
        RECT 156.935 177.825 157.455 178.365 ;
        RECT 157.625 177.995 158.145 178.535 ;
        RECT 156.935 176.735 158.145 177.825 ;
        RECT 2.750 176.565 158.230 176.735 ;
        RECT 2.835 175.475 4.045 176.565 ;
        RECT 5.140 175.895 5.395 176.395 ;
        RECT 5.565 176.065 5.895 176.565 ;
        RECT 5.140 175.725 5.890 175.895 ;
        RECT 2.835 174.765 3.355 175.305 ;
        RECT 3.525 174.935 4.045 175.475 ;
        RECT 5.140 174.905 5.490 175.555 ;
        RECT 2.835 174.015 4.045 174.765 ;
        RECT 5.660 174.735 5.890 175.725 ;
        RECT 5.140 174.565 5.890 174.735 ;
        RECT 5.140 174.275 5.395 174.565 ;
        RECT 5.565 174.015 5.895 174.395 ;
        RECT 6.065 174.275 6.235 176.395 ;
        RECT 6.405 175.595 6.730 176.380 ;
        RECT 6.900 176.105 7.150 176.565 ;
        RECT 7.320 176.065 7.570 176.395 ;
        RECT 7.785 176.065 8.465 176.395 ;
        RECT 7.320 175.935 7.490 176.065 ;
        RECT 7.095 175.765 7.490 175.935 ;
        RECT 6.465 174.545 6.925 175.595 ;
        RECT 7.095 174.405 7.265 175.765 ;
        RECT 7.660 175.505 8.125 175.895 ;
        RECT 7.435 174.695 7.785 175.315 ;
        RECT 7.955 174.915 8.125 175.505 ;
        RECT 8.295 175.285 8.465 176.065 ;
        RECT 8.635 175.965 8.805 176.305 ;
        RECT 9.040 176.135 9.370 176.565 ;
        RECT 9.540 175.965 9.710 176.305 ;
        RECT 10.005 176.105 10.375 176.565 ;
        RECT 8.635 175.795 9.710 175.965 ;
        RECT 10.545 175.935 10.715 176.395 ;
        RECT 10.950 176.055 11.820 176.395 ;
        RECT 11.990 176.105 12.240 176.565 ;
        RECT 10.155 175.765 10.715 175.935 ;
        RECT 10.155 175.625 10.325 175.765 ;
        RECT 8.825 175.455 10.325 175.625 ;
        RECT 11.020 175.595 11.480 175.885 ;
        RECT 8.295 175.115 9.985 175.285 ;
        RECT 7.955 174.695 8.310 174.915 ;
        RECT 8.480 174.405 8.650 175.115 ;
        RECT 8.855 174.695 9.645 174.945 ;
        RECT 9.815 174.935 9.985 175.115 ;
        RECT 10.155 174.765 10.325 175.455 ;
        RECT 6.595 174.015 6.925 174.375 ;
        RECT 7.095 174.235 7.590 174.405 ;
        RECT 7.795 174.235 8.650 174.405 ;
        RECT 9.525 174.015 9.855 174.475 ;
        RECT 10.065 174.375 10.325 174.765 ;
        RECT 10.515 175.585 11.480 175.595 ;
        RECT 11.650 175.675 11.820 176.055 ;
        RECT 12.410 176.015 12.580 176.305 ;
        RECT 12.760 176.185 13.090 176.565 ;
        RECT 12.410 175.845 13.210 176.015 ;
        RECT 10.515 175.425 11.190 175.585 ;
        RECT 11.650 175.505 12.870 175.675 ;
        RECT 10.515 174.635 10.725 175.425 ;
        RECT 11.650 175.415 11.820 175.505 ;
        RECT 10.895 174.635 11.245 175.255 ;
        RECT 11.415 175.245 11.820 175.415 ;
        RECT 11.415 174.465 11.585 175.245 ;
        RECT 11.755 174.795 11.975 175.075 ;
        RECT 12.155 174.965 12.695 175.335 ;
        RECT 13.040 175.255 13.210 175.845 ;
        RECT 13.430 175.425 13.735 176.565 ;
        RECT 13.905 175.375 14.160 176.255 ;
        RECT 14.335 175.475 15.545 176.565 ;
        RECT 13.040 175.225 13.780 175.255 ;
        RECT 11.755 174.625 12.285 174.795 ;
        RECT 10.065 174.205 10.415 174.375 ;
        RECT 10.635 174.185 11.585 174.465 ;
        RECT 11.755 174.015 11.945 174.455 ;
        RECT 12.115 174.395 12.285 174.625 ;
        RECT 12.455 174.565 12.695 174.965 ;
        RECT 12.865 174.925 13.780 175.225 ;
        RECT 12.865 174.750 13.190 174.925 ;
        RECT 12.865 174.395 13.185 174.750 ;
        RECT 13.950 174.725 14.160 175.375 ;
        RECT 12.115 174.225 13.185 174.395 ;
        RECT 13.430 174.015 13.735 174.475 ;
        RECT 13.905 174.195 14.160 174.725 ;
        RECT 14.335 174.765 14.855 175.305 ;
        RECT 15.025 174.935 15.545 175.475 ;
        RECT 15.715 175.400 16.005 176.565 ;
        RECT 16.175 175.475 17.385 176.565 ;
        RECT 16.175 174.765 16.695 175.305 ;
        RECT 16.865 174.935 17.385 175.475 ;
        RECT 17.645 175.635 17.815 176.395 ;
        RECT 17.995 175.805 18.325 176.565 ;
        RECT 17.645 175.465 18.310 175.635 ;
        RECT 18.495 175.490 18.765 176.395 ;
        RECT 18.140 175.320 18.310 175.465 ;
        RECT 17.575 174.915 17.905 175.285 ;
        RECT 18.140 174.990 18.425 175.320 ;
        RECT 14.335 174.015 15.545 174.765 ;
        RECT 15.715 174.015 16.005 174.740 ;
        RECT 16.175 174.015 17.385 174.765 ;
        RECT 18.140 174.735 18.310 174.990 ;
        RECT 17.645 174.565 18.310 174.735 ;
        RECT 18.595 174.690 18.765 175.490 ;
        RECT 18.940 176.175 19.275 176.395 ;
        RECT 20.280 176.185 20.635 176.565 ;
        RECT 18.940 175.555 19.195 176.175 ;
        RECT 19.445 176.015 19.675 176.055 ;
        RECT 20.805 176.015 21.055 176.395 ;
        RECT 19.445 175.815 21.055 176.015 ;
        RECT 19.445 175.725 19.630 175.815 ;
        RECT 20.220 175.805 21.055 175.815 ;
        RECT 21.305 175.785 21.555 176.565 ;
        RECT 21.725 175.715 21.985 176.395 ;
        RECT 19.785 175.615 20.115 175.645 ;
        RECT 19.785 175.555 21.585 175.615 ;
        RECT 18.940 175.445 21.645 175.555 ;
        RECT 18.940 175.385 20.115 175.445 ;
        RECT 21.445 175.410 21.645 175.445 ;
        RECT 18.935 175.005 19.425 175.205 ;
        RECT 19.615 175.005 20.090 175.215 ;
        RECT 17.645 174.185 17.815 174.565 ;
        RECT 17.995 174.015 18.325 174.395 ;
        RECT 18.505 174.185 18.765 174.690 ;
        RECT 18.940 174.015 19.395 174.780 ;
        RECT 19.870 174.605 20.090 175.005 ;
        RECT 20.335 175.005 20.665 175.215 ;
        RECT 20.335 174.605 20.545 175.005 ;
        RECT 20.835 174.970 21.245 175.275 ;
        RECT 21.475 174.835 21.645 175.410 ;
        RECT 21.375 174.715 21.645 174.835 ;
        RECT 20.800 174.670 21.645 174.715 ;
        RECT 20.800 174.545 21.555 174.670 ;
        RECT 20.800 174.395 20.970 174.545 ;
        RECT 21.815 174.525 21.985 175.715 ;
        RECT 22.155 175.805 22.670 176.215 ;
        RECT 22.905 175.805 23.075 176.565 ;
        RECT 23.245 176.225 25.275 176.395 ;
        RECT 22.155 174.995 22.495 175.805 ;
        RECT 23.245 175.560 23.415 176.225 ;
        RECT 23.810 175.885 24.935 176.055 ;
        RECT 22.665 175.370 23.415 175.560 ;
        RECT 23.585 175.545 24.595 175.715 ;
        RECT 22.155 174.825 23.385 174.995 ;
        RECT 21.755 174.515 21.985 174.525 ;
        RECT 19.670 174.185 20.970 174.395 ;
        RECT 21.225 174.015 21.555 174.375 ;
        RECT 21.725 174.185 21.985 174.515 ;
        RECT 22.430 174.220 22.675 174.825 ;
        RECT 22.895 174.015 23.405 174.550 ;
        RECT 23.585 174.185 23.775 175.545 ;
        RECT 23.945 175.205 24.220 175.345 ;
        RECT 23.945 175.035 24.225 175.205 ;
        RECT 23.945 174.185 24.220 175.035 ;
        RECT 24.425 174.745 24.595 175.545 ;
        RECT 24.765 174.755 24.935 175.885 ;
        RECT 25.105 175.255 25.275 176.225 ;
        RECT 25.445 175.425 25.615 176.565 ;
        RECT 25.785 175.425 26.120 176.395 ;
        RECT 26.295 176.130 31.640 176.565 ;
        RECT 25.105 174.925 25.300 175.255 ;
        RECT 25.525 174.925 25.780 175.255 ;
        RECT 25.525 174.755 25.695 174.925 ;
        RECT 25.950 174.755 26.120 175.425 ;
        RECT 24.765 174.585 25.695 174.755 ;
        RECT 24.765 174.550 24.940 174.585 ;
        RECT 24.410 174.185 24.940 174.550 ;
        RECT 25.365 174.015 25.695 174.415 ;
        RECT 25.865 174.185 26.120 174.755 ;
        RECT 27.880 174.560 28.220 175.390 ;
        RECT 29.700 174.880 30.050 176.130 ;
        RECT 31.815 175.475 33.025 176.565 ;
        RECT 33.250 175.695 33.535 176.565 ;
        RECT 33.705 175.935 33.965 176.395 ;
        RECT 34.140 176.105 34.395 176.565 ;
        RECT 34.565 175.935 34.825 176.395 ;
        RECT 33.705 175.765 34.825 175.935 ;
        RECT 34.995 175.765 35.305 176.565 ;
        RECT 33.705 175.515 33.965 175.765 ;
        RECT 35.475 175.595 35.785 176.395 ;
        RECT 31.815 174.765 32.335 175.305 ;
        RECT 32.505 174.935 33.025 175.475 ;
        RECT 33.210 175.345 33.965 175.515 ;
        RECT 34.755 175.425 35.785 175.595 ;
        RECT 33.210 174.835 33.615 175.345 ;
        RECT 34.755 175.175 34.925 175.425 ;
        RECT 33.785 175.005 34.925 175.175 ;
        RECT 26.295 174.015 31.640 174.560 ;
        RECT 31.815 174.015 33.025 174.765 ;
        RECT 33.210 174.665 34.860 174.835 ;
        RECT 35.095 174.685 35.445 175.255 ;
        RECT 33.255 174.015 33.535 174.495 ;
        RECT 33.705 174.275 33.965 174.665 ;
        RECT 34.140 174.015 34.395 174.495 ;
        RECT 34.565 174.275 34.860 174.665 ;
        RECT 35.615 174.515 35.785 175.425 ;
        RECT 35.040 174.015 35.315 174.495 ;
        RECT 35.485 174.185 35.785 174.515 ;
        RECT 35.960 175.425 36.295 176.395 ;
        RECT 36.465 175.425 36.635 176.565 ;
        RECT 36.805 176.225 38.835 176.395 ;
        RECT 35.960 174.755 36.130 175.425 ;
        RECT 36.805 175.255 36.975 176.225 ;
        RECT 36.300 174.925 36.555 175.255 ;
        RECT 36.780 174.925 36.975 175.255 ;
        RECT 37.145 175.885 38.270 176.055 ;
        RECT 36.385 174.755 36.555 174.925 ;
        RECT 37.145 174.755 37.315 175.885 ;
        RECT 35.960 174.185 36.215 174.755 ;
        RECT 36.385 174.585 37.315 174.755 ;
        RECT 37.485 175.545 38.495 175.715 ;
        RECT 37.485 174.745 37.655 175.545 ;
        RECT 37.140 174.550 37.315 174.585 ;
        RECT 36.385 174.015 36.715 174.415 ;
        RECT 37.140 174.185 37.670 174.550 ;
        RECT 37.860 174.525 38.135 175.345 ;
        RECT 37.855 174.355 38.135 174.525 ;
        RECT 37.860 174.185 38.135 174.355 ;
        RECT 38.305 174.185 38.495 175.545 ;
        RECT 38.665 175.560 38.835 176.225 ;
        RECT 39.005 175.805 39.175 176.565 ;
        RECT 39.410 175.805 39.925 176.215 ;
        RECT 38.665 175.370 39.415 175.560 ;
        RECT 39.585 174.995 39.925 175.805 ;
        RECT 40.095 175.475 41.305 176.565 ;
        RECT 38.695 174.825 39.925 174.995 ;
        RECT 38.675 174.015 39.185 174.550 ;
        RECT 39.405 174.220 39.650 174.825 ;
        RECT 40.095 174.765 40.615 175.305 ;
        RECT 40.785 174.935 41.305 175.475 ;
        RECT 41.475 175.400 41.765 176.565 ;
        RECT 41.940 175.425 42.275 176.395 ;
        RECT 42.445 175.425 42.615 176.565 ;
        RECT 42.785 176.225 44.815 176.395 ;
        RECT 40.095 174.015 41.305 174.765 ;
        RECT 41.940 174.755 42.110 175.425 ;
        RECT 42.785 175.255 42.955 176.225 ;
        RECT 42.280 174.925 42.535 175.255 ;
        RECT 42.760 174.925 42.955 175.255 ;
        RECT 43.125 175.885 44.250 176.055 ;
        RECT 42.365 174.755 42.535 174.925 ;
        RECT 43.125 174.755 43.295 175.885 ;
        RECT 41.475 174.015 41.765 174.740 ;
        RECT 41.940 174.185 42.195 174.755 ;
        RECT 42.365 174.585 43.295 174.755 ;
        RECT 43.465 175.545 44.475 175.715 ;
        RECT 43.465 174.745 43.635 175.545 ;
        RECT 43.120 174.550 43.295 174.585 ;
        RECT 42.365 174.015 42.695 174.415 ;
        RECT 43.120 174.185 43.650 174.550 ;
        RECT 43.840 174.525 44.115 175.345 ;
        RECT 43.835 174.355 44.115 174.525 ;
        RECT 43.840 174.185 44.115 174.355 ;
        RECT 44.285 174.185 44.475 175.545 ;
        RECT 44.645 175.560 44.815 176.225 ;
        RECT 44.985 175.805 45.155 176.565 ;
        RECT 45.390 175.805 45.905 176.215 ;
        RECT 44.645 175.370 45.395 175.560 ;
        RECT 45.565 174.995 45.905 175.805 ;
        RECT 46.625 175.555 46.795 176.395 ;
        RECT 46.965 176.225 48.135 176.395 ;
        RECT 46.965 175.725 47.295 176.225 ;
        RECT 47.805 176.185 48.135 176.225 ;
        RECT 48.325 176.145 48.680 176.565 ;
        RECT 47.465 175.965 47.695 176.055 ;
        RECT 48.850 175.965 49.100 176.395 ;
        RECT 47.465 175.725 49.100 175.965 ;
        RECT 49.270 175.805 49.600 176.565 ;
        RECT 49.770 175.725 50.025 176.395 ;
        RECT 49.815 175.715 50.025 175.725 ;
        RECT 46.625 175.385 49.685 175.555 ;
        RECT 46.540 175.005 46.890 175.215 ;
        RECT 47.060 175.005 47.505 175.205 ;
        RECT 47.675 175.005 48.150 175.205 ;
        RECT 44.675 174.825 45.905 174.995 ;
        RECT 44.655 174.015 45.165 174.550 ;
        RECT 45.385 174.220 45.630 174.825 ;
        RECT 46.625 174.665 47.690 174.835 ;
        RECT 46.625 174.185 46.795 174.665 ;
        RECT 46.965 174.015 47.295 174.495 ;
        RECT 47.520 174.435 47.690 174.665 ;
        RECT 47.870 174.605 48.150 175.005 ;
        RECT 48.420 175.005 48.750 175.205 ;
        RECT 48.920 175.035 49.295 175.205 ;
        RECT 48.920 175.005 49.285 175.035 ;
        RECT 48.420 174.605 48.705 175.005 ;
        RECT 49.515 174.835 49.685 175.385 ;
        RECT 48.885 174.665 49.685 174.835 ;
        RECT 48.885 174.435 49.055 174.665 ;
        RECT 49.855 174.595 50.025 175.715 ;
        RECT 49.840 174.515 50.025 174.595 ;
        RECT 47.520 174.185 49.055 174.435 ;
        RECT 49.225 174.015 49.555 174.495 ;
        RECT 49.770 174.185 50.025 174.515 ;
        RECT 50.250 175.775 50.785 176.395 ;
        RECT 50.250 174.755 50.565 175.775 ;
        RECT 50.955 175.765 51.285 176.565 ;
        RECT 51.770 175.595 52.160 175.770 ;
        RECT 50.735 175.425 52.160 175.595 ;
        RECT 52.670 175.555 52.970 176.395 ;
        RECT 53.165 175.725 53.415 176.565 ;
        RECT 54.005 175.975 54.810 176.395 ;
        RECT 53.585 175.805 55.150 175.975 ;
        RECT 53.585 175.555 53.755 175.805 ;
        RECT 50.735 174.925 50.905 175.425 ;
        RECT 50.250 174.185 50.865 174.755 ;
        RECT 51.155 174.695 51.420 175.255 ;
        RECT 51.590 174.525 51.760 175.425 ;
        RECT 52.670 175.385 53.755 175.555 ;
        RECT 51.930 174.695 52.285 175.255 ;
        RECT 52.515 174.925 52.845 175.215 ;
        RECT 53.015 174.755 53.185 175.385 ;
        RECT 53.925 175.255 54.245 175.635 ;
        RECT 54.435 175.545 54.810 175.635 ;
        RECT 54.415 175.375 54.810 175.545 ;
        RECT 54.980 175.555 55.150 175.805 ;
        RECT 55.320 175.725 55.650 176.565 ;
        RECT 55.820 175.805 56.485 176.395 ;
        RECT 54.980 175.385 55.900 175.555 ;
        RECT 53.355 175.005 53.685 175.215 ;
        RECT 53.865 175.005 54.245 175.255 ;
        RECT 54.435 175.215 54.810 175.375 ;
        RECT 55.730 175.215 55.900 175.385 ;
        RECT 54.435 175.005 54.920 175.215 ;
        RECT 55.110 175.005 55.560 175.215 ;
        RECT 55.730 175.005 56.065 175.215 ;
        RECT 56.235 174.835 56.485 175.805 ;
        RECT 56.660 175.895 56.915 176.395 ;
        RECT 57.085 176.065 57.415 176.565 ;
        RECT 56.660 175.725 57.410 175.895 ;
        RECT 56.660 174.905 57.010 175.555 ;
        RECT 52.675 174.575 53.185 174.755 ;
        RECT 53.590 174.665 55.290 174.835 ;
        RECT 53.590 174.575 53.975 174.665 ;
        RECT 51.035 174.015 51.250 174.525 ;
        RECT 51.480 174.195 51.760 174.525 ;
        RECT 51.940 174.015 52.180 174.525 ;
        RECT 52.675 174.185 53.005 174.575 ;
        RECT 53.175 174.235 54.360 174.405 ;
        RECT 54.620 174.015 54.790 174.485 ;
        RECT 54.960 174.200 55.290 174.665 ;
        RECT 55.460 174.015 55.630 174.835 ;
        RECT 55.800 174.195 56.485 174.835 ;
        RECT 57.180 174.735 57.410 175.725 ;
        RECT 56.660 174.565 57.410 174.735 ;
        RECT 56.660 174.275 56.915 174.565 ;
        RECT 57.085 174.015 57.415 174.395 ;
        RECT 57.585 174.275 57.755 176.395 ;
        RECT 57.925 175.595 58.250 176.380 ;
        RECT 58.420 176.105 58.670 176.565 ;
        RECT 58.840 176.065 59.090 176.395 ;
        RECT 59.305 176.065 59.985 176.395 ;
        RECT 58.840 175.935 59.010 176.065 ;
        RECT 58.615 175.765 59.010 175.935 ;
        RECT 57.985 174.545 58.445 175.595 ;
        RECT 58.615 174.405 58.785 175.765 ;
        RECT 59.180 175.505 59.645 175.895 ;
        RECT 58.955 174.695 59.305 175.315 ;
        RECT 59.475 174.915 59.645 175.505 ;
        RECT 59.815 175.285 59.985 176.065 ;
        RECT 60.155 175.965 60.325 176.305 ;
        RECT 60.560 176.135 60.890 176.565 ;
        RECT 61.060 175.965 61.230 176.305 ;
        RECT 61.525 176.105 61.895 176.565 ;
        RECT 60.155 175.795 61.230 175.965 ;
        RECT 62.065 175.935 62.235 176.395 ;
        RECT 62.470 176.055 63.340 176.395 ;
        RECT 63.510 176.105 63.760 176.565 ;
        RECT 61.675 175.765 62.235 175.935 ;
        RECT 61.675 175.625 61.845 175.765 ;
        RECT 60.345 175.455 61.845 175.625 ;
        RECT 62.540 175.595 63.000 175.885 ;
        RECT 59.815 175.115 61.505 175.285 ;
        RECT 59.475 174.695 59.830 174.915 ;
        RECT 60.000 174.405 60.170 175.115 ;
        RECT 60.375 174.695 61.165 174.945 ;
        RECT 61.335 174.935 61.505 175.115 ;
        RECT 61.675 174.765 61.845 175.455 ;
        RECT 58.115 174.015 58.445 174.375 ;
        RECT 58.615 174.235 59.110 174.405 ;
        RECT 59.315 174.235 60.170 174.405 ;
        RECT 61.045 174.015 61.375 174.475 ;
        RECT 61.585 174.375 61.845 174.765 ;
        RECT 62.035 175.585 63.000 175.595 ;
        RECT 63.170 175.675 63.340 176.055 ;
        RECT 63.930 176.015 64.100 176.305 ;
        RECT 64.280 176.185 64.610 176.565 ;
        RECT 63.930 175.845 64.730 176.015 ;
        RECT 62.035 175.425 62.710 175.585 ;
        RECT 63.170 175.505 64.390 175.675 ;
        RECT 62.035 174.635 62.245 175.425 ;
        RECT 63.170 175.415 63.340 175.505 ;
        RECT 62.415 174.635 62.765 175.255 ;
        RECT 62.935 175.245 63.340 175.415 ;
        RECT 62.935 174.465 63.105 175.245 ;
        RECT 63.275 174.795 63.495 175.075 ;
        RECT 63.675 174.965 64.215 175.335 ;
        RECT 64.560 175.255 64.730 175.845 ;
        RECT 64.950 175.425 65.255 176.565 ;
        RECT 65.425 175.375 65.675 176.255 ;
        RECT 65.845 175.425 66.095 176.565 ;
        RECT 67.235 175.400 67.525 176.565 ;
        RECT 67.695 175.475 68.905 176.565 ;
        RECT 69.075 175.800 69.540 176.395 ;
        RECT 69.710 176.000 69.910 176.395 ;
        RECT 70.080 176.170 70.410 176.565 ;
        RECT 70.580 176.000 70.750 176.395 ;
        RECT 69.710 175.800 70.750 176.000 ;
        RECT 70.920 175.630 71.170 176.395 ;
        RECT 71.340 176.000 71.670 176.395 ;
        RECT 72.320 176.170 72.650 176.565 ;
        RECT 72.820 176.000 72.990 176.395 ;
        RECT 71.340 175.800 72.990 176.000 ;
        RECT 64.560 175.225 65.300 175.255 ;
        RECT 63.275 174.625 63.805 174.795 ;
        RECT 61.585 174.205 61.935 174.375 ;
        RECT 62.155 174.185 63.105 174.465 ;
        RECT 63.275 174.015 63.465 174.455 ;
        RECT 63.635 174.395 63.805 174.625 ;
        RECT 63.975 174.565 64.215 174.965 ;
        RECT 64.385 174.925 65.300 175.225 ;
        RECT 64.385 174.750 64.710 174.925 ;
        RECT 64.385 174.395 64.705 174.750 ;
        RECT 65.470 174.725 65.675 175.375 ;
        RECT 63.635 174.225 64.705 174.395 ;
        RECT 64.950 174.015 65.255 174.475 ;
        RECT 65.425 174.195 65.675 174.725 ;
        RECT 65.845 174.015 66.095 174.770 ;
        RECT 67.695 174.765 68.215 175.305 ;
        RECT 68.385 174.935 68.905 175.475 ;
        RECT 69.075 175.460 70.750 175.630 ;
        RECT 70.920 175.460 72.110 175.630 ;
        RECT 69.075 174.985 69.790 175.460 ;
        RECT 70.460 175.290 70.750 175.460 ;
        RECT 69.960 174.985 70.290 175.290 ;
        RECT 70.460 174.985 71.165 175.290 ;
        RECT 71.335 174.985 71.665 175.290 ;
        RECT 72.280 175.285 72.650 175.625 ;
        RECT 71.855 174.985 72.650 175.285 ;
        RECT 72.820 175.220 72.990 175.800 ;
        RECT 73.180 175.390 73.510 176.565 ;
        RECT 73.680 175.595 73.865 176.395 ;
        RECT 74.035 175.765 74.365 176.565 ;
        RECT 74.535 175.595 74.750 176.395 ;
        RECT 74.920 175.765 75.345 176.565 ;
        RECT 75.605 175.595 75.775 176.395 ;
        RECT 76.065 175.935 76.315 176.355 ;
        RECT 76.505 176.105 76.835 176.565 ;
        RECT 77.045 175.935 77.295 176.355 ;
        RECT 76.005 175.765 77.295 175.935 ;
        RECT 77.465 175.765 77.715 176.565 ;
        RECT 77.885 175.935 78.055 176.395 ;
        RECT 78.265 176.105 78.515 176.565 ;
        RECT 77.885 175.765 78.560 175.935 ;
        RECT 73.680 175.390 75.345 175.595 ;
        RECT 75.605 175.425 78.095 175.595 ;
        RECT 74.655 175.375 75.345 175.390 ;
        RECT 72.820 174.985 74.525 175.220 ;
        RECT 72.820 174.815 72.990 174.985 ;
        RECT 74.695 174.815 75.345 175.375 ;
        RECT 67.235 174.015 67.525 174.740 ;
        RECT 67.695 174.015 68.905 174.765 ;
        RECT 69.075 174.565 72.050 174.815 ;
        RECT 72.220 174.565 72.990 174.815 ;
        RECT 69.075 174.185 69.490 174.565 ;
        RECT 69.660 174.015 69.990 174.375 ;
        RECT 70.160 174.185 70.330 174.565 ;
        RECT 70.500 174.015 70.830 174.375 ;
        RECT 71.000 174.185 71.170 174.565 ;
        RECT 71.860 174.395 72.050 174.565 ;
        RECT 71.340 174.015 71.670 174.375 ;
        RECT 71.860 174.185 72.990 174.395 ;
        RECT 73.180 174.015 73.495 174.815 ;
        RECT 73.665 174.645 75.345 174.815 ;
        RECT 75.560 174.685 75.755 175.255 ;
        RECT 73.665 174.585 74.750 174.645 ;
        RECT 73.665 174.185 73.865 174.585 ;
        RECT 74.035 174.015 74.365 174.415 ;
        RECT 74.535 174.185 74.750 174.585 ;
        RECT 74.920 174.015 75.345 174.475 ;
        RECT 75.515 174.015 75.775 174.495 ;
        RECT 75.945 174.435 76.115 175.425 ;
        RECT 76.295 174.800 76.465 175.255 ;
        RECT 76.855 175.175 77.025 175.190 ;
        RECT 76.695 175.005 77.025 175.175 ;
        RECT 76.295 174.630 76.685 174.800 ;
        RECT 75.945 174.265 76.275 174.435 ;
        RECT 76.475 174.345 76.685 174.630 ;
        RECT 76.855 174.795 77.025 175.005 ;
        RECT 77.255 174.925 77.585 175.255 ;
        RECT 77.925 175.175 78.095 175.425 ;
        RECT 77.765 175.005 78.095 175.175 ;
        RECT 76.855 174.625 77.120 174.795 ;
        RECT 77.380 174.690 77.585 174.925 ;
        RECT 78.305 174.815 78.560 175.765 ;
        RECT 78.740 175.895 78.995 176.395 ;
        RECT 79.165 176.065 79.495 176.565 ;
        RECT 78.740 175.725 79.490 175.895 ;
        RECT 78.740 174.905 79.090 175.555 ;
        RECT 76.950 174.525 77.120 174.625 ;
        RECT 77.885 174.645 78.560 174.815 ;
        RECT 79.260 174.735 79.490 175.725 ;
        RECT 76.950 174.355 77.125 174.525 ;
        RECT 77.465 174.395 77.635 174.475 ;
        RECT 76.950 174.330 77.120 174.355 ;
        RECT 75.945 174.185 76.190 174.265 ;
        RECT 77.365 174.015 77.695 174.395 ;
        RECT 77.885 174.185 78.055 174.645 ;
        RECT 78.740 174.565 79.490 174.735 ;
        RECT 78.305 174.015 78.560 174.475 ;
        RECT 78.740 174.275 78.995 174.565 ;
        RECT 79.165 174.015 79.495 174.395 ;
        RECT 79.665 174.275 79.835 176.395 ;
        RECT 80.005 175.595 80.330 176.380 ;
        RECT 80.500 176.105 80.750 176.565 ;
        RECT 80.920 176.065 81.170 176.395 ;
        RECT 81.385 176.065 82.065 176.395 ;
        RECT 80.920 175.935 81.090 176.065 ;
        RECT 80.695 175.765 81.090 175.935 ;
        RECT 80.065 174.545 80.525 175.595 ;
        RECT 80.695 174.405 80.865 175.765 ;
        RECT 81.260 175.505 81.725 175.895 ;
        RECT 81.035 174.695 81.385 175.315 ;
        RECT 81.555 174.915 81.725 175.505 ;
        RECT 81.895 175.285 82.065 176.065 ;
        RECT 82.235 175.965 82.405 176.305 ;
        RECT 82.640 176.135 82.970 176.565 ;
        RECT 83.140 175.965 83.310 176.305 ;
        RECT 83.605 176.105 83.975 176.565 ;
        RECT 82.235 175.795 83.310 175.965 ;
        RECT 84.145 175.935 84.315 176.395 ;
        RECT 84.550 176.055 85.420 176.395 ;
        RECT 85.590 176.105 85.840 176.565 ;
        RECT 83.755 175.765 84.315 175.935 ;
        RECT 83.755 175.625 83.925 175.765 ;
        RECT 82.425 175.455 83.925 175.625 ;
        RECT 84.620 175.595 85.080 175.885 ;
        RECT 81.895 175.115 83.585 175.285 ;
        RECT 81.555 174.695 81.910 174.915 ;
        RECT 82.080 174.405 82.250 175.115 ;
        RECT 82.455 174.695 83.245 174.945 ;
        RECT 83.415 174.935 83.585 175.115 ;
        RECT 83.755 174.765 83.925 175.455 ;
        RECT 80.195 174.015 80.525 174.375 ;
        RECT 80.695 174.235 81.190 174.405 ;
        RECT 81.395 174.235 82.250 174.405 ;
        RECT 83.125 174.015 83.455 174.475 ;
        RECT 83.665 174.375 83.925 174.765 ;
        RECT 84.115 175.585 85.080 175.595 ;
        RECT 85.250 175.675 85.420 176.055 ;
        RECT 86.010 176.015 86.180 176.305 ;
        RECT 86.360 176.185 86.690 176.565 ;
        RECT 86.010 175.845 86.810 176.015 ;
        RECT 84.115 175.425 84.790 175.585 ;
        RECT 85.250 175.505 86.470 175.675 ;
        RECT 84.115 174.635 84.325 175.425 ;
        RECT 85.250 175.415 85.420 175.505 ;
        RECT 84.495 174.635 84.845 175.255 ;
        RECT 85.015 175.245 85.420 175.415 ;
        RECT 85.015 174.465 85.185 175.245 ;
        RECT 85.355 174.795 85.575 175.075 ;
        RECT 85.755 174.965 86.295 175.335 ;
        RECT 86.640 175.255 86.810 175.845 ;
        RECT 87.030 175.425 87.335 176.565 ;
        RECT 87.505 175.375 87.760 176.255 ;
        RECT 86.640 175.225 87.380 175.255 ;
        RECT 85.355 174.625 85.885 174.795 ;
        RECT 83.665 174.205 84.015 174.375 ;
        RECT 84.235 174.185 85.185 174.465 ;
        RECT 85.355 174.015 85.545 174.455 ;
        RECT 85.715 174.395 85.885 174.625 ;
        RECT 86.055 174.565 86.295 174.965 ;
        RECT 86.465 174.925 87.380 175.225 ;
        RECT 86.465 174.750 86.790 174.925 ;
        RECT 86.465 174.395 86.785 174.750 ;
        RECT 87.550 174.725 87.760 175.375 ;
        RECT 85.715 174.225 86.785 174.395 ;
        RECT 87.030 174.015 87.335 174.475 ;
        RECT 87.505 174.195 87.760 174.725 ;
        RECT 87.935 175.425 88.320 176.395 ;
        RECT 88.490 176.105 88.815 176.565 ;
        RECT 89.335 175.935 89.615 176.395 ;
        RECT 88.490 175.715 89.615 175.935 ;
        RECT 87.935 174.755 88.215 175.425 ;
        RECT 88.490 175.255 88.940 175.715 ;
        RECT 89.805 175.545 90.205 176.395 ;
        RECT 90.605 176.105 90.875 176.565 ;
        RECT 91.045 175.935 91.330 176.395 ;
        RECT 88.385 174.925 88.940 175.255 ;
        RECT 89.110 174.985 90.205 175.545 ;
        RECT 88.490 174.815 88.940 174.925 ;
        RECT 87.935 174.185 88.320 174.755 ;
        RECT 88.490 174.645 89.615 174.815 ;
        RECT 88.490 174.015 88.815 174.475 ;
        RECT 89.335 174.185 89.615 174.645 ;
        RECT 89.805 174.185 90.205 174.985 ;
        RECT 90.375 175.715 91.330 175.935 ;
        RECT 90.375 174.815 90.585 175.715 ;
        RECT 90.755 174.985 91.445 175.545 ;
        RECT 91.615 175.425 91.895 176.565 ;
        RECT 92.065 175.415 92.395 176.395 ;
        RECT 92.565 175.425 92.825 176.565 ;
        RECT 91.625 174.985 91.960 175.255 ;
        RECT 92.130 174.815 92.300 175.415 ;
        RECT 92.995 175.400 93.285 176.565 ;
        RECT 93.460 175.695 93.725 176.395 ;
        RECT 93.895 175.865 94.225 176.565 ;
        RECT 94.395 175.695 95.065 176.395 ;
        RECT 95.570 175.865 96.000 176.565 ;
        RECT 96.180 176.005 96.370 176.395 ;
        RECT 96.540 176.185 96.870 176.565 ;
        RECT 97.135 176.060 97.765 176.565 ;
        RECT 96.180 175.835 96.910 176.005 ;
        RECT 93.460 175.440 96.035 175.695 ;
        RECT 92.470 175.005 92.805 175.255 ;
        RECT 93.455 174.925 93.730 175.255 ;
        RECT 90.375 174.645 91.330 174.815 ;
        RECT 90.605 174.015 90.875 174.475 ;
        RECT 91.045 174.185 91.330 174.645 ;
        RECT 91.615 174.015 91.925 174.815 ;
        RECT 92.130 174.185 92.825 174.815 ;
        RECT 93.900 174.755 94.080 175.440 ;
        RECT 95.865 175.255 96.035 175.440 ;
        RECT 94.250 174.925 94.610 175.255 ;
        RECT 94.900 175.205 95.190 175.255 ;
        RECT 94.895 175.035 95.190 175.205 ;
        RECT 94.900 174.925 95.190 175.035 ;
        RECT 95.360 174.925 95.695 175.255 ;
        RECT 95.865 174.925 96.545 175.255 ;
        RECT 92.995 174.015 93.285 174.740 ;
        RECT 93.465 174.355 94.080 174.755 ;
        RECT 94.250 174.565 95.520 174.755 ;
        RECT 96.715 174.715 96.910 175.835 ;
        RECT 97.150 175.525 97.405 175.890 ;
        RECT 97.575 175.885 97.765 176.060 ;
        RECT 97.945 176.055 98.420 176.395 ;
        RECT 97.575 175.695 97.905 175.885 ;
        RECT 98.130 175.525 98.380 175.820 ;
        RECT 98.605 175.720 98.820 176.565 ;
        RECT 99.020 175.725 99.295 176.395 ;
        RECT 97.150 175.355 98.940 175.525 ;
        RECT 99.125 175.375 99.295 175.725 ;
        RECT 99.465 175.555 99.725 176.565 ;
        RECT 96.090 174.545 96.910 174.715 ;
        RECT 97.135 174.695 97.520 175.175 ;
        RECT 93.465 174.185 93.800 174.355 ;
        RECT 94.760 174.015 95.095 174.395 ;
        RECT 95.685 174.015 95.920 174.455 ;
        RECT 96.090 174.185 96.420 174.545 ;
        RECT 97.690 174.500 97.945 175.355 ;
        RECT 96.590 174.015 96.920 174.375 ;
        RECT 97.155 174.235 97.945 174.500 ;
        RECT 98.115 174.680 98.525 175.175 ;
        RECT 98.710 174.925 98.940 175.355 ;
        RECT 99.110 174.855 99.725 175.375 ;
        RECT 99.895 175.360 100.185 176.565 ;
        RECT 100.355 175.425 100.630 176.395 ;
        RECT 100.840 175.765 101.120 176.565 ;
        RECT 101.290 176.055 102.485 176.345 ;
        RECT 102.660 176.055 104.315 176.345 ;
        RECT 101.300 175.715 102.465 175.885 ;
        RECT 101.300 175.595 101.470 175.715 ;
        RECT 100.800 175.425 101.470 175.595 ;
        RECT 98.115 174.235 98.345 174.680 ;
        RECT 99.110 174.645 99.280 174.855 ;
        RECT 98.525 174.015 98.855 174.510 ;
        RECT 99.030 174.185 99.280 174.645 ;
        RECT 99.450 174.015 99.725 174.675 ;
        RECT 99.895 174.015 100.185 174.845 ;
        RECT 100.355 174.690 100.525 175.425 ;
        RECT 100.800 175.255 100.970 175.425 ;
        RECT 101.740 175.255 101.965 175.545 ;
        RECT 102.135 175.425 102.465 175.715 ;
        RECT 102.660 175.715 104.250 175.885 ;
        RECT 104.485 175.765 104.765 176.565 ;
        RECT 102.660 175.425 102.980 175.715 ;
        RECT 104.080 175.595 104.250 175.715 ;
        RECT 100.695 174.925 100.970 175.255 ;
        RECT 101.140 174.925 101.965 175.255 ;
        RECT 102.135 174.925 102.485 175.255 ;
        RECT 100.800 174.755 100.970 174.925 ;
        RECT 100.355 174.345 100.630 174.690 ;
        RECT 100.800 174.585 102.465 174.755 ;
        RECT 102.660 174.685 103.010 175.255 ;
        RECT 103.180 174.925 103.890 175.545 ;
        RECT 104.080 175.425 104.805 175.595 ;
        RECT 104.975 175.425 105.245 176.395 ;
        RECT 105.415 176.055 106.605 176.345 ;
        RECT 105.435 175.715 106.605 175.885 ;
        RECT 106.775 175.765 107.055 176.565 ;
        RECT 105.435 175.425 105.760 175.715 ;
        RECT 106.435 175.595 106.605 175.715 ;
        RECT 104.635 175.255 104.805 175.425 ;
        RECT 104.060 174.925 104.465 175.255 ;
        RECT 104.635 174.925 104.905 175.255 ;
        RECT 104.635 174.755 104.805 174.925 ;
        RECT 100.820 174.015 101.200 174.415 ;
        RECT 101.370 174.235 101.540 174.585 ;
        RECT 101.710 174.015 102.040 174.415 ;
        RECT 102.210 174.235 102.465 174.585 ;
        RECT 103.195 174.585 104.805 174.755 ;
        RECT 105.075 174.690 105.245 175.425 ;
        RECT 105.930 175.255 106.125 175.545 ;
        RECT 106.435 175.425 107.095 175.595 ;
        RECT 107.265 175.425 107.540 176.395 ;
        RECT 107.725 175.425 108.055 176.565 ;
        RECT 108.585 175.595 108.915 176.380 ;
        RECT 108.235 175.425 108.915 175.595 ;
        RECT 106.925 175.255 107.095 175.425 ;
        RECT 105.415 174.925 105.760 175.255 ;
        RECT 105.930 174.925 106.755 175.255 ;
        RECT 106.925 174.925 107.200 175.255 ;
        RECT 106.925 174.755 107.095 174.925 ;
        RECT 102.665 174.015 102.995 174.515 ;
        RECT 103.195 174.235 103.365 174.585 ;
        RECT 103.565 174.015 103.895 174.415 ;
        RECT 104.065 174.235 104.235 174.585 ;
        RECT 104.405 174.015 104.785 174.415 ;
        RECT 104.975 174.345 105.245 174.690 ;
        RECT 105.430 174.585 107.095 174.755 ;
        RECT 107.370 174.690 107.540 175.425 ;
        RECT 107.715 175.005 108.065 175.255 ;
        RECT 108.235 174.825 108.405 175.425 ;
        RECT 110.020 175.415 110.280 176.565 ;
        RECT 110.455 175.490 110.710 176.395 ;
        RECT 110.880 175.805 111.210 176.565 ;
        RECT 111.425 175.635 111.595 176.395 ;
        RECT 108.575 175.005 108.925 175.255 ;
        RECT 105.430 174.235 105.685 174.585 ;
        RECT 105.855 174.015 106.185 174.415 ;
        RECT 106.355 174.235 106.525 174.585 ;
        RECT 106.695 174.015 107.075 174.415 ;
        RECT 107.265 174.345 107.540 174.690 ;
        RECT 107.725 174.015 107.995 174.825 ;
        RECT 108.165 174.185 108.495 174.825 ;
        RECT 108.665 174.015 108.905 174.825 ;
        RECT 110.020 174.015 110.280 174.855 ;
        RECT 110.455 174.760 110.625 175.490 ;
        RECT 110.880 175.465 111.595 175.635 ;
        RECT 112.775 175.595 113.085 176.395 ;
        RECT 113.255 175.765 113.565 176.565 ;
        RECT 113.735 175.935 113.995 176.395 ;
        RECT 114.165 176.105 114.420 176.565 ;
        RECT 114.595 175.935 114.855 176.395 ;
        RECT 113.735 175.765 114.855 175.935 ;
        RECT 110.880 175.255 111.050 175.465 ;
        RECT 112.775 175.425 113.805 175.595 ;
        RECT 110.795 174.925 111.050 175.255 ;
        RECT 110.455 174.185 110.710 174.760 ;
        RECT 110.880 174.735 111.050 174.925 ;
        RECT 111.330 174.915 111.685 175.285 ;
        RECT 110.880 174.565 111.595 174.735 ;
        RECT 110.880 174.015 111.210 174.395 ;
        RECT 111.425 174.185 111.595 174.565 ;
        RECT 112.775 174.515 112.945 175.425 ;
        RECT 113.115 174.685 113.465 175.255 ;
        RECT 113.635 175.175 113.805 175.425 ;
        RECT 114.595 175.515 114.855 175.765 ;
        RECT 115.025 175.695 115.310 176.565 ;
        RECT 115.535 176.010 116.140 176.565 ;
        RECT 116.315 176.055 116.795 176.395 ;
        RECT 116.965 176.020 117.220 176.565 ;
        RECT 115.535 175.910 116.150 176.010 ;
        RECT 115.965 175.885 116.150 175.910 ;
        RECT 114.595 175.345 115.350 175.515 ;
        RECT 113.635 175.005 114.775 175.175 ;
        RECT 114.945 174.835 115.350 175.345 ;
        RECT 115.535 175.290 115.795 175.740 ;
        RECT 115.965 175.640 116.295 175.885 ;
        RECT 116.465 175.565 117.220 175.815 ;
        RECT 117.390 175.695 117.665 176.395 ;
        RECT 116.450 175.530 117.220 175.565 ;
        RECT 116.435 175.520 117.220 175.530 ;
        RECT 116.430 175.505 117.325 175.520 ;
        RECT 116.410 175.490 117.325 175.505 ;
        RECT 116.390 175.480 117.325 175.490 ;
        RECT 116.365 175.470 117.325 175.480 ;
        RECT 116.295 175.440 117.325 175.470 ;
        RECT 116.275 175.410 117.325 175.440 ;
        RECT 116.255 175.380 117.325 175.410 ;
        RECT 116.225 175.355 117.325 175.380 ;
        RECT 116.190 175.320 117.325 175.355 ;
        RECT 116.160 175.315 117.325 175.320 ;
        RECT 116.160 175.310 116.550 175.315 ;
        RECT 116.160 175.300 116.525 175.310 ;
        RECT 116.160 175.295 116.510 175.300 ;
        RECT 116.160 175.290 116.495 175.295 ;
        RECT 115.535 175.285 116.495 175.290 ;
        RECT 115.535 175.275 116.485 175.285 ;
        RECT 115.535 175.270 116.475 175.275 ;
        RECT 115.535 175.260 116.465 175.270 ;
        RECT 115.535 175.250 116.460 175.260 ;
        RECT 115.535 175.245 116.455 175.250 ;
        RECT 115.535 175.230 116.445 175.245 ;
        RECT 115.535 175.215 116.440 175.230 ;
        RECT 115.535 175.190 116.430 175.215 ;
        RECT 115.535 175.120 116.425 175.190 ;
        RECT 113.700 174.665 115.350 174.835 ;
        RECT 112.775 174.185 113.075 174.515 ;
        RECT 113.245 174.015 113.520 174.495 ;
        RECT 113.700 174.275 113.995 174.665 ;
        RECT 114.165 174.015 114.420 174.495 ;
        RECT 114.595 174.275 114.855 174.665 ;
        RECT 115.535 174.565 116.085 174.950 ;
        RECT 115.025 174.015 115.305 174.495 ;
        RECT 116.255 174.395 116.425 175.120 ;
        RECT 115.535 174.225 116.425 174.395 ;
        RECT 116.595 174.720 116.925 175.145 ;
        RECT 117.095 174.920 117.325 175.315 ;
        RECT 116.595 174.235 116.815 174.720 ;
        RECT 117.495 174.665 117.665 175.695 ;
        RECT 118.755 175.400 119.045 176.565 ;
        RECT 119.215 175.595 119.525 176.395 ;
        RECT 119.695 175.765 120.005 176.565 ;
        RECT 120.175 175.935 120.435 176.395 ;
        RECT 120.605 176.105 120.860 176.565 ;
        RECT 121.035 175.935 121.295 176.395 ;
        RECT 120.175 175.765 121.295 175.935 ;
        RECT 119.215 175.425 120.245 175.595 ;
        RECT 116.985 174.015 117.235 174.555 ;
        RECT 117.405 174.185 117.665 174.665 ;
        RECT 118.755 174.015 119.045 174.740 ;
        RECT 119.215 174.515 119.385 175.425 ;
        RECT 119.555 174.685 119.905 175.255 ;
        RECT 120.075 175.175 120.245 175.425 ;
        RECT 121.035 175.515 121.295 175.765 ;
        RECT 121.465 175.695 121.750 176.565 ;
        RECT 121.035 175.345 121.790 175.515 ;
        RECT 121.980 175.415 122.240 176.565 ;
        RECT 122.415 175.490 122.670 176.395 ;
        RECT 122.840 175.805 123.170 176.565 ;
        RECT 123.385 175.635 123.555 176.395 ;
        RECT 123.815 176.060 124.445 176.565 ;
        RECT 120.075 175.005 121.215 175.175 ;
        RECT 121.385 174.835 121.790 175.345 ;
        RECT 120.140 174.665 121.790 174.835 ;
        RECT 119.215 174.185 119.515 174.515 ;
        RECT 119.685 174.015 119.960 174.495 ;
        RECT 120.140 174.275 120.435 174.665 ;
        RECT 120.605 174.015 120.860 174.495 ;
        RECT 121.035 174.275 121.295 174.665 ;
        RECT 121.465 174.015 121.745 174.495 ;
        RECT 121.980 174.015 122.240 174.855 ;
        RECT 122.415 174.760 122.585 175.490 ;
        RECT 122.840 175.465 123.555 175.635 ;
        RECT 123.830 175.525 124.085 175.890 ;
        RECT 124.255 175.885 124.445 176.060 ;
        RECT 124.625 176.055 125.100 176.395 ;
        RECT 124.255 175.695 124.585 175.885 ;
        RECT 124.810 175.525 125.060 175.820 ;
        RECT 125.285 175.720 125.500 176.565 ;
        RECT 125.700 175.725 125.975 176.395 ;
        RECT 122.840 175.255 123.010 175.465 ;
        RECT 123.830 175.355 125.620 175.525 ;
        RECT 125.805 175.375 125.975 175.725 ;
        RECT 126.145 175.555 126.405 176.565 ;
        RECT 126.595 175.675 126.855 176.385 ;
        RECT 127.025 175.855 127.355 176.565 ;
        RECT 127.525 175.675 127.755 176.385 ;
        RECT 126.595 175.435 127.755 175.675 ;
        RECT 127.935 175.655 128.205 176.385 ;
        RECT 128.385 175.835 128.725 176.565 ;
        RECT 127.935 175.435 128.705 175.655 ;
        RECT 122.755 174.925 123.010 175.255 ;
        RECT 122.415 174.185 122.670 174.760 ;
        RECT 122.840 174.735 123.010 174.925 ;
        RECT 123.290 174.915 123.645 175.285 ;
        RECT 122.840 174.565 123.555 174.735 ;
        RECT 123.815 174.695 124.200 175.175 ;
        RECT 122.840 174.015 123.170 174.395 ;
        RECT 123.385 174.185 123.555 174.565 ;
        RECT 124.370 174.500 124.625 175.355 ;
        RECT 123.835 174.235 124.625 174.500 ;
        RECT 124.795 174.680 125.205 175.175 ;
        RECT 125.390 174.925 125.620 175.355 ;
        RECT 125.790 174.855 126.405 175.375 ;
        RECT 126.585 174.925 126.885 175.255 ;
        RECT 127.065 174.945 127.590 175.255 ;
        RECT 127.770 174.945 128.235 175.255 ;
        RECT 124.795 174.235 125.025 174.680 ;
        RECT 125.790 174.645 125.960 174.855 ;
        RECT 125.205 174.015 125.535 174.510 ;
        RECT 125.710 174.185 125.960 174.645 ;
        RECT 126.130 174.015 126.405 174.675 ;
        RECT 126.595 174.015 126.885 174.745 ;
        RECT 127.065 174.305 127.295 174.945 ;
        RECT 128.415 174.765 128.705 175.435 ;
        RECT 127.475 174.565 128.705 174.765 ;
        RECT 127.475 174.195 127.785 174.565 ;
        RECT 127.965 174.015 128.635 174.385 ;
        RECT 128.895 174.195 129.155 176.385 ;
        RECT 129.335 175.475 131.005 176.565 ;
        RECT 131.820 175.765 131.990 176.565 ;
        RECT 132.160 175.935 132.490 176.395 ;
        RECT 132.660 176.105 132.830 176.565 ;
        RECT 133.000 175.935 133.330 176.395 ;
        RECT 132.160 175.765 133.330 175.935 ;
        RECT 133.540 175.765 133.710 176.565 ;
        RECT 132.160 175.595 132.490 175.765 ;
        RECT 134.255 175.595 134.615 176.395 ;
        RECT 129.335 174.785 130.085 175.305 ;
        RECT 130.255 174.955 131.005 175.475 ;
        RECT 131.635 175.425 132.490 175.595 ;
        RECT 133.155 175.425 134.615 175.595 ;
        RECT 134.855 175.475 136.065 176.565 ;
        RECT 131.635 174.835 131.980 175.425 ;
        RECT 133.155 175.175 133.360 175.425 ;
        RECT 132.150 175.005 133.360 175.175 ;
        RECT 133.530 174.925 133.905 175.255 ;
        RECT 129.335 174.015 131.005 174.785 ;
        RECT 131.635 174.665 133.330 174.835 ;
        RECT 134.075 174.755 134.255 175.425 ;
        RECT 131.820 174.015 131.990 174.495 ;
        RECT 132.160 174.195 132.490 174.665 ;
        RECT 132.660 174.015 132.830 174.495 ;
        RECT 133.000 174.195 133.330 174.665 ;
        RECT 133.540 174.015 133.710 174.755 ;
        RECT 133.925 174.220 134.255 174.755 ;
        RECT 134.425 174.695 134.680 175.255 ;
        RECT 134.855 174.765 135.375 175.305 ;
        RECT 135.545 174.935 136.065 175.475 ;
        RECT 136.240 175.425 136.560 176.565 ;
        RECT 136.740 175.255 136.935 176.305 ;
        RECT 137.115 175.715 137.445 176.395 ;
        RECT 137.645 175.765 137.900 176.565 ;
        RECT 137.115 175.435 137.465 175.715 ;
        RECT 138.545 175.615 138.820 176.385 ;
        RECT 138.990 175.955 139.320 176.385 ;
        RECT 139.490 176.125 139.685 176.565 ;
        RECT 139.865 175.955 140.195 176.385 ;
        RECT 138.990 175.785 140.195 175.955 ;
        RECT 136.300 175.205 136.560 175.255 ;
        RECT 136.295 175.035 136.560 175.205 ;
        RECT 136.300 174.925 136.560 175.035 ;
        RECT 136.740 174.925 137.125 175.255 ;
        RECT 137.295 175.055 137.465 175.435 ;
        RECT 137.655 175.225 137.900 175.585 ;
        RECT 138.545 175.425 139.130 175.615 ;
        RECT 139.300 175.455 140.195 175.785 ;
        RECT 140.375 175.475 143.885 176.565 ;
        RECT 137.295 174.885 137.815 175.055 ;
        RECT 134.425 174.015 134.665 174.525 ;
        RECT 134.855 174.015 136.065 174.765 ;
        RECT 136.240 174.545 137.455 174.715 ;
        RECT 136.240 174.195 136.530 174.545 ;
        RECT 136.725 174.015 137.055 174.375 ;
        RECT 137.225 174.240 137.455 174.545 ;
        RECT 137.645 174.320 137.815 174.885 ;
        RECT 138.545 174.605 138.785 175.255 ;
        RECT 138.955 174.755 139.130 175.425 ;
        RECT 139.300 174.925 139.715 175.255 ;
        RECT 139.895 174.925 140.190 175.255 ;
        RECT 138.955 174.575 139.285 174.755 ;
        RECT 138.560 174.015 138.890 174.405 ;
        RECT 139.060 174.195 139.285 174.575 ;
        RECT 139.485 174.305 139.715 174.925 ;
        RECT 140.375 174.785 142.025 175.305 ;
        RECT 142.195 174.955 143.885 175.475 ;
        RECT 144.515 175.400 144.805 176.565 ;
        RECT 144.975 175.475 148.485 176.565 ;
        RECT 149.575 176.055 150.765 176.345 ;
        RECT 144.975 174.785 146.625 175.305 ;
        RECT 146.795 174.955 148.485 175.475 ;
        RECT 149.595 175.715 150.765 175.885 ;
        RECT 150.935 175.765 151.215 176.565 ;
        RECT 149.595 175.425 149.920 175.715 ;
        RECT 150.595 175.595 150.765 175.715 ;
        RECT 150.090 175.255 150.285 175.545 ;
        RECT 150.595 175.425 151.255 175.595 ;
        RECT 151.425 175.425 151.700 176.395 ;
        RECT 151.875 175.475 155.385 176.565 ;
        RECT 155.555 175.475 156.765 176.565 ;
        RECT 151.085 175.255 151.255 175.425 ;
        RECT 149.575 174.925 149.920 175.255 ;
        RECT 150.090 174.925 150.915 175.255 ;
        RECT 151.085 174.925 151.360 175.255 ;
        RECT 139.895 174.015 140.195 174.745 ;
        RECT 140.375 174.015 143.885 174.785 ;
        RECT 144.515 174.015 144.805 174.740 ;
        RECT 144.975 174.015 148.485 174.785 ;
        RECT 151.085 174.755 151.255 174.925 ;
        RECT 149.590 174.585 151.255 174.755 ;
        RECT 151.530 174.690 151.700 175.425 ;
        RECT 149.590 174.235 149.845 174.585 ;
        RECT 150.015 174.015 150.345 174.415 ;
        RECT 150.515 174.235 150.685 174.585 ;
        RECT 150.855 174.015 151.235 174.415 ;
        RECT 151.425 174.345 151.700 174.690 ;
        RECT 151.875 174.785 153.525 175.305 ;
        RECT 153.695 174.955 155.385 175.475 ;
        RECT 151.875 174.015 155.385 174.785 ;
        RECT 155.555 174.765 156.075 175.305 ;
        RECT 156.245 174.935 156.765 175.475 ;
        RECT 156.935 175.475 158.145 176.565 ;
        RECT 156.935 174.935 157.455 175.475 ;
        RECT 157.625 174.765 158.145 175.305 ;
        RECT 155.555 174.015 156.765 174.765 ;
        RECT 156.935 174.015 158.145 174.765 ;
        RECT 2.750 173.845 158.230 174.015 ;
        RECT 2.835 173.095 4.045 173.845 ;
        RECT 2.835 172.555 3.355 173.095 ;
        RECT 4.215 173.075 6.805 173.845 ;
        RECT 7.435 173.170 7.695 173.675 ;
        RECT 7.875 173.465 8.205 173.845 ;
        RECT 8.385 173.295 8.555 173.675 ;
        RECT 3.525 172.385 4.045 172.925 ;
        RECT 4.215 172.555 5.425 173.075 ;
        RECT 5.595 172.385 6.805 172.905 ;
        RECT 2.835 171.295 4.045 172.385 ;
        RECT 4.215 171.295 6.805 172.385 ;
        RECT 7.435 172.370 7.605 173.170 ;
        RECT 7.890 173.125 8.555 173.295 ;
        RECT 7.890 172.870 8.060 173.125 ;
        RECT 8.815 173.095 10.025 173.845 ;
        RECT 10.200 173.105 10.455 173.675 ;
        RECT 10.625 173.445 10.955 173.845 ;
        RECT 11.380 173.310 11.910 173.675 ;
        RECT 11.380 173.275 11.555 173.310 ;
        RECT 10.625 173.105 11.555 173.275 ;
        RECT 12.100 173.165 12.375 173.675 ;
        RECT 7.775 172.540 8.060 172.870 ;
        RECT 8.295 172.575 8.625 172.945 ;
        RECT 8.815 172.555 9.335 173.095 ;
        RECT 7.890 172.395 8.060 172.540 ;
        RECT 7.435 171.465 7.705 172.370 ;
        RECT 7.890 172.225 8.555 172.395 ;
        RECT 9.505 172.385 10.025 172.925 ;
        RECT 7.875 171.295 8.205 172.055 ;
        RECT 8.385 171.465 8.555 172.225 ;
        RECT 8.815 171.295 10.025 172.385 ;
        RECT 10.200 172.435 10.370 173.105 ;
        RECT 10.625 172.935 10.795 173.105 ;
        RECT 10.540 172.605 10.795 172.935 ;
        RECT 11.020 172.605 11.215 172.935 ;
        RECT 10.200 171.465 10.535 172.435 ;
        RECT 10.705 171.295 10.875 172.435 ;
        RECT 11.045 171.635 11.215 172.605 ;
        RECT 11.385 171.975 11.555 173.105 ;
        RECT 11.725 172.315 11.895 173.115 ;
        RECT 12.095 172.995 12.375 173.165 ;
        RECT 12.100 172.515 12.375 172.995 ;
        RECT 12.545 172.315 12.735 173.675 ;
        RECT 12.915 173.310 13.425 173.845 ;
        RECT 13.645 173.035 13.890 173.640 ;
        RECT 14.335 173.075 17.845 173.845 ;
        RECT 18.940 173.080 19.395 173.845 ;
        RECT 19.670 173.465 20.970 173.675 ;
        RECT 21.225 173.485 21.555 173.845 ;
        RECT 20.800 173.315 20.970 173.465 ;
        RECT 21.725 173.345 21.985 173.675 ;
        RECT 12.935 172.865 14.165 173.035 ;
        RECT 11.725 172.145 12.735 172.315 ;
        RECT 12.905 172.300 13.655 172.490 ;
        RECT 11.385 171.805 12.510 171.975 ;
        RECT 12.905 171.635 13.075 172.300 ;
        RECT 13.825 172.055 14.165 172.865 ;
        RECT 14.335 172.555 15.985 173.075 ;
        RECT 16.155 172.385 17.845 172.905 ;
        RECT 19.870 172.855 20.090 173.255 ;
        RECT 18.935 172.655 19.425 172.855 ;
        RECT 19.615 172.645 20.090 172.855 ;
        RECT 20.335 172.855 20.545 173.255 ;
        RECT 20.800 173.190 21.555 173.315 ;
        RECT 20.800 173.145 21.645 173.190 ;
        RECT 21.375 173.025 21.645 173.145 ;
        RECT 20.335 172.645 20.665 172.855 ;
        RECT 20.835 172.585 21.245 172.890 ;
        RECT 11.045 171.465 13.075 171.635 ;
        RECT 13.245 171.295 13.415 172.055 ;
        RECT 13.650 171.645 14.165 172.055 ;
        RECT 14.335 171.295 17.845 172.385 ;
        RECT 18.940 172.415 20.115 172.475 ;
        RECT 21.475 172.450 21.645 173.025 ;
        RECT 21.445 172.415 21.645 172.450 ;
        RECT 18.940 172.305 21.645 172.415 ;
        RECT 18.940 171.685 19.195 172.305 ;
        RECT 19.785 172.245 21.585 172.305 ;
        RECT 19.785 172.215 20.115 172.245 ;
        RECT 21.815 172.145 21.985 173.345 ;
        RECT 22.430 173.035 22.675 173.640 ;
        RECT 22.895 173.310 23.405 173.845 ;
        RECT 19.445 172.045 19.630 172.135 ;
        RECT 20.220 172.045 21.055 172.055 ;
        RECT 19.445 171.845 21.055 172.045 ;
        RECT 19.445 171.805 19.675 171.845 ;
        RECT 18.940 171.465 19.275 171.685 ;
        RECT 20.280 171.295 20.635 171.675 ;
        RECT 20.805 171.465 21.055 171.845 ;
        RECT 21.305 171.295 21.555 172.075 ;
        RECT 21.725 171.465 21.985 172.145 ;
        RECT 22.155 172.865 23.385 173.035 ;
        RECT 22.155 172.055 22.495 172.865 ;
        RECT 22.665 172.300 23.415 172.490 ;
        RECT 22.155 171.645 22.670 172.055 ;
        RECT 22.905 171.295 23.075 172.055 ;
        RECT 23.245 171.635 23.415 172.300 ;
        RECT 23.585 172.315 23.775 173.675 ;
        RECT 23.945 173.505 24.220 173.675 ;
        RECT 23.945 173.335 24.225 173.505 ;
        RECT 23.945 172.515 24.220 173.335 ;
        RECT 24.410 173.310 24.940 173.675 ;
        RECT 25.365 173.445 25.695 173.845 ;
        RECT 24.765 173.275 24.940 173.310 ;
        RECT 24.425 172.315 24.595 173.115 ;
        RECT 23.585 172.145 24.595 172.315 ;
        RECT 24.765 173.105 25.695 173.275 ;
        RECT 25.865 173.105 26.120 173.675 ;
        RECT 24.765 171.975 24.935 173.105 ;
        RECT 25.525 172.935 25.695 173.105 ;
        RECT 23.810 171.805 24.935 171.975 ;
        RECT 25.105 172.605 25.300 172.935 ;
        RECT 25.525 172.605 25.780 172.935 ;
        RECT 25.105 171.635 25.275 172.605 ;
        RECT 25.950 172.435 26.120 173.105 ;
        RECT 26.295 173.075 27.965 173.845 ;
        RECT 28.595 173.120 28.885 173.845 ;
        RECT 29.515 173.170 29.775 173.675 ;
        RECT 29.955 173.465 30.285 173.845 ;
        RECT 30.465 173.295 30.635 173.675 ;
        RECT 26.295 172.555 27.045 173.075 ;
        RECT 23.245 171.465 25.275 171.635 ;
        RECT 25.445 171.295 25.615 172.435 ;
        RECT 25.785 171.465 26.120 172.435 ;
        RECT 27.215 172.385 27.965 172.905 ;
        RECT 26.295 171.295 27.965 172.385 ;
        RECT 28.595 171.295 28.885 172.460 ;
        RECT 29.515 172.370 29.685 173.170 ;
        RECT 29.970 173.125 30.635 173.295 ;
        RECT 29.970 172.870 30.140 173.125 ;
        RECT 30.900 173.105 31.155 173.675 ;
        RECT 31.325 173.445 31.655 173.845 ;
        RECT 32.080 173.310 32.610 173.675 ;
        RECT 32.080 173.275 32.255 173.310 ;
        RECT 31.325 173.105 32.255 173.275 ;
        RECT 29.855 172.540 30.140 172.870 ;
        RECT 30.375 172.575 30.705 172.945 ;
        RECT 29.970 172.395 30.140 172.540 ;
        RECT 30.900 172.435 31.070 173.105 ;
        RECT 31.325 172.935 31.495 173.105 ;
        RECT 31.240 172.605 31.495 172.935 ;
        RECT 31.720 172.605 31.915 172.935 ;
        RECT 29.515 171.465 29.785 172.370 ;
        RECT 29.970 172.225 30.635 172.395 ;
        RECT 29.955 171.295 30.285 172.055 ;
        RECT 30.465 171.465 30.635 172.225 ;
        RECT 30.900 171.465 31.235 172.435 ;
        RECT 31.405 171.295 31.575 172.435 ;
        RECT 31.745 171.635 31.915 172.605 ;
        RECT 32.085 171.975 32.255 173.105 ;
        RECT 32.425 172.315 32.595 173.115 ;
        RECT 32.800 172.825 33.075 173.675 ;
        RECT 32.795 172.655 33.075 172.825 ;
        RECT 32.800 172.515 33.075 172.655 ;
        RECT 33.245 172.315 33.435 173.675 ;
        RECT 33.615 173.310 34.125 173.845 ;
        RECT 34.345 173.035 34.590 173.640 ;
        RECT 35.035 173.075 36.705 173.845 ;
        RECT 37.340 173.295 37.595 173.585 ;
        RECT 37.765 173.465 38.095 173.845 ;
        RECT 37.340 173.125 38.090 173.295 ;
        RECT 33.635 172.865 34.865 173.035 ;
        RECT 32.425 172.145 33.435 172.315 ;
        RECT 33.605 172.300 34.355 172.490 ;
        RECT 32.085 171.805 33.210 171.975 ;
        RECT 33.605 171.635 33.775 172.300 ;
        RECT 34.525 172.055 34.865 172.865 ;
        RECT 35.035 172.555 35.785 173.075 ;
        RECT 35.955 172.385 36.705 172.905 ;
        RECT 31.745 171.465 33.775 171.635 ;
        RECT 33.945 171.295 34.115 172.055 ;
        RECT 34.350 171.645 34.865 172.055 ;
        RECT 35.035 171.295 36.705 172.385 ;
        RECT 37.340 172.305 37.690 172.955 ;
        RECT 37.860 172.135 38.090 173.125 ;
        RECT 37.340 171.965 38.090 172.135 ;
        RECT 37.340 171.465 37.595 171.965 ;
        RECT 37.765 171.295 38.095 171.795 ;
        RECT 38.265 171.465 38.435 173.585 ;
        RECT 38.795 173.485 39.125 173.845 ;
        RECT 39.295 173.455 39.790 173.625 ;
        RECT 39.995 173.455 40.850 173.625 ;
        RECT 38.665 172.265 39.125 173.315 ;
        RECT 38.605 171.480 38.930 172.265 ;
        RECT 39.295 172.095 39.465 173.455 ;
        RECT 39.635 172.545 39.985 173.165 ;
        RECT 40.155 172.945 40.510 173.165 ;
        RECT 40.155 172.355 40.325 172.945 ;
        RECT 40.680 172.745 40.850 173.455 ;
        RECT 41.725 173.385 42.055 173.845 ;
        RECT 42.265 173.485 42.615 173.655 ;
        RECT 41.055 172.915 41.845 173.165 ;
        RECT 42.265 173.095 42.525 173.485 ;
        RECT 42.835 173.395 43.785 173.675 ;
        RECT 43.955 173.405 44.145 173.845 ;
        RECT 44.315 173.465 45.385 173.635 ;
        RECT 42.015 172.745 42.185 172.925 ;
        RECT 39.295 171.925 39.690 172.095 ;
        RECT 39.860 171.965 40.325 172.355 ;
        RECT 40.495 172.575 42.185 172.745 ;
        RECT 39.520 171.795 39.690 171.925 ;
        RECT 40.495 171.795 40.665 172.575 ;
        RECT 42.355 172.405 42.525 173.095 ;
        RECT 41.025 172.235 42.525 172.405 ;
        RECT 42.715 172.435 42.925 173.225 ;
        RECT 43.095 172.605 43.445 173.225 ;
        RECT 43.615 172.615 43.785 173.395 ;
        RECT 44.315 173.235 44.485 173.465 ;
        RECT 43.955 173.065 44.485 173.235 ;
        RECT 43.955 172.785 44.175 173.065 ;
        RECT 44.655 172.895 44.895 173.295 ;
        RECT 43.615 172.445 44.020 172.615 ;
        RECT 44.355 172.525 44.895 172.895 ;
        RECT 45.065 173.110 45.385 173.465 ;
        RECT 45.630 173.385 45.935 173.845 ;
        RECT 46.105 173.135 46.360 173.665 ;
        RECT 45.065 172.935 45.390 173.110 ;
        RECT 45.065 172.635 45.980 172.935 ;
        RECT 45.240 172.605 45.980 172.635 ;
        RECT 42.715 172.275 43.390 172.435 ;
        RECT 43.850 172.355 44.020 172.445 ;
        RECT 42.715 172.265 43.680 172.275 ;
        RECT 42.355 172.095 42.525 172.235 ;
        RECT 39.100 171.295 39.350 171.755 ;
        RECT 39.520 171.465 39.770 171.795 ;
        RECT 39.985 171.465 40.665 171.795 ;
        RECT 40.835 171.895 41.910 172.065 ;
        RECT 42.355 171.925 42.915 172.095 ;
        RECT 43.220 171.975 43.680 172.265 ;
        RECT 43.850 172.185 45.070 172.355 ;
        RECT 40.835 171.555 41.005 171.895 ;
        RECT 41.240 171.295 41.570 171.725 ;
        RECT 41.740 171.555 41.910 171.895 ;
        RECT 42.205 171.295 42.575 171.755 ;
        RECT 42.745 171.465 42.915 171.925 ;
        RECT 43.850 171.805 44.020 172.185 ;
        RECT 45.240 172.015 45.410 172.605 ;
        RECT 46.150 172.485 46.360 173.135 ;
        RECT 43.150 171.465 44.020 171.805 ;
        RECT 44.610 171.845 45.410 172.015 ;
        RECT 44.190 171.295 44.440 171.755 ;
        RECT 44.610 171.555 44.780 171.845 ;
        RECT 44.960 171.295 45.290 171.675 ;
        RECT 45.630 171.295 45.935 172.435 ;
        RECT 46.105 171.605 46.360 172.485 ;
        RECT 46.535 173.345 46.835 173.675 ;
        RECT 47.005 173.365 47.280 173.845 ;
        RECT 46.535 172.435 46.705 173.345 ;
        RECT 47.460 173.195 47.755 173.585 ;
        RECT 47.925 173.365 48.180 173.845 ;
        RECT 48.355 173.195 48.615 173.585 ;
        RECT 48.785 173.365 49.065 173.845 ;
        RECT 46.875 172.605 47.225 173.175 ;
        RECT 47.460 173.025 49.110 173.195 ;
        RECT 49.305 173.035 49.575 173.845 ;
        RECT 49.745 173.035 50.075 173.675 ;
        RECT 50.245 173.035 50.485 173.845 ;
        RECT 50.765 173.195 50.935 173.675 ;
        RECT 51.105 173.365 51.435 173.845 ;
        RECT 51.660 173.425 53.195 173.675 ;
        RECT 51.660 173.195 51.830 173.425 ;
        RECT 47.395 172.685 48.535 172.855 ;
        RECT 47.395 172.435 47.565 172.685 ;
        RECT 48.705 172.515 49.110 173.025 ;
        RECT 49.295 172.605 49.645 172.855 ;
        RECT 46.535 172.265 47.565 172.435 ;
        RECT 48.355 172.345 49.110 172.515 ;
        RECT 49.815 172.435 49.985 173.035 ;
        RECT 50.765 173.025 51.830 173.195 ;
        RECT 52.010 172.855 52.290 173.255 ;
        RECT 50.155 172.605 50.505 172.855 ;
        RECT 50.680 172.645 51.030 172.855 ;
        RECT 51.200 172.655 51.645 172.855 ;
        RECT 51.815 172.655 52.290 172.855 ;
        RECT 52.560 172.855 52.845 173.255 ;
        RECT 53.025 173.195 53.195 173.425 ;
        RECT 53.365 173.365 53.695 173.845 ;
        RECT 53.910 173.345 54.165 173.675 ;
        RECT 53.980 173.265 54.165 173.345 ;
        RECT 53.025 173.025 53.825 173.195 ;
        RECT 52.560 172.655 52.890 172.855 ;
        RECT 53.060 172.655 53.425 172.855 ;
        RECT 53.655 172.475 53.825 173.025 ;
        RECT 46.535 171.465 46.845 172.265 ;
        RECT 48.355 172.095 48.615 172.345 ;
        RECT 47.015 171.295 47.325 172.095 ;
        RECT 47.495 171.925 48.615 172.095 ;
        RECT 47.495 171.465 47.755 171.925 ;
        RECT 47.925 171.295 48.180 171.755 ;
        RECT 48.355 171.465 48.615 171.925 ;
        RECT 48.785 171.295 49.070 172.165 ;
        RECT 49.305 171.295 49.635 172.435 ;
        RECT 49.815 172.265 50.495 172.435 ;
        RECT 50.165 171.480 50.495 172.265 ;
        RECT 50.765 172.305 53.825 172.475 ;
        RECT 50.765 171.465 50.935 172.305 ;
        RECT 53.995 172.135 54.165 173.265 ;
        RECT 54.355 173.120 54.645 173.845 ;
        RECT 55.895 173.285 56.225 173.675 ;
        RECT 56.395 173.455 57.580 173.625 ;
        RECT 57.840 173.375 58.010 173.845 ;
        RECT 55.895 173.105 56.405 173.285 ;
        RECT 55.735 172.645 56.065 172.935 ;
        RECT 56.235 172.475 56.405 173.105 ;
        RECT 56.810 173.195 57.195 173.285 ;
        RECT 58.180 173.195 58.510 173.660 ;
        RECT 56.810 173.025 58.510 173.195 ;
        RECT 58.680 173.025 58.850 173.845 ;
        RECT 59.020 173.025 59.705 173.665 ;
        RECT 60.910 173.215 61.195 173.675 ;
        RECT 61.365 173.385 61.635 173.845 ;
        RECT 60.910 173.045 61.865 173.215 ;
        RECT 56.575 172.645 56.905 172.855 ;
        RECT 57.085 172.605 57.465 172.855 ;
        RECT 57.655 172.825 58.140 172.855 ;
        RECT 57.635 172.655 58.140 172.825 ;
        RECT 51.105 171.635 51.435 172.135 ;
        RECT 51.605 171.895 53.240 172.135 ;
        RECT 51.605 171.805 51.835 171.895 ;
        RECT 51.945 171.635 52.275 171.675 ;
        RECT 51.105 171.465 52.275 171.635 ;
        RECT 52.465 171.295 52.820 171.715 ;
        RECT 52.990 171.465 53.240 171.895 ;
        RECT 53.410 171.295 53.740 172.055 ;
        RECT 53.910 171.465 54.165 172.135 ;
        RECT 54.355 171.295 54.645 172.460 ;
        RECT 55.890 172.305 56.975 172.475 ;
        RECT 55.890 171.465 56.190 172.305 ;
        RECT 56.385 171.295 56.635 172.135 ;
        RECT 56.805 172.055 56.975 172.305 ;
        RECT 57.145 172.225 57.465 172.605 ;
        RECT 57.655 172.645 58.140 172.655 ;
        RECT 58.330 172.645 58.780 172.855 ;
        RECT 58.950 172.645 59.285 172.855 ;
        RECT 57.655 172.225 58.030 172.645 ;
        RECT 58.950 172.475 59.120 172.645 ;
        RECT 58.200 172.305 59.120 172.475 ;
        RECT 58.200 172.055 58.370 172.305 ;
        RECT 56.805 171.885 58.370 172.055 ;
        RECT 57.225 171.465 58.030 171.885 ;
        RECT 58.540 171.295 58.870 172.135 ;
        RECT 59.455 172.055 59.705 173.025 ;
        RECT 60.795 172.315 61.485 172.875 ;
        RECT 61.655 172.145 61.865 173.045 ;
        RECT 59.040 171.465 59.705 172.055 ;
        RECT 60.910 171.925 61.865 172.145 ;
        RECT 62.035 172.875 62.435 173.675 ;
        RECT 62.625 173.215 62.905 173.675 ;
        RECT 63.425 173.385 63.750 173.845 ;
        RECT 62.625 173.045 63.750 173.215 ;
        RECT 63.920 173.105 64.305 173.675 ;
        RECT 63.300 172.935 63.750 173.045 ;
        RECT 62.035 172.315 63.130 172.875 ;
        RECT 63.300 172.605 63.855 172.935 ;
        RECT 60.910 171.465 61.195 171.925 ;
        RECT 61.365 171.295 61.635 171.755 ;
        RECT 62.035 171.465 62.435 172.315 ;
        RECT 63.300 172.145 63.750 172.605 ;
        RECT 64.025 172.435 64.305 173.105 ;
        RECT 64.590 173.215 64.875 173.675 ;
        RECT 65.045 173.385 65.315 173.845 ;
        RECT 64.590 173.045 65.545 173.215 ;
        RECT 62.625 171.925 63.750 172.145 ;
        RECT 62.625 171.465 62.905 171.925 ;
        RECT 63.425 171.295 63.750 171.755 ;
        RECT 63.920 171.465 64.305 172.435 ;
        RECT 64.475 172.315 65.165 172.875 ;
        RECT 65.335 172.145 65.545 173.045 ;
        RECT 64.590 171.925 65.545 172.145 ;
        RECT 65.715 172.875 66.115 173.675 ;
        RECT 66.305 173.215 66.585 173.675 ;
        RECT 67.105 173.385 67.430 173.845 ;
        RECT 66.305 173.045 67.430 173.215 ;
        RECT 67.600 173.105 67.985 173.675 ;
        RECT 68.190 173.345 68.440 173.845 ;
        RECT 68.770 173.275 68.940 173.625 ;
        RECT 69.140 173.445 69.470 173.845 ;
        RECT 69.640 173.275 69.810 173.625 ;
        RECT 70.030 173.445 70.410 173.845 ;
        RECT 66.980 172.935 67.430 173.045 ;
        RECT 65.715 172.315 66.810 172.875 ;
        RECT 66.980 172.605 67.535 172.935 ;
        RECT 64.590 171.465 64.875 171.925 ;
        RECT 65.045 171.295 65.315 171.755 ;
        RECT 65.715 171.465 66.115 172.315 ;
        RECT 66.980 172.145 67.430 172.605 ;
        RECT 67.705 172.435 67.985 173.105 ;
        RECT 68.155 172.605 68.440 173.175 ;
        RECT 68.610 173.105 70.420 173.275 ;
        RECT 68.610 172.435 68.780 173.105 ;
        RECT 66.305 171.925 67.430 172.145 ;
        RECT 66.305 171.465 66.585 171.925 ;
        RECT 67.105 171.295 67.430 171.755 ;
        RECT 67.600 171.465 67.985 172.435 ;
        RECT 68.185 172.265 68.780 172.435 ;
        RECT 68.950 172.310 69.120 172.935 ;
        RECT 69.350 172.480 69.680 172.935 ;
        RECT 68.185 171.480 68.520 172.265 ;
        RECT 68.950 171.555 69.300 172.310 ;
        RECT 69.470 172.145 69.680 172.480 ;
        RECT 69.910 172.485 70.080 172.935 ;
        RECT 70.250 172.855 70.420 173.105 ;
        RECT 70.590 173.205 70.840 173.675 ;
        RECT 71.010 173.375 71.180 173.845 ;
        RECT 71.350 173.205 71.680 173.675 ;
        RECT 71.850 173.375 72.020 173.845 ;
        RECT 73.220 173.215 73.555 173.675 ;
        RECT 73.725 173.385 73.895 173.845 ;
        RECT 74.065 173.215 74.395 173.675 ;
        RECT 74.565 173.385 74.735 173.845 ;
        RECT 74.905 173.465 76.915 173.675 ;
        RECT 77.815 173.465 78.705 173.635 ;
        RECT 74.905 173.215 75.155 173.465 ;
        RECT 70.590 173.025 72.125 173.205 ;
        RECT 73.220 173.025 75.155 173.215 ;
        RECT 75.325 173.125 76.495 173.295 ;
        RECT 70.250 172.685 71.710 172.855 ;
        RECT 69.910 172.315 70.345 172.485 ;
        RECT 71.880 172.475 72.125 173.025 ;
        RECT 75.325 172.855 75.575 173.125 ;
        RECT 76.665 173.045 76.915 173.465 ;
        RECT 77.815 172.910 78.365 173.295 ;
        RECT 73.240 172.605 74.860 172.855 ;
        RECT 70.550 172.305 72.125 172.475 ;
        RECT 75.040 172.435 75.575 172.855 ;
        RECT 75.745 172.605 77.185 172.855 ;
        RECT 78.535 172.740 78.705 173.465 ;
        RECT 77.815 172.670 78.705 172.740 ;
        RECT 78.875 173.165 79.095 173.625 ;
        RECT 79.265 173.305 79.515 173.845 ;
        RECT 79.685 173.195 79.945 173.675 ;
        RECT 78.875 173.140 79.125 173.165 ;
        RECT 78.875 172.715 79.205 173.140 ;
        RECT 77.815 172.645 78.710 172.670 ;
        RECT 77.815 172.630 78.720 172.645 ;
        RECT 77.815 172.615 78.725 172.630 ;
        RECT 77.815 172.610 78.735 172.615 ;
        RECT 77.815 172.600 78.740 172.610 ;
        RECT 77.815 172.590 78.745 172.600 ;
        RECT 77.815 172.585 78.755 172.590 ;
        RECT 77.815 172.575 78.765 172.585 ;
        RECT 77.815 172.570 78.775 172.575 ;
        RECT 69.470 171.555 69.790 172.145 ;
        RECT 70.075 171.295 70.325 172.135 ;
        RECT 70.550 171.465 70.800 172.305 ;
        RECT 70.970 171.295 71.220 172.135 ;
        RECT 71.390 171.465 71.640 172.305 ;
        RECT 71.810 171.295 72.060 172.135 ;
        RECT 73.220 171.295 73.475 172.435 ;
        RECT 73.645 172.265 76.495 172.435 ;
        RECT 73.645 171.465 73.975 172.265 ;
        RECT 74.145 171.295 74.315 172.095 ;
        RECT 74.485 171.465 74.815 172.265 ;
        RECT 74.985 171.295 75.155 172.095 ;
        RECT 75.325 171.465 75.655 172.265 ;
        RECT 75.825 171.295 75.995 172.095 ;
        RECT 76.165 171.465 76.495 172.265 ;
        RECT 77.815 172.120 78.075 172.570 ;
        RECT 78.440 172.565 78.775 172.570 ;
        RECT 78.440 172.560 78.790 172.565 ;
        RECT 78.440 172.550 78.805 172.560 ;
        RECT 78.440 172.545 78.830 172.550 ;
        RECT 79.375 172.545 79.605 172.940 ;
        RECT 78.440 172.540 79.605 172.545 ;
        RECT 78.470 172.505 79.605 172.540 ;
        RECT 78.505 172.480 79.605 172.505 ;
        RECT 78.535 172.450 79.605 172.480 ;
        RECT 78.555 172.420 79.605 172.450 ;
        RECT 78.575 172.390 79.605 172.420 ;
        RECT 78.645 172.380 79.605 172.390 ;
        RECT 78.670 172.370 79.605 172.380 ;
        RECT 78.690 172.355 79.605 172.370 ;
        RECT 78.710 172.340 79.605 172.355 ;
        RECT 78.715 172.330 79.500 172.340 ;
        RECT 78.730 172.295 79.500 172.330 ;
        RECT 76.665 171.295 76.915 172.095 ;
        RECT 78.245 171.975 78.575 172.220 ;
        RECT 78.745 172.045 79.500 172.295 ;
        RECT 79.775 172.165 79.945 173.195 ;
        RECT 80.115 173.120 80.405 173.845 ;
        RECT 80.575 173.365 80.835 173.845 ;
        RECT 81.005 173.595 81.250 173.675 ;
        RECT 81.005 173.425 81.335 173.595 ;
        RECT 80.620 172.605 80.815 173.175 ;
        RECT 78.245 171.950 78.430 171.975 ;
        RECT 77.815 171.850 78.430 171.950 ;
        RECT 77.815 171.295 78.420 171.850 ;
        RECT 78.595 171.465 79.075 171.805 ;
        RECT 79.245 171.295 79.500 171.840 ;
        RECT 79.670 171.465 79.945 172.165 ;
        RECT 80.115 171.295 80.405 172.460 ;
        RECT 81.005 172.435 81.175 173.425 ;
        RECT 81.535 173.230 81.745 173.515 ;
        RECT 82.010 173.505 82.180 173.530 ;
        RECT 82.010 173.335 82.185 173.505 ;
        RECT 82.425 173.465 82.755 173.845 ;
        RECT 82.525 173.385 82.695 173.465 ;
        RECT 82.010 173.235 82.180 173.335 ;
        RECT 81.355 173.060 81.745 173.230 ;
        RECT 81.915 173.065 82.180 173.235 ;
        RECT 82.945 173.215 83.115 173.675 ;
        RECT 83.365 173.385 83.620 173.845 ;
        RECT 81.355 172.605 81.525 173.060 ;
        RECT 81.915 172.855 82.085 173.065 ;
        RECT 82.440 172.935 82.645 173.170 ;
        RECT 82.945 173.045 83.620 173.215 ;
        RECT 81.755 172.685 82.085 172.855 ;
        RECT 81.915 172.670 82.085 172.685 ;
        RECT 82.315 172.605 82.645 172.935 ;
        RECT 82.825 172.685 83.155 172.855 ;
        RECT 82.985 172.435 83.155 172.685 ;
        RECT 80.665 172.265 83.155 172.435 ;
        RECT 80.665 171.465 80.835 172.265 ;
        RECT 83.365 172.095 83.620 173.045 ;
        RECT 81.065 171.925 82.355 172.095 ;
        RECT 81.125 171.505 81.375 171.925 ;
        RECT 81.565 171.295 81.895 171.755 ;
        RECT 82.105 171.505 82.355 171.925 ;
        RECT 82.525 171.295 82.775 172.095 ;
        RECT 82.945 171.925 83.620 172.095 ;
        RECT 83.795 173.170 84.055 173.675 ;
        RECT 84.235 173.465 84.565 173.845 ;
        RECT 84.745 173.295 84.915 173.675 ;
        RECT 83.795 172.370 83.965 173.170 ;
        RECT 84.250 173.125 84.915 173.295 ;
        RECT 84.250 172.870 84.420 173.125 ;
        RECT 85.655 173.115 85.945 173.845 ;
        RECT 84.135 172.540 84.420 172.870 ;
        RECT 84.655 172.575 84.985 172.945 ;
        RECT 85.645 172.605 85.945 172.935 ;
        RECT 86.125 172.915 86.355 173.555 ;
        RECT 86.535 173.295 86.845 173.665 ;
        RECT 87.025 173.475 87.695 173.845 ;
        RECT 86.535 173.095 87.765 173.295 ;
        RECT 86.125 172.605 86.650 172.915 ;
        RECT 86.830 172.605 87.295 172.915 ;
        RECT 84.250 172.395 84.420 172.540 ;
        RECT 87.475 172.425 87.765 173.095 ;
        RECT 82.945 171.465 83.115 171.925 ;
        RECT 83.325 171.295 83.575 171.755 ;
        RECT 83.795 171.465 84.065 172.370 ;
        RECT 84.250 172.225 84.915 172.395 ;
        RECT 84.235 171.295 84.565 172.055 ;
        RECT 84.745 171.465 84.915 172.225 ;
        RECT 85.655 172.185 86.815 172.425 ;
        RECT 85.655 171.475 85.915 172.185 ;
        RECT 86.085 171.295 86.415 172.005 ;
        RECT 86.585 171.475 86.815 172.185 ;
        RECT 86.995 172.205 87.765 172.425 ;
        RECT 86.995 171.475 87.265 172.205 ;
        RECT 87.445 171.295 87.785 172.025 ;
        RECT 87.955 171.475 88.215 173.665 ;
        RECT 88.455 173.365 88.735 173.845 ;
        RECT 88.905 173.195 89.165 173.585 ;
        RECT 89.340 173.365 89.595 173.845 ;
        RECT 89.765 173.195 90.060 173.585 ;
        RECT 90.240 173.365 90.515 173.845 ;
        RECT 90.685 173.345 90.985 173.675 ;
        RECT 88.410 173.025 90.060 173.195 ;
        RECT 88.410 172.515 88.815 173.025 ;
        RECT 88.985 172.685 90.125 172.855 ;
        RECT 88.410 172.345 89.165 172.515 ;
        RECT 88.450 171.295 88.735 172.165 ;
        RECT 88.905 172.095 89.165 172.345 ;
        RECT 89.955 172.435 90.125 172.685 ;
        RECT 90.295 172.605 90.645 173.175 ;
        RECT 90.815 172.435 90.985 173.345 ;
        RECT 91.155 173.045 91.465 173.845 ;
        RECT 91.670 173.045 92.365 173.675 ;
        RECT 92.620 173.345 93.115 173.675 ;
        RECT 91.165 172.605 91.500 172.875 ;
        RECT 91.670 172.445 91.840 173.045 ;
        RECT 92.010 172.605 92.345 172.855 ;
        RECT 89.955 172.265 90.985 172.435 ;
        RECT 88.905 171.925 90.025 172.095 ;
        RECT 88.905 171.465 89.165 171.925 ;
        RECT 89.340 171.295 89.595 171.755 ;
        RECT 89.765 171.465 90.025 171.925 ;
        RECT 90.195 171.295 90.505 172.095 ;
        RECT 90.675 171.465 90.985 172.265 ;
        RECT 91.155 171.295 91.435 172.435 ;
        RECT 91.605 171.465 91.935 172.445 ;
        RECT 92.105 171.295 92.365 172.435 ;
        RECT 92.535 171.855 92.775 173.165 ;
        RECT 92.945 172.435 93.115 173.345 ;
        RECT 93.335 172.605 93.685 173.570 ;
        RECT 93.865 172.605 94.165 173.575 ;
        RECT 94.345 172.605 94.625 173.575 ;
        RECT 94.805 173.045 95.075 173.845 ;
        RECT 95.245 173.125 95.585 173.635 ;
        RECT 97.005 173.445 97.335 173.845 ;
        RECT 97.505 173.275 97.835 173.615 ;
        RECT 98.885 173.445 99.215 173.845 ;
        RECT 94.820 172.605 95.150 172.855 ;
        RECT 94.820 172.435 95.135 172.605 ;
        RECT 92.945 172.265 95.135 172.435 ;
        RECT 92.540 171.295 92.875 171.675 ;
        RECT 93.045 171.465 93.295 172.265 ;
        RECT 93.515 171.295 93.845 172.015 ;
        RECT 94.030 171.465 94.280 172.265 ;
        RECT 94.745 171.295 95.075 172.095 ;
        RECT 95.325 171.725 95.585 173.125 ;
        RECT 96.850 173.105 99.215 173.275 ;
        RECT 99.385 173.120 99.715 173.630 ;
        RECT 96.850 172.105 97.020 173.105 ;
        RECT 99.045 172.935 99.215 173.105 ;
        RECT 97.190 172.275 97.435 172.935 ;
        RECT 97.650 172.275 97.915 172.935 ;
        RECT 98.110 172.275 98.395 172.935 ;
        RECT 98.570 172.605 98.875 172.935 ;
        RECT 99.045 172.605 99.355 172.935 ;
        RECT 98.570 172.275 98.785 172.605 ;
        RECT 96.850 171.935 97.305 172.105 ;
        RECT 95.245 171.465 95.585 171.725 ;
        RECT 96.975 171.505 97.305 171.935 ;
        RECT 97.485 171.935 98.775 172.105 ;
        RECT 97.485 171.515 97.735 171.935 ;
        RECT 97.965 171.295 98.295 171.765 ;
        RECT 98.525 171.515 98.775 171.935 ;
        RECT 98.965 171.295 99.215 172.435 ;
        RECT 99.525 172.355 99.715 173.120 ;
        RECT 99.385 171.505 99.715 172.355 ;
        RECT 99.895 173.105 100.385 173.675 ;
        RECT 100.555 173.275 100.785 173.675 ;
        RECT 100.955 173.445 101.375 173.845 ;
        RECT 101.545 173.275 101.715 173.675 ;
        RECT 100.555 173.105 101.715 173.275 ;
        RECT 101.885 173.105 102.335 173.845 ;
        RECT 102.505 173.105 102.945 173.665 ;
        RECT 99.895 172.435 100.065 173.105 ;
        RECT 100.235 172.605 100.640 172.935 ;
        RECT 99.895 172.265 100.665 172.435 ;
        RECT 99.905 171.295 100.235 172.095 ;
        RECT 100.415 171.635 100.665 172.265 ;
        RECT 100.855 171.805 101.105 172.935 ;
        RECT 101.305 172.605 101.550 172.935 ;
        RECT 101.735 172.655 102.125 172.935 ;
        RECT 101.305 171.805 101.505 172.605 ;
        RECT 102.295 172.485 102.465 172.935 ;
        RECT 101.675 172.315 102.465 172.485 ;
        RECT 101.675 171.635 101.845 172.315 ;
        RECT 100.415 171.465 101.845 171.635 ;
        RECT 102.015 171.295 102.330 172.145 ;
        RECT 102.635 172.095 102.945 173.105 ;
        RECT 103.115 173.095 104.325 173.845 ;
        RECT 103.115 172.555 103.635 173.095 ;
        RECT 104.555 173.025 104.765 173.845 ;
        RECT 104.935 173.045 105.265 173.675 ;
        RECT 103.805 172.385 104.325 172.925 ;
        RECT 104.935 172.445 105.185 173.045 ;
        RECT 105.435 173.025 105.665 173.845 ;
        RECT 105.875 173.120 106.165 173.845 ;
        RECT 106.795 173.345 107.135 173.845 ;
        RECT 105.355 172.605 105.685 172.855 ;
        RECT 106.795 172.605 107.135 173.175 ;
        RECT 107.305 172.935 107.550 173.625 ;
        RECT 107.745 173.345 108.075 173.845 ;
        RECT 108.275 173.275 108.445 173.625 ;
        RECT 108.620 173.445 108.950 173.845 ;
        RECT 109.120 173.275 109.290 173.625 ;
        RECT 109.460 173.445 109.840 173.845 ;
        RECT 108.275 173.105 109.860 173.275 ;
        RECT 110.030 173.170 110.305 173.515 ;
        RECT 109.690 172.935 109.860 173.105 ;
        RECT 107.305 172.605 107.960 172.935 ;
        RECT 102.505 171.465 102.945 172.095 ;
        RECT 103.115 171.295 104.325 172.385 ;
        RECT 104.555 171.295 104.765 172.435 ;
        RECT 104.935 171.465 105.265 172.445 ;
        RECT 105.435 171.295 105.665 172.435 ;
        RECT 105.875 171.295 106.165 172.460 ;
        RECT 106.795 171.295 107.135 172.370 ;
        RECT 107.305 172.010 107.545 172.605 ;
        RECT 107.740 172.145 108.060 172.435 ;
        RECT 108.230 172.315 108.970 172.935 ;
        RECT 109.140 172.605 109.520 172.935 ;
        RECT 109.690 172.605 109.965 172.935 ;
        RECT 109.690 172.435 109.860 172.605 ;
        RECT 110.135 172.435 110.305 173.170 ;
        RECT 109.200 172.265 109.860 172.435 ;
        RECT 109.200 172.145 109.370 172.265 ;
        RECT 107.740 171.975 109.370 172.145 ;
        RECT 107.320 171.515 109.370 171.805 ;
        RECT 109.540 171.295 109.820 172.095 ;
        RECT 110.030 171.465 110.305 172.435 ;
        RECT 110.475 173.170 110.750 173.515 ;
        RECT 110.940 173.445 111.320 173.845 ;
        RECT 111.490 173.275 111.660 173.625 ;
        RECT 111.830 173.445 112.160 173.845 ;
        RECT 112.335 173.275 112.505 173.625 ;
        RECT 112.705 173.345 113.035 173.845 ;
        RECT 110.475 172.435 110.645 173.170 ;
        RECT 110.920 173.105 112.505 173.275 ;
        RECT 110.920 172.935 111.090 173.105 ;
        RECT 113.230 172.935 113.475 173.625 ;
        RECT 113.645 173.345 113.985 173.845 ;
        RECT 110.815 172.605 111.090 172.935 ;
        RECT 111.260 172.605 111.640 172.935 ;
        RECT 110.920 172.435 111.090 172.605 ;
        RECT 110.475 171.465 110.750 172.435 ;
        RECT 110.920 172.265 111.580 172.435 ;
        RECT 111.810 172.315 112.550 172.935 ;
        RECT 112.820 172.605 113.475 172.935 ;
        RECT 113.645 172.605 113.985 173.175 ;
        RECT 114.155 173.105 114.540 173.675 ;
        RECT 114.710 173.385 115.035 173.845 ;
        RECT 115.555 173.215 115.835 173.675 ;
        RECT 111.410 172.145 111.580 172.265 ;
        RECT 112.720 172.145 113.040 172.435 ;
        RECT 110.960 171.295 111.240 172.095 ;
        RECT 111.410 171.975 113.040 172.145 ;
        RECT 113.235 172.010 113.475 172.605 ;
        RECT 114.155 172.435 114.435 173.105 ;
        RECT 114.710 173.045 115.835 173.215 ;
        RECT 114.710 172.935 115.160 173.045 ;
        RECT 114.605 172.605 115.160 172.935 ;
        RECT 116.025 172.875 116.425 173.675 ;
        RECT 116.825 173.385 117.095 173.845 ;
        RECT 117.265 173.215 117.550 173.675 ;
        RECT 117.845 173.345 118.175 173.845 ;
        RECT 111.410 171.515 113.460 171.805 ;
        RECT 113.645 171.295 113.985 172.370 ;
        RECT 114.155 171.465 114.540 172.435 ;
        RECT 114.710 172.145 115.160 172.605 ;
        RECT 115.330 172.315 116.425 172.875 ;
        RECT 114.710 171.925 115.835 172.145 ;
        RECT 114.710 171.295 115.035 171.755 ;
        RECT 115.555 171.465 115.835 171.925 ;
        RECT 116.025 171.465 116.425 172.315 ;
        RECT 116.595 173.045 117.550 173.215 ;
        RECT 118.375 173.275 118.545 173.625 ;
        RECT 118.745 173.445 119.075 173.845 ;
        RECT 119.245 173.275 119.415 173.625 ;
        RECT 119.585 173.445 119.965 173.845 ;
        RECT 116.595 172.145 116.805 173.045 ;
        RECT 116.975 172.315 117.665 172.875 ;
        RECT 117.840 172.605 118.190 173.175 ;
        RECT 118.375 173.105 119.985 173.275 ;
        RECT 120.155 173.170 120.425 173.515 ;
        RECT 119.815 172.935 119.985 173.105 ;
        RECT 117.840 172.145 118.160 172.435 ;
        RECT 118.360 172.315 119.070 172.935 ;
        RECT 119.240 172.605 119.645 172.935 ;
        RECT 119.815 172.605 120.085 172.935 ;
        RECT 119.815 172.435 119.985 172.605 ;
        RECT 120.255 172.435 120.425 173.170 ;
        RECT 120.595 173.120 120.935 173.845 ;
        RECT 121.105 172.935 121.310 173.535 ;
        RECT 121.540 173.330 122.490 173.515 ;
        RECT 119.260 172.265 119.985 172.435 ;
        RECT 119.260 172.145 119.430 172.265 ;
        RECT 116.595 171.925 117.550 172.145 ;
        RECT 117.840 171.975 119.430 172.145 ;
        RECT 116.825 171.295 117.095 171.755 ;
        RECT 117.265 171.465 117.550 171.925 ;
        RECT 117.840 171.515 119.495 171.805 ;
        RECT 119.665 171.295 119.945 172.095 ;
        RECT 120.155 171.465 120.425 172.435 ;
        RECT 120.620 172.305 120.875 172.935 ;
        RECT 121.105 172.305 121.485 172.935 ;
        RECT 121.745 172.605 121.965 173.330 ;
        RECT 122.660 173.195 123.075 173.630 ;
        RECT 123.265 173.365 123.595 173.845 ;
        RECT 123.765 173.370 124.105 173.630 ;
        RECT 122.660 173.120 123.675 173.195 ;
        RECT 122.855 173.025 123.675 173.120 ;
        RECT 122.275 172.825 122.655 172.935 ;
        RECT 122.275 172.655 122.665 172.825 ;
        RECT 122.275 172.605 122.655 172.655 ;
        RECT 122.355 172.310 122.655 172.605 ;
        RECT 122.855 172.295 123.185 172.855 ;
        RECT 120.685 171.965 122.655 172.135 ;
        RECT 123.505 172.105 123.675 173.025 ;
        RECT 120.685 171.465 120.855 171.965 ;
        RECT 121.095 171.295 121.345 171.755 ;
        RECT 121.645 171.465 121.815 171.965 ;
        RECT 122.025 171.295 122.275 171.755 ;
        RECT 122.485 171.465 122.655 171.965 ;
        RECT 122.825 171.935 123.675 172.105 ;
        RECT 122.825 171.505 123.155 171.935 ;
        RECT 123.845 171.765 124.105 173.370 ;
        RECT 124.275 173.185 124.550 173.845 ;
        RECT 124.720 173.215 124.970 173.675 ;
        RECT 125.145 173.350 125.475 173.845 ;
        RECT 124.720 173.005 124.890 173.215 ;
        RECT 125.655 173.180 125.885 173.625 ;
        RECT 124.275 172.485 124.890 173.005 ;
        RECT 125.060 172.505 125.290 172.935 ;
        RECT 125.475 172.685 125.885 173.180 ;
        RECT 126.055 173.360 126.845 173.625 ;
        RECT 126.055 172.505 126.310 173.360 ;
        RECT 127.035 173.195 127.295 173.675 ;
        RECT 127.465 173.305 127.715 173.845 ;
        RECT 126.480 172.685 126.865 173.165 ;
        RECT 123.345 171.295 123.595 171.755 ;
        RECT 123.765 171.505 124.105 171.765 ;
        RECT 124.275 171.295 124.535 172.305 ;
        RECT 124.705 172.135 124.875 172.485 ;
        RECT 125.060 172.335 126.850 172.505 ;
        RECT 124.705 171.465 124.980 172.135 ;
        RECT 125.180 171.295 125.395 172.140 ;
        RECT 125.620 172.040 125.870 172.335 ;
        RECT 126.095 171.975 126.425 172.165 ;
        RECT 125.580 171.465 126.055 171.805 ;
        RECT 126.235 171.800 126.425 171.975 ;
        RECT 126.595 171.970 126.850 172.335 ;
        RECT 127.035 172.165 127.205 173.195 ;
        RECT 127.885 173.140 128.105 173.625 ;
        RECT 127.375 172.545 127.605 172.940 ;
        RECT 127.775 172.715 128.105 173.140 ;
        RECT 128.275 173.465 129.165 173.635 ;
        RECT 128.275 172.740 128.445 173.465 ;
        RECT 128.615 172.910 129.165 173.295 ;
        RECT 129.335 173.075 131.005 173.845 ;
        RECT 131.635 173.120 131.925 173.845 ;
        RECT 132.095 173.075 134.685 173.845 ;
        RECT 134.855 173.105 135.240 173.675 ;
        RECT 135.410 173.385 135.735 173.845 ;
        RECT 136.255 173.215 136.535 173.675 ;
        RECT 128.275 172.670 129.165 172.740 ;
        RECT 128.270 172.645 129.165 172.670 ;
        RECT 128.260 172.630 129.165 172.645 ;
        RECT 128.255 172.615 129.165 172.630 ;
        RECT 128.245 172.610 129.165 172.615 ;
        RECT 128.240 172.600 129.165 172.610 ;
        RECT 128.235 172.590 129.165 172.600 ;
        RECT 128.225 172.585 129.165 172.590 ;
        RECT 128.215 172.575 129.165 172.585 ;
        RECT 128.205 172.570 129.165 172.575 ;
        RECT 128.205 172.565 128.540 172.570 ;
        RECT 128.190 172.560 128.540 172.565 ;
        RECT 128.175 172.550 128.540 172.560 ;
        RECT 128.150 172.545 128.540 172.550 ;
        RECT 127.375 172.540 128.540 172.545 ;
        RECT 127.375 172.505 128.510 172.540 ;
        RECT 127.375 172.480 128.475 172.505 ;
        RECT 127.375 172.450 128.445 172.480 ;
        RECT 127.375 172.420 128.425 172.450 ;
        RECT 127.375 172.390 128.405 172.420 ;
        RECT 127.375 172.380 128.335 172.390 ;
        RECT 127.375 172.370 128.310 172.380 ;
        RECT 127.375 172.355 128.290 172.370 ;
        RECT 127.375 172.340 128.270 172.355 ;
        RECT 127.480 172.330 128.265 172.340 ;
        RECT 127.480 172.295 128.250 172.330 ;
        RECT 126.235 171.295 126.865 171.800 ;
        RECT 127.035 171.465 127.310 172.165 ;
        RECT 127.480 172.045 128.235 172.295 ;
        RECT 128.405 171.975 128.735 172.220 ;
        RECT 128.905 172.120 129.165 172.570 ;
        RECT 129.335 172.555 130.085 173.075 ;
        RECT 130.255 172.385 131.005 172.905 ;
        RECT 132.095 172.555 133.305 173.075 ;
        RECT 128.550 171.950 128.735 171.975 ;
        RECT 128.550 171.850 129.165 171.950 ;
        RECT 127.480 171.295 127.735 171.840 ;
        RECT 127.905 171.465 128.385 171.805 ;
        RECT 128.560 171.295 129.165 171.850 ;
        RECT 129.335 171.295 131.005 172.385 ;
        RECT 131.635 171.295 131.925 172.460 ;
        RECT 133.475 172.385 134.685 172.905 ;
        RECT 132.095 171.295 134.685 172.385 ;
        RECT 134.855 172.435 135.135 173.105 ;
        RECT 135.410 173.045 136.535 173.215 ;
        RECT 135.410 172.935 135.860 173.045 ;
        RECT 135.305 172.605 135.860 172.935 ;
        RECT 136.725 172.875 137.125 173.675 ;
        RECT 137.525 173.385 137.795 173.845 ;
        RECT 137.965 173.215 138.250 173.675 ;
        RECT 138.535 173.300 143.880 173.845 ;
        RECT 144.055 173.300 149.400 173.845 ;
        RECT 149.575 173.300 154.920 173.845 ;
        RECT 134.855 171.465 135.240 172.435 ;
        RECT 135.410 172.145 135.860 172.605 ;
        RECT 136.030 172.315 137.125 172.875 ;
        RECT 135.410 171.925 136.535 172.145 ;
        RECT 135.410 171.295 135.735 171.755 ;
        RECT 136.255 171.465 136.535 171.925 ;
        RECT 136.725 171.465 137.125 172.315 ;
        RECT 137.295 173.045 138.250 173.215 ;
        RECT 137.295 172.145 137.505 173.045 ;
        RECT 137.675 172.315 138.365 172.875 ;
        RECT 140.120 172.470 140.460 173.300 ;
        RECT 137.295 171.925 138.250 172.145 ;
        RECT 137.525 171.295 137.795 171.755 ;
        RECT 137.965 171.465 138.250 171.925 ;
        RECT 141.940 171.730 142.290 172.980 ;
        RECT 145.640 172.470 145.980 173.300 ;
        RECT 147.460 171.730 147.810 172.980 ;
        RECT 151.160 172.470 151.500 173.300 ;
        RECT 155.095 173.075 156.765 173.845 ;
        RECT 156.935 173.095 158.145 173.845 ;
        RECT 152.980 171.730 153.330 172.980 ;
        RECT 155.095 172.555 155.845 173.075 ;
        RECT 156.015 172.385 156.765 172.905 ;
        RECT 138.535 171.295 143.880 171.730 ;
        RECT 144.055 171.295 149.400 171.730 ;
        RECT 149.575 171.295 154.920 171.730 ;
        RECT 155.095 171.295 156.765 172.385 ;
        RECT 156.935 172.385 157.455 172.925 ;
        RECT 157.625 172.555 158.145 173.095 ;
        RECT 156.935 171.295 158.145 172.385 ;
        RECT 2.750 171.125 158.230 171.295 ;
        RECT 2.835 170.035 4.045 171.125 ;
        RECT 4.220 170.455 4.475 170.955 ;
        RECT 4.645 170.625 4.975 171.125 ;
        RECT 4.220 170.285 4.970 170.455 ;
        RECT 2.835 169.325 3.355 169.865 ;
        RECT 3.525 169.495 4.045 170.035 ;
        RECT 4.220 169.465 4.570 170.115 ;
        RECT 2.835 168.575 4.045 169.325 ;
        RECT 4.740 169.295 4.970 170.285 ;
        RECT 4.220 169.125 4.970 169.295 ;
        RECT 4.220 168.835 4.475 169.125 ;
        RECT 4.645 168.575 4.975 168.955 ;
        RECT 5.145 168.835 5.315 170.955 ;
        RECT 5.485 170.155 5.810 170.940 ;
        RECT 5.980 170.665 6.230 171.125 ;
        RECT 6.400 170.625 6.650 170.955 ;
        RECT 6.865 170.625 7.545 170.955 ;
        RECT 6.400 170.495 6.570 170.625 ;
        RECT 6.175 170.325 6.570 170.495 ;
        RECT 5.545 169.105 6.005 170.155 ;
        RECT 6.175 168.965 6.345 170.325 ;
        RECT 6.740 170.065 7.205 170.455 ;
        RECT 6.515 169.255 6.865 169.875 ;
        RECT 7.035 169.475 7.205 170.065 ;
        RECT 7.375 169.845 7.545 170.625 ;
        RECT 7.715 170.525 7.885 170.865 ;
        RECT 8.120 170.695 8.450 171.125 ;
        RECT 8.620 170.525 8.790 170.865 ;
        RECT 9.085 170.665 9.455 171.125 ;
        RECT 7.715 170.355 8.790 170.525 ;
        RECT 9.625 170.495 9.795 170.955 ;
        RECT 10.030 170.615 10.900 170.955 ;
        RECT 11.070 170.665 11.320 171.125 ;
        RECT 9.235 170.325 9.795 170.495 ;
        RECT 9.235 170.185 9.405 170.325 ;
        RECT 7.905 170.015 9.405 170.185 ;
        RECT 10.100 170.155 10.560 170.445 ;
        RECT 7.375 169.675 9.065 169.845 ;
        RECT 7.035 169.255 7.390 169.475 ;
        RECT 7.560 168.965 7.730 169.675 ;
        RECT 7.935 169.255 8.725 169.505 ;
        RECT 8.895 169.495 9.065 169.675 ;
        RECT 9.235 169.325 9.405 170.015 ;
        RECT 5.675 168.575 6.005 168.935 ;
        RECT 6.175 168.795 6.670 168.965 ;
        RECT 6.875 168.795 7.730 168.965 ;
        RECT 8.605 168.575 8.935 169.035 ;
        RECT 9.145 168.935 9.405 169.325 ;
        RECT 9.595 170.145 10.560 170.155 ;
        RECT 10.730 170.235 10.900 170.615 ;
        RECT 11.490 170.575 11.660 170.865 ;
        RECT 11.840 170.745 12.170 171.125 ;
        RECT 11.490 170.405 12.290 170.575 ;
        RECT 9.595 169.985 10.270 170.145 ;
        RECT 10.730 170.065 11.950 170.235 ;
        RECT 9.595 169.195 9.805 169.985 ;
        RECT 10.730 169.975 10.900 170.065 ;
        RECT 9.975 169.195 10.325 169.815 ;
        RECT 10.495 169.805 10.900 169.975 ;
        RECT 10.495 169.025 10.665 169.805 ;
        RECT 10.835 169.355 11.055 169.635 ;
        RECT 11.235 169.525 11.775 169.895 ;
        RECT 12.120 169.815 12.290 170.405 ;
        RECT 12.510 169.985 12.815 171.125 ;
        RECT 12.985 169.935 13.240 170.815 ;
        RECT 14.425 170.195 14.595 170.955 ;
        RECT 14.775 170.365 15.105 171.125 ;
        RECT 14.425 170.025 15.090 170.195 ;
        RECT 15.275 170.050 15.545 170.955 ;
        RECT 12.120 169.785 12.860 169.815 ;
        RECT 10.835 169.185 11.365 169.355 ;
        RECT 9.145 168.765 9.495 168.935 ;
        RECT 9.715 168.745 10.665 169.025 ;
        RECT 10.835 168.575 11.025 169.015 ;
        RECT 11.195 168.955 11.365 169.185 ;
        RECT 11.535 169.125 11.775 169.525 ;
        RECT 11.945 169.485 12.860 169.785 ;
        RECT 11.945 169.310 12.270 169.485 ;
        RECT 11.945 168.955 12.265 169.310 ;
        RECT 13.030 169.285 13.240 169.935 ;
        RECT 14.920 169.880 15.090 170.025 ;
        RECT 14.355 169.475 14.685 169.845 ;
        RECT 14.920 169.550 15.205 169.880 ;
        RECT 14.920 169.295 15.090 169.550 ;
        RECT 11.195 168.785 12.265 168.955 ;
        RECT 12.510 168.575 12.815 169.035 ;
        RECT 12.985 168.755 13.240 169.285 ;
        RECT 14.425 169.125 15.090 169.295 ;
        RECT 15.375 169.250 15.545 170.050 ;
        RECT 15.715 169.960 16.005 171.125 ;
        RECT 16.265 170.455 16.435 170.955 ;
        RECT 16.605 170.625 16.935 171.125 ;
        RECT 16.265 170.285 16.930 170.455 ;
        RECT 16.180 169.465 16.530 170.115 ;
        RECT 14.425 168.745 14.595 169.125 ;
        RECT 14.775 168.575 15.105 168.955 ;
        RECT 15.285 168.745 15.545 169.250 ;
        RECT 15.715 168.575 16.005 169.300 ;
        RECT 16.700 169.295 16.930 170.285 ;
        RECT 16.265 169.125 16.930 169.295 ;
        RECT 16.265 168.835 16.435 169.125 ;
        RECT 16.605 168.575 16.935 168.955 ;
        RECT 17.105 168.835 17.330 170.955 ;
        RECT 17.545 170.625 17.875 171.125 ;
        RECT 18.045 170.455 18.215 170.955 ;
        RECT 18.450 170.740 19.280 170.910 ;
        RECT 19.520 170.745 19.900 171.125 ;
        RECT 17.520 170.285 18.215 170.455 ;
        RECT 17.520 169.315 17.690 170.285 ;
        RECT 17.860 169.495 18.270 170.115 ;
        RECT 18.440 170.065 18.940 170.445 ;
        RECT 17.520 169.125 18.215 169.315 ;
        RECT 18.440 169.195 18.660 170.065 ;
        RECT 19.110 169.895 19.280 170.740 ;
        RECT 20.080 170.575 20.250 170.865 ;
        RECT 20.420 170.745 20.750 171.125 ;
        RECT 21.220 170.655 21.850 170.905 ;
        RECT 22.030 170.745 22.450 171.125 ;
        RECT 21.680 170.575 21.850 170.655 ;
        RECT 22.650 170.575 22.890 170.865 ;
        RECT 19.450 170.325 20.820 170.575 ;
        RECT 19.450 170.065 19.700 170.325 ;
        RECT 20.210 169.895 20.460 170.055 ;
        RECT 19.110 169.725 20.460 169.895 ;
        RECT 19.110 169.685 19.530 169.725 ;
        RECT 18.840 169.135 19.190 169.505 ;
        RECT 17.545 168.575 17.875 168.955 ;
        RECT 18.045 168.795 18.215 169.125 ;
        RECT 19.360 168.955 19.530 169.685 ;
        RECT 20.630 169.555 20.820 170.325 ;
        RECT 19.700 169.225 20.110 169.555 ;
        RECT 20.400 169.215 20.820 169.555 ;
        RECT 20.990 170.145 21.510 170.455 ;
        RECT 21.680 170.405 22.890 170.575 ;
        RECT 23.120 170.435 23.450 171.125 ;
        RECT 20.990 169.385 21.160 170.145 ;
        RECT 21.330 169.555 21.510 169.965 ;
        RECT 21.680 169.895 21.850 170.405 ;
        RECT 23.620 170.255 23.790 170.865 ;
        RECT 24.060 170.405 24.390 170.915 ;
        RECT 23.620 170.235 23.940 170.255 ;
        RECT 22.020 170.065 23.940 170.235 ;
        RECT 21.680 169.725 23.580 169.895 ;
        RECT 21.910 169.385 22.240 169.505 ;
        RECT 20.990 169.215 22.240 169.385 ;
        RECT 18.515 168.755 19.530 168.955 ;
        RECT 19.700 168.575 20.110 169.015 ;
        RECT 20.400 168.785 20.650 169.215 ;
        RECT 20.850 168.575 21.170 169.035 ;
        RECT 22.410 168.965 22.580 169.725 ;
        RECT 23.250 169.665 23.580 169.725 ;
        RECT 22.770 169.495 23.100 169.555 ;
        RECT 22.770 169.225 23.430 169.495 ;
        RECT 23.750 169.170 23.940 170.065 ;
        RECT 21.730 168.795 22.580 168.965 ;
        RECT 22.780 168.575 23.440 169.055 ;
        RECT 23.620 168.840 23.940 169.170 ;
        RECT 24.140 169.815 24.390 170.405 ;
        RECT 24.570 170.325 24.855 171.125 ;
        RECT 25.035 170.785 25.290 170.815 ;
        RECT 25.035 170.615 25.375 170.785 ;
        RECT 25.035 170.145 25.290 170.615 ;
        RECT 24.140 169.485 24.940 169.815 ;
        RECT 24.140 168.835 24.390 169.485 ;
        RECT 25.110 169.285 25.290 170.145 ;
        RECT 25.835 170.035 28.425 171.125 ;
        RECT 28.600 170.455 28.855 170.955 ;
        RECT 29.025 170.625 29.355 171.125 ;
        RECT 28.600 170.285 29.350 170.455 ;
        RECT 24.570 168.575 24.855 169.035 ;
        RECT 25.035 168.755 25.290 169.285 ;
        RECT 25.835 169.345 27.045 169.865 ;
        RECT 27.215 169.515 28.425 170.035 ;
        RECT 28.600 169.465 28.950 170.115 ;
        RECT 25.835 168.575 28.425 169.345 ;
        RECT 29.120 169.295 29.350 170.285 ;
        RECT 28.600 169.125 29.350 169.295 ;
        RECT 28.600 168.835 28.855 169.125 ;
        RECT 29.025 168.575 29.355 168.955 ;
        RECT 29.525 168.835 29.695 170.955 ;
        RECT 29.865 170.155 30.190 170.940 ;
        RECT 30.360 170.665 30.610 171.125 ;
        RECT 30.780 170.625 31.030 170.955 ;
        RECT 31.245 170.625 31.925 170.955 ;
        RECT 30.780 170.495 30.950 170.625 ;
        RECT 30.555 170.325 30.950 170.495 ;
        RECT 29.925 169.105 30.385 170.155 ;
        RECT 30.555 168.965 30.725 170.325 ;
        RECT 31.120 170.065 31.585 170.455 ;
        RECT 30.895 169.255 31.245 169.875 ;
        RECT 31.415 169.475 31.585 170.065 ;
        RECT 31.755 169.845 31.925 170.625 ;
        RECT 32.095 170.525 32.265 170.865 ;
        RECT 32.500 170.695 32.830 171.125 ;
        RECT 33.000 170.525 33.170 170.865 ;
        RECT 33.465 170.665 33.835 171.125 ;
        RECT 32.095 170.355 33.170 170.525 ;
        RECT 34.005 170.495 34.175 170.955 ;
        RECT 34.410 170.615 35.280 170.955 ;
        RECT 35.450 170.665 35.700 171.125 ;
        RECT 33.615 170.325 34.175 170.495 ;
        RECT 33.615 170.185 33.785 170.325 ;
        RECT 32.285 170.015 33.785 170.185 ;
        RECT 34.480 170.155 34.940 170.445 ;
        RECT 31.755 169.675 33.445 169.845 ;
        RECT 31.415 169.255 31.770 169.475 ;
        RECT 31.940 168.965 32.110 169.675 ;
        RECT 32.315 169.255 33.105 169.505 ;
        RECT 33.275 169.495 33.445 169.675 ;
        RECT 33.615 169.325 33.785 170.015 ;
        RECT 30.055 168.575 30.385 168.935 ;
        RECT 30.555 168.795 31.050 168.965 ;
        RECT 31.255 168.795 32.110 168.965 ;
        RECT 32.985 168.575 33.315 169.035 ;
        RECT 33.525 168.935 33.785 169.325 ;
        RECT 33.975 170.145 34.940 170.155 ;
        RECT 35.110 170.235 35.280 170.615 ;
        RECT 35.870 170.575 36.040 170.865 ;
        RECT 36.220 170.745 36.550 171.125 ;
        RECT 35.870 170.405 36.670 170.575 ;
        RECT 33.975 169.985 34.650 170.145 ;
        RECT 35.110 170.065 36.330 170.235 ;
        RECT 33.975 169.195 34.185 169.985 ;
        RECT 35.110 169.975 35.280 170.065 ;
        RECT 34.355 169.195 34.705 169.815 ;
        RECT 34.875 169.805 35.280 169.975 ;
        RECT 34.875 169.025 35.045 169.805 ;
        RECT 35.215 169.355 35.435 169.635 ;
        RECT 35.615 169.525 36.155 169.895 ;
        RECT 36.500 169.815 36.670 170.405 ;
        RECT 36.890 169.985 37.195 171.125 ;
        RECT 37.365 169.935 37.620 170.815 ;
        RECT 36.500 169.785 37.240 169.815 ;
        RECT 35.215 169.185 35.745 169.355 ;
        RECT 33.525 168.765 33.875 168.935 ;
        RECT 34.095 168.745 35.045 169.025 ;
        RECT 35.215 168.575 35.405 169.015 ;
        RECT 35.575 168.955 35.745 169.185 ;
        RECT 35.915 169.125 36.155 169.525 ;
        RECT 36.325 169.485 37.240 169.785 ;
        RECT 36.325 169.310 36.650 169.485 ;
        RECT 36.325 168.955 36.645 169.310 ;
        RECT 37.410 169.285 37.620 169.935 ;
        RECT 35.575 168.785 36.645 168.955 ;
        RECT 36.890 168.575 37.195 169.035 ;
        RECT 37.365 168.755 37.620 169.285 ;
        RECT 38.715 170.050 38.985 170.955 ;
        RECT 39.155 170.365 39.485 171.125 ;
        RECT 39.665 170.195 39.835 170.955 ;
        RECT 38.715 169.250 38.885 170.050 ;
        RECT 39.170 170.025 39.835 170.195 ;
        RECT 40.185 170.195 40.355 170.955 ;
        RECT 40.535 170.365 40.865 171.125 ;
        RECT 40.185 170.025 40.850 170.195 ;
        RECT 41.035 170.050 41.305 170.955 ;
        RECT 39.170 169.880 39.340 170.025 ;
        RECT 39.055 169.550 39.340 169.880 ;
        RECT 40.680 169.880 40.850 170.025 ;
        RECT 39.170 169.295 39.340 169.550 ;
        RECT 39.575 169.475 39.905 169.845 ;
        RECT 40.115 169.475 40.445 169.845 ;
        RECT 40.680 169.550 40.965 169.880 ;
        RECT 40.680 169.295 40.850 169.550 ;
        RECT 38.715 168.745 38.975 169.250 ;
        RECT 39.170 169.125 39.835 169.295 ;
        RECT 39.155 168.575 39.485 168.955 ;
        RECT 39.665 168.745 39.835 169.125 ;
        RECT 40.185 169.125 40.850 169.295 ;
        RECT 41.135 169.250 41.305 170.050 ;
        RECT 41.475 169.960 41.765 171.125 ;
        RECT 41.935 170.365 42.450 170.775 ;
        RECT 42.685 170.365 42.855 171.125 ;
        RECT 43.025 170.785 45.055 170.955 ;
        RECT 41.935 169.555 42.275 170.365 ;
        RECT 43.025 170.120 43.195 170.785 ;
        RECT 43.590 170.445 44.715 170.615 ;
        RECT 42.445 169.930 43.195 170.120 ;
        RECT 43.365 170.105 44.375 170.275 ;
        RECT 41.935 169.385 43.165 169.555 ;
        RECT 40.185 168.745 40.355 169.125 ;
        RECT 40.535 168.575 40.865 168.955 ;
        RECT 41.045 168.745 41.305 169.250 ;
        RECT 41.475 168.575 41.765 169.300 ;
        RECT 42.210 168.780 42.455 169.385 ;
        RECT 42.675 168.575 43.185 169.110 ;
        RECT 43.365 168.745 43.555 170.105 ;
        RECT 43.725 169.425 44.000 169.905 ;
        RECT 43.725 169.255 44.005 169.425 ;
        RECT 44.205 169.305 44.375 170.105 ;
        RECT 44.545 169.315 44.715 170.445 ;
        RECT 44.885 169.815 45.055 170.785 ;
        RECT 45.225 169.985 45.395 171.125 ;
        RECT 45.565 169.985 45.900 170.955 ;
        RECT 46.085 170.515 46.415 170.945 ;
        RECT 46.595 170.685 46.790 171.125 ;
        RECT 46.960 170.515 47.290 170.945 ;
        RECT 46.085 170.345 47.290 170.515 ;
        RECT 46.085 170.015 46.980 170.345 ;
        RECT 47.460 170.175 47.735 170.945 ;
        RECT 44.885 169.485 45.080 169.815 ;
        RECT 45.305 169.485 45.560 169.815 ;
        RECT 45.305 169.315 45.475 169.485 ;
        RECT 45.730 169.315 45.900 169.985 ;
        RECT 47.150 169.985 47.735 170.175 ;
        RECT 47.955 170.175 48.245 170.945 ;
        RECT 48.815 170.585 49.075 170.945 ;
        RECT 49.245 170.755 49.575 171.125 ;
        RECT 49.745 170.585 50.005 170.945 ;
        RECT 48.815 170.355 50.005 170.585 ;
        RECT 50.195 170.405 50.525 171.125 ;
        RECT 50.695 170.175 50.960 170.945 ;
        RECT 47.955 169.995 50.450 170.175 ;
        RECT 46.090 169.485 46.385 169.815 ;
        RECT 46.565 169.485 46.980 169.815 ;
        RECT 43.725 168.745 44.000 169.255 ;
        RECT 44.545 169.145 45.475 169.315 ;
        RECT 44.545 169.110 44.720 169.145 ;
        RECT 44.190 168.745 44.720 169.110 ;
        RECT 45.145 168.575 45.475 168.975 ;
        RECT 45.645 168.745 45.900 169.315 ;
        RECT 46.085 168.575 46.385 169.305 ;
        RECT 46.565 168.865 46.795 169.485 ;
        RECT 47.150 169.315 47.325 169.985 ;
        RECT 46.995 169.135 47.325 169.315 ;
        RECT 47.495 169.165 47.735 169.815 ;
        RECT 47.925 169.485 48.195 169.815 ;
        RECT 48.375 169.485 48.810 169.815 ;
        RECT 48.990 169.485 49.565 169.815 ;
        RECT 49.745 169.485 50.025 169.815 ;
        RECT 50.225 169.305 50.450 169.995 ;
        RECT 46.995 168.755 47.220 169.135 ;
        RECT 47.965 169.115 50.450 169.305 ;
        RECT 47.390 168.575 47.720 168.965 ;
        RECT 47.965 168.755 48.190 169.115 ;
        RECT 48.370 168.575 48.700 168.945 ;
        RECT 48.880 168.755 49.135 169.115 ;
        RECT 49.700 168.575 50.445 168.945 ;
        RECT 50.625 168.755 50.960 170.175 ;
        RECT 51.145 170.155 51.475 170.940 ;
        RECT 51.145 169.985 51.825 170.155 ;
        RECT 52.005 169.985 52.335 171.125 ;
        RECT 52.525 170.175 52.800 170.945 ;
        RECT 52.970 170.515 53.300 170.945 ;
        RECT 53.470 170.685 53.665 171.125 ;
        RECT 53.845 170.515 54.175 170.945 ;
        RECT 54.355 170.615 56.015 170.905 ;
        RECT 52.970 170.345 54.175 170.515 ;
        RECT 52.525 169.985 53.110 170.175 ;
        RECT 53.280 170.015 54.175 170.345 ;
        RECT 54.355 170.275 55.950 170.445 ;
        RECT 56.185 170.325 56.465 171.125 ;
        RECT 54.355 169.985 54.680 170.275 ;
        RECT 55.780 170.155 55.950 170.275 ;
        RECT 51.135 169.565 51.485 169.815 ;
        RECT 51.655 169.385 51.825 169.985 ;
        RECT 51.995 169.565 52.345 169.815 ;
        RECT 51.155 168.575 51.395 169.385 ;
        RECT 51.565 168.745 51.895 169.385 ;
        RECT 52.065 168.575 52.335 169.385 ;
        RECT 52.525 169.165 52.765 169.815 ;
        RECT 52.935 169.315 53.110 169.985 ;
        RECT 53.280 169.485 53.695 169.815 ;
        RECT 53.875 169.485 54.170 169.815 ;
        RECT 52.935 169.135 53.265 169.315 ;
        RECT 52.540 168.575 52.870 168.965 ;
        RECT 53.040 168.755 53.265 169.135 ;
        RECT 53.465 168.865 53.695 169.485 ;
        RECT 53.875 168.575 54.175 169.305 ;
        RECT 54.355 169.245 54.710 169.815 ;
        RECT 54.880 169.485 55.590 170.105 ;
        RECT 55.780 169.985 56.505 170.155 ;
        RECT 56.675 169.985 56.950 170.955 ;
        RECT 56.335 169.815 56.505 169.985 ;
        RECT 55.760 169.485 56.165 169.815 ;
        RECT 56.335 169.485 56.610 169.815 ;
        RECT 56.335 169.315 56.505 169.485 ;
        RECT 54.895 169.145 56.505 169.315 ;
        RECT 56.780 169.250 56.950 169.985 ;
        RECT 57.120 169.945 57.290 171.125 ;
        RECT 57.730 170.115 58.030 170.955 ;
        RECT 58.225 170.285 58.475 171.125 ;
        RECT 59.065 170.535 59.870 170.955 ;
        RECT 58.645 170.365 60.210 170.535 ;
        RECT 58.645 170.115 58.815 170.365 ;
        RECT 57.730 169.945 58.815 170.115 ;
        RECT 54.360 168.575 54.695 169.075 ;
        RECT 54.895 168.795 55.065 169.145 ;
        RECT 55.265 168.575 55.595 168.975 ;
        RECT 55.765 168.795 55.935 169.145 ;
        RECT 56.105 168.575 56.485 168.975 ;
        RECT 56.675 168.905 56.950 169.250 ;
        RECT 57.120 168.575 57.290 169.490 ;
        RECT 57.575 169.485 57.905 169.775 ;
        RECT 58.075 169.315 58.245 169.945 ;
        RECT 58.985 169.815 59.305 170.195 ;
        RECT 58.415 169.565 58.745 169.775 ;
        RECT 58.925 169.565 59.305 169.815 ;
        RECT 59.495 169.775 59.870 170.195 ;
        RECT 60.040 170.115 60.210 170.365 ;
        RECT 60.380 170.285 60.710 171.125 ;
        RECT 60.880 170.365 61.545 170.955 ;
        RECT 60.040 169.945 60.960 170.115 ;
        RECT 60.790 169.775 60.960 169.945 ;
        RECT 59.495 169.765 59.980 169.775 ;
        RECT 59.475 169.595 59.980 169.765 ;
        RECT 59.495 169.565 59.980 169.595 ;
        RECT 60.170 169.565 60.620 169.775 ;
        RECT 60.790 169.565 61.125 169.775 ;
        RECT 61.295 169.395 61.545 170.365 ;
        RECT 61.715 170.035 62.925 171.125 ;
        RECT 57.735 169.135 58.245 169.315 ;
        RECT 58.650 169.225 60.350 169.395 ;
        RECT 58.650 169.135 59.035 169.225 ;
        RECT 57.735 168.745 58.065 169.135 ;
        RECT 58.235 168.795 59.420 168.965 ;
        RECT 59.680 168.575 59.850 169.045 ;
        RECT 60.020 168.760 60.350 169.225 ;
        RECT 60.520 168.575 60.690 169.395 ;
        RECT 60.860 168.755 61.545 169.395 ;
        RECT 61.715 169.325 62.235 169.865 ;
        RECT 62.405 169.495 62.925 170.035 ;
        RECT 63.250 170.115 63.550 170.955 ;
        RECT 63.745 170.285 63.995 171.125 ;
        RECT 64.585 170.535 65.390 170.955 ;
        RECT 64.165 170.365 65.730 170.535 ;
        RECT 64.165 170.115 64.335 170.365 ;
        RECT 63.250 169.945 64.335 170.115 ;
        RECT 63.095 169.485 63.425 169.775 ;
        RECT 61.715 168.575 62.925 169.325 ;
        RECT 63.595 169.315 63.765 169.945 ;
        RECT 64.505 169.815 64.825 170.195 ;
        RECT 63.935 169.565 64.265 169.775 ;
        RECT 64.445 169.565 64.825 169.815 ;
        RECT 65.015 169.775 65.390 170.195 ;
        RECT 65.560 170.115 65.730 170.365 ;
        RECT 65.900 170.285 66.230 171.125 ;
        RECT 66.400 170.365 67.065 170.955 ;
        RECT 65.560 169.945 66.480 170.115 ;
        RECT 66.310 169.775 66.480 169.945 ;
        RECT 65.015 169.765 65.500 169.775 ;
        RECT 64.995 169.595 65.500 169.765 ;
        RECT 65.015 169.565 65.500 169.595 ;
        RECT 65.690 169.565 66.140 169.775 ;
        RECT 66.310 169.565 66.645 169.775 ;
        RECT 66.815 169.395 67.065 170.365 ;
        RECT 67.235 169.960 67.525 171.125 ;
        RECT 67.700 170.455 67.955 170.955 ;
        RECT 68.125 170.625 68.455 171.125 ;
        RECT 67.700 170.285 68.450 170.455 ;
        RECT 67.700 169.465 68.050 170.115 ;
        RECT 63.255 169.135 63.765 169.315 ;
        RECT 64.170 169.225 65.870 169.395 ;
        RECT 64.170 169.135 64.555 169.225 ;
        RECT 63.255 168.745 63.585 169.135 ;
        RECT 63.755 168.795 64.940 168.965 ;
        RECT 65.200 168.575 65.370 169.045 ;
        RECT 65.540 168.760 65.870 169.225 ;
        RECT 66.040 168.575 66.210 169.395 ;
        RECT 66.380 168.755 67.065 169.395 ;
        RECT 67.235 168.575 67.525 169.300 ;
        RECT 68.220 169.295 68.450 170.285 ;
        RECT 67.700 169.125 68.450 169.295 ;
        RECT 67.700 168.835 67.955 169.125 ;
        RECT 68.125 168.575 68.455 168.955 ;
        RECT 68.625 168.835 68.795 170.955 ;
        RECT 68.965 170.155 69.290 170.940 ;
        RECT 69.460 170.665 69.710 171.125 ;
        RECT 69.880 170.625 70.130 170.955 ;
        RECT 70.345 170.625 71.025 170.955 ;
        RECT 69.880 170.495 70.050 170.625 ;
        RECT 69.655 170.325 70.050 170.495 ;
        RECT 69.025 169.105 69.485 170.155 ;
        RECT 69.655 168.965 69.825 170.325 ;
        RECT 70.220 170.065 70.685 170.455 ;
        RECT 69.995 169.255 70.345 169.875 ;
        RECT 70.515 169.475 70.685 170.065 ;
        RECT 70.855 169.845 71.025 170.625 ;
        RECT 71.195 170.525 71.365 170.865 ;
        RECT 71.600 170.695 71.930 171.125 ;
        RECT 72.100 170.525 72.270 170.865 ;
        RECT 72.565 170.665 72.935 171.125 ;
        RECT 71.195 170.355 72.270 170.525 ;
        RECT 73.105 170.495 73.275 170.955 ;
        RECT 73.510 170.615 74.380 170.955 ;
        RECT 74.550 170.665 74.800 171.125 ;
        RECT 72.715 170.325 73.275 170.495 ;
        RECT 72.715 170.185 72.885 170.325 ;
        RECT 71.385 170.015 72.885 170.185 ;
        RECT 73.580 170.155 74.040 170.445 ;
        RECT 70.855 169.675 72.545 169.845 ;
        RECT 70.515 169.255 70.870 169.475 ;
        RECT 71.040 168.965 71.210 169.675 ;
        RECT 71.415 169.255 72.205 169.505 ;
        RECT 72.375 169.495 72.545 169.675 ;
        RECT 72.715 169.325 72.885 170.015 ;
        RECT 69.155 168.575 69.485 168.935 ;
        RECT 69.655 168.795 70.150 168.965 ;
        RECT 70.355 168.795 71.210 168.965 ;
        RECT 72.085 168.575 72.415 169.035 ;
        RECT 72.625 168.935 72.885 169.325 ;
        RECT 73.075 170.145 74.040 170.155 ;
        RECT 74.210 170.235 74.380 170.615 ;
        RECT 74.970 170.575 75.140 170.865 ;
        RECT 75.320 170.745 75.650 171.125 ;
        RECT 74.970 170.405 75.770 170.575 ;
        RECT 73.075 169.985 73.750 170.145 ;
        RECT 74.210 170.065 75.430 170.235 ;
        RECT 73.075 169.195 73.285 169.985 ;
        RECT 74.210 169.975 74.380 170.065 ;
        RECT 73.455 169.195 73.805 169.815 ;
        RECT 73.975 169.805 74.380 169.975 ;
        RECT 73.975 169.025 74.145 169.805 ;
        RECT 74.315 169.355 74.535 169.635 ;
        RECT 74.715 169.525 75.255 169.895 ;
        RECT 75.600 169.815 75.770 170.405 ;
        RECT 75.990 169.985 76.295 171.125 ;
        RECT 76.465 169.935 76.715 170.815 ;
        RECT 76.885 169.985 77.135 171.125 ;
        RECT 77.355 170.695 77.695 170.955 ;
        RECT 75.600 169.785 76.340 169.815 ;
        RECT 74.315 169.185 74.845 169.355 ;
        RECT 72.625 168.765 72.975 168.935 ;
        RECT 73.195 168.745 74.145 169.025 ;
        RECT 74.315 168.575 74.505 169.015 ;
        RECT 74.675 168.955 74.845 169.185 ;
        RECT 75.015 169.125 75.255 169.525 ;
        RECT 75.425 169.485 76.340 169.785 ;
        RECT 75.425 169.310 75.750 169.485 ;
        RECT 75.425 168.955 75.745 169.310 ;
        RECT 76.510 169.285 76.715 169.935 ;
        RECT 74.675 168.785 75.745 168.955 ;
        RECT 75.990 168.575 76.295 169.035 ;
        RECT 76.465 168.755 76.715 169.285 ;
        RECT 76.885 168.575 77.135 169.330 ;
        RECT 77.355 169.295 77.615 170.695 ;
        RECT 77.865 170.325 78.195 171.125 ;
        RECT 78.660 170.155 78.910 170.955 ;
        RECT 79.095 170.405 79.425 171.125 ;
        RECT 79.645 170.155 79.895 170.955 ;
        RECT 80.065 170.745 80.400 171.125 ;
        RECT 77.805 169.985 79.995 170.155 ;
        RECT 77.805 169.815 78.120 169.985 ;
        RECT 77.790 169.565 78.120 169.815 ;
        RECT 77.355 168.785 77.695 169.295 ;
        RECT 77.865 168.575 78.135 169.375 ;
        RECT 78.315 168.845 78.595 169.815 ;
        RECT 78.775 168.845 79.075 169.815 ;
        RECT 79.255 168.850 79.605 169.815 ;
        RECT 79.825 169.075 79.995 169.985 ;
        RECT 80.165 169.255 80.405 170.565 ;
        RECT 80.575 170.405 81.035 170.955 ;
        RECT 81.225 170.405 81.555 171.125 ;
        RECT 79.825 168.745 80.320 169.075 ;
        RECT 80.575 169.035 80.825 170.405 ;
        RECT 81.755 170.235 82.055 170.785 ;
        RECT 82.225 170.455 82.505 171.125 ;
        RECT 81.115 170.065 82.055 170.235 ;
        RECT 82.965 170.195 83.135 170.955 ;
        RECT 83.350 170.365 83.680 171.125 ;
        RECT 81.115 169.815 81.285 170.065 ;
        RECT 82.425 169.815 82.690 170.175 ;
        RECT 82.965 170.025 83.680 170.195 ;
        RECT 83.850 170.050 84.105 170.955 ;
        RECT 80.995 169.485 81.285 169.815 ;
        RECT 81.455 169.565 81.795 169.815 ;
        RECT 82.015 169.565 82.690 169.815 ;
        RECT 81.115 169.395 81.285 169.485 ;
        RECT 82.875 169.475 83.230 169.845 ;
        RECT 83.510 169.815 83.680 170.025 ;
        RECT 83.510 169.485 83.765 169.815 ;
        RECT 81.115 169.205 82.505 169.395 ;
        RECT 83.510 169.295 83.680 169.485 ;
        RECT 83.935 169.320 84.105 170.050 ;
        RECT 84.280 169.975 84.540 171.125 ;
        RECT 85.185 170.745 85.515 171.125 ;
        RECT 80.575 168.745 81.135 169.035 ;
        RECT 81.305 168.575 81.555 169.035 ;
        RECT 82.175 168.845 82.505 169.205 ;
        RECT 82.965 169.125 83.680 169.295 ;
        RECT 82.965 168.745 83.135 169.125 ;
        RECT 83.350 168.575 83.680 168.955 ;
        RECT 83.850 168.745 84.105 169.320 ;
        RECT 84.280 168.575 84.540 169.415 ;
        RECT 85.215 169.245 85.420 170.565 ;
        RECT 85.690 170.155 85.940 170.955 ;
        RECT 86.160 170.405 86.490 171.125 ;
        RECT 86.675 170.155 86.925 170.955 ;
        RECT 87.325 170.325 87.655 171.125 ;
        RECT 87.825 170.785 88.160 170.955 ;
        RECT 87.825 170.615 88.165 170.785 ;
        RECT 85.590 169.985 87.645 170.155 ;
        RECT 87.825 169.985 88.160 170.615 ;
        RECT 88.335 170.325 88.665 171.125 ;
        RECT 88.855 169.985 89.135 171.125 ;
        RECT 85.590 169.075 85.760 169.985 ;
        RECT 85.265 168.745 85.760 169.075 ;
        RECT 85.980 168.910 86.335 169.815 ;
        RECT 86.510 169.795 86.680 169.815 ;
        RECT 86.510 168.905 86.810 169.795 ;
        RECT 86.990 168.905 87.250 169.815 ;
        RECT 87.420 169.805 87.645 169.985 ;
        RECT 87.420 169.565 87.815 169.805 ;
        RECT 87.420 168.575 87.655 169.380 ;
        RECT 87.985 169.295 88.160 169.985 ;
        RECT 89.305 169.975 89.635 170.955 ;
        RECT 89.805 169.985 90.065 171.125 ;
        RECT 91.160 169.975 91.420 171.125 ;
        RECT 91.595 170.050 91.850 170.955 ;
        RECT 92.020 170.365 92.350 171.125 ;
        RECT 92.565 170.195 92.735 170.955 ;
        RECT 88.865 169.545 89.200 169.815 ;
        RECT 89.370 169.375 89.540 169.975 ;
        RECT 89.710 169.565 90.045 169.815 ;
        RECT 87.825 168.830 88.160 169.295 ;
        RECT 87.825 168.785 88.155 168.830 ;
        RECT 88.345 168.575 88.675 169.300 ;
        RECT 88.855 168.575 89.165 169.375 ;
        RECT 89.370 168.745 90.065 169.375 ;
        RECT 91.160 168.575 91.420 169.415 ;
        RECT 91.595 169.320 91.765 170.050 ;
        RECT 92.020 170.025 92.735 170.195 ;
        RECT 92.020 169.815 92.190 170.025 ;
        RECT 92.995 169.960 93.285 171.125 ;
        RECT 93.545 170.445 93.715 170.955 ;
        RECT 93.885 170.615 94.215 171.125 ;
        RECT 94.385 170.445 94.555 170.955 ;
        RECT 94.725 170.615 95.055 171.125 ;
        RECT 95.225 170.445 95.395 170.955 ;
        RECT 95.565 170.615 95.895 171.125 ;
        RECT 96.185 170.785 97.195 170.955 ;
        RECT 96.185 170.445 96.355 170.785 ;
        RECT 93.545 170.275 96.355 170.445 ;
        RECT 96.525 170.115 96.855 170.605 ;
        RECT 97.025 170.285 97.195 170.785 ;
        RECT 97.465 170.615 97.795 171.125 ;
        RECT 97.965 170.445 98.135 170.955 ;
        RECT 98.305 170.615 98.635 171.125 ;
        RECT 98.805 170.445 98.975 170.955 ;
        RECT 99.145 170.615 99.475 171.125 ;
        RECT 97.905 170.275 99.665 170.445 ;
        RECT 93.515 169.935 96.225 170.105 ;
        RECT 91.935 169.485 92.190 169.815 ;
        RECT 91.595 168.745 91.850 169.320 ;
        RECT 92.020 169.295 92.190 169.485 ;
        RECT 92.470 169.475 92.825 169.845 ;
        RECT 93.520 169.565 93.895 169.935 ;
        RECT 94.095 169.565 94.425 169.735 ;
        RECT 94.725 169.565 95.075 169.765 ;
        RECT 95.355 169.565 95.685 169.765 ;
        RECT 95.895 169.565 96.225 169.935 ;
        RECT 96.525 169.945 97.765 170.115 ;
        RECT 94.175 169.395 94.345 169.565 ;
        RECT 95.355 169.395 95.540 169.565 ;
        RECT 92.020 169.125 92.735 169.295 ;
        RECT 92.020 168.575 92.350 168.955 ;
        RECT 92.565 168.745 92.735 169.125 ;
        RECT 92.995 168.575 93.285 169.300 ;
        RECT 93.545 168.575 93.715 169.395 ;
        RECT 94.175 169.225 95.540 169.395 ;
        RECT 96.525 169.360 96.715 169.945 ;
        RECT 97.595 169.815 97.765 169.945 ;
        RECT 96.945 169.565 97.400 169.775 ;
        RECT 95.720 169.295 96.715 169.360 ;
        RECT 95.720 169.190 96.855 169.295 ;
        RECT 97.185 169.235 97.400 169.565 ;
        RECT 97.595 169.485 99.305 169.815 ;
        RECT 99.495 169.315 99.665 170.275 ;
        RECT 99.985 170.155 100.155 170.955 ;
        RECT 100.445 170.495 100.695 170.915 ;
        RECT 100.885 170.665 101.215 171.125 ;
        RECT 101.425 170.495 101.675 170.915 ;
        RECT 100.385 170.325 101.675 170.495 ;
        RECT 101.845 170.325 102.095 171.125 ;
        RECT 102.265 170.495 102.435 170.955 ;
        RECT 102.645 170.665 102.895 171.125 ;
        RECT 102.265 170.325 102.940 170.495 ;
        RECT 103.125 170.325 103.455 171.125 ;
        RECT 103.635 170.785 105.065 170.955 ;
        RECT 99.985 169.985 102.475 170.155 ;
        RECT 95.720 169.055 95.890 169.190 ;
        RECT 94.725 168.885 95.890 169.055 ;
        RECT 96.070 168.575 96.355 169.020 ;
        RECT 96.525 168.785 96.855 169.190 ;
        RECT 97.875 169.145 99.665 169.315 ;
        RECT 99.940 169.245 100.135 169.815 ;
        RECT 97.105 168.575 97.635 169.055 ;
        RECT 98.305 168.575 98.635 168.975 ;
        RECT 99.145 168.575 99.475 168.975 ;
        RECT 99.895 168.575 100.155 169.055 ;
        RECT 100.325 168.995 100.495 169.985 ;
        RECT 100.675 169.360 100.845 169.815 ;
        RECT 101.235 169.735 101.405 169.750 ;
        RECT 101.075 169.565 101.405 169.735 ;
        RECT 100.675 169.190 101.065 169.360 ;
        RECT 100.325 168.825 100.655 168.995 ;
        RECT 100.855 168.905 101.065 169.190 ;
        RECT 101.235 169.355 101.405 169.565 ;
        RECT 101.635 169.485 101.965 169.815 ;
        RECT 102.305 169.735 102.475 169.985 ;
        RECT 102.145 169.565 102.475 169.735 ;
        RECT 101.235 169.185 101.500 169.355 ;
        RECT 101.760 169.250 101.965 169.485 ;
        RECT 102.685 169.375 102.940 170.325 ;
        RECT 103.635 170.155 103.885 170.785 ;
        RECT 101.330 169.085 101.500 169.185 ;
        RECT 102.265 169.205 102.940 169.375 ;
        RECT 103.115 169.985 103.885 170.155 ;
        RECT 103.115 169.315 103.285 169.985 ;
        RECT 103.455 169.485 103.860 169.815 ;
        RECT 104.075 169.485 104.325 170.615 ;
        RECT 104.525 169.815 104.725 170.615 ;
        RECT 104.895 170.105 105.065 170.785 ;
        RECT 105.235 170.275 105.550 171.125 ;
        RECT 105.725 170.325 106.165 170.955 ;
        RECT 104.895 169.935 105.685 170.105 ;
        RECT 104.525 169.485 104.770 169.815 ;
        RECT 104.955 169.485 105.345 169.765 ;
        RECT 105.515 169.485 105.685 169.935 ;
        RECT 105.855 169.315 106.165 170.325 ;
        RECT 106.795 169.935 107.055 171.125 ;
        RECT 107.225 170.105 107.555 170.955 ;
        RECT 107.725 170.325 107.895 171.125 ;
        RECT 108.065 170.105 108.395 170.955 ;
        RECT 108.565 170.325 108.815 171.125 ;
        RECT 109.005 170.785 110.935 170.955 ;
        RECT 109.005 170.275 109.255 170.785 ;
        RECT 109.425 170.105 109.755 170.615 ;
        RECT 109.925 170.275 110.095 170.785 ;
        RECT 110.265 170.105 110.595 170.615 ;
        RECT 107.225 169.935 110.595 170.105 ;
        RECT 110.765 170.105 110.935 170.785 ;
        RECT 111.105 170.785 114.395 170.955 ;
        RECT 111.105 170.275 111.355 170.785 ;
        RECT 111.525 170.105 111.855 170.615 ;
        RECT 112.025 170.275 112.195 170.785 ;
        RECT 112.365 170.105 112.695 170.615 ;
        RECT 110.765 169.935 112.695 170.105 ;
        RECT 112.885 170.105 113.215 170.615 ;
        RECT 113.385 170.275 113.555 170.785 ;
        RECT 113.725 170.105 114.055 170.615 ;
        RECT 114.225 170.275 114.395 170.785 ;
        RECT 114.565 170.105 114.895 170.955 ;
        RECT 115.065 170.325 115.235 171.125 ;
        RECT 115.405 170.105 115.735 170.955 ;
        RECT 115.905 170.325 116.075 171.125 ;
        RECT 116.245 170.105 116.575 170.955 ;
        RECT 112.885 169.935 116.575 170.105 ;
        RECT 116.915 170.035 118.585 171.125 ;
        RECT 106.815 169.565 108.410 169.765 ;
        RECT 108.580 169.395 108.870 169.935 ;
        RECT 109.060 169.565 110.730 169.765 ;
        RECT 111.020 169.565 112.690 169.765 ;
        RECT 112.880 169.565 114.650 169.765 ;
        RECT 114.865 169.565 116.745 169.765 ;
        RECT 101.330 168.915 101.505 169.085 ;
        RECT 101.845 168.955 102.015 169.035 ;
        RECT 101.330 168.890 101.500 168.915 ;
        RECT 100.325 168.745 100.570 168.825 ;
        RECT 101.745 168.575 102.075 168.955 ;
        RECT 102.265 168.745 102.435 169.205 ;
        RECT 102.685 168.575 102.940 169.035 ;
        RECT 103.115 168.745 103.605 169.315 ;
        RECT 103.775 169.145 104.935 169.315 ;
        RECT 103.775 168.745 104.005 169.145 ;
        RECT 104.175 168.575 104.595 168.975 ;
        RECT 104.765 168.745 104.935 169.145 ;
        RECT 105.105 168.575 105.555 169.315 ;
        RECT 105.725 168.755 106.165 169.315 ;
        RECT 106.795 168.955 107.055 169.395 ;
        RECT 107.225 169.125 108.870 169.395 ;
        RECT 109.060 169.225 116.575 169.395 ;
        RECT 109.060 168.955 109.335 169.225 ;
        RECT 106.795 168.745 109.335 168.955 ;
        RECT 109.505 168.575 109.675 169.035 ;
        RECT 109.845 168.745 110.175 169.225 ;
        RECT 110.345 168.575 110.515 169.035 ;
        RECT 110.685 168.745 111.015 169.225 ;
        RECT 111.185 168.575 111.355 169.035 ;
        RECT 111.525 168.745 111.855 169.225 ;
        RECT 112.025 168.575 112.195 169.035 ;
        RECT 112.365 168.745 112.695 169.225 ;
        RECT 112.885 168.750 113.215 169.225 ;
        RECT 113.385 168.575 113.555 169.035 ;
        RECT 113.725 168.750 114.055 169.225 ;
        RECT 114.225 168.575 114.395 169.035 ;
        RECT 114.565 168.750 114.895 169.225 ;
        RECT 115.065 168.575 115.235 169.035 ;
        RECT 115.405 168.750 115.735 169.225 ;
        RECT 115.905 168.575 116.075 169.035 ;
        RECT 116.245 168.750 116.575 169.225 ;
        RECT 116.915 169.345 117.665 169.865 ;
        RECT 117.835 169.515 118.585 170.035 ;
        RECT 118.755 169.960 119.045 171.125 ;
        RECT 119.270 170.255 119.555 171.125 ;
        RECT 119.725 170.495 119.985 170.955 ;
        RECT 120.160 170.665 120.415 171.125 ;
        RECT 120.585 170.495 120.845 170.955 ;
        RECT 119.725 170.325 120.845 170.495 ;
        RECT 121.015 170.325 121.325 171.125 ;
        RECT 119.725 170.075 119.985 170.325 ;
        RECT 121.495 170.155 121.805 170.955 ;
        RECT 119.230 169.905 119.985 170.075 ;
        RECT 120.775 169.985 121.805 170.155 ;
        RECT 119.230 169.395 119.635 169.905 ;
        RECT 120.775 169.735 120.945 169.985 ;
        RECT 119.805 169.565 120.945 169.735 ;
        RECT 116.915 168.575 118.585 169.345 ;
        RECT 118.755 168.575 119.045 169.300 ;
        RECT 119.230 169.225 120.880 169.395 ;
        RECT 121.115 169.245 121.465 169.815 ;
        RECT 119.275 168.575 119.555 169.055 ;
        RECT 119.725 168.835 119.985 169.225 ;
        RECT 120.160 168.575 120.415 169.055 ;
        RECT 120.585 168.835 120.880 169.225 ;
        RECT 121.635 169.075 121.805 169.985 ;
        RECT 121.060 168.575 121.335 169.055 ;
        RECT 121.505 168.745 121.805 169.075 ;
        RECT 121.975 170.155 122.285 170.955 ;
        RECT 122.455 170.325 122.765 171.125 ;
        RECT 122.935 170.495 123.195 170.955 ;
        RECT 123.365 170.665 123.620 171.125 ;
        RECT 123.795 170.495 124.055 170.955 ;
        RECT 122.935 170.325 124.055 170.495 ;
        RECT 121.975 169.985 123.005 170.155 ;
        RECT 121.975 169.075 122.145 169.985 ;
        RECT 122.315 169.245 122.665 169.815 ;
        RECT 122.835 169.735 123.005 169.985 ;
        RECT 123.795 170.075 124.055 170.325 ;
        RECT 124.225 170.255 124.510 171.125 ;
        RECT 124.825 170.455 124.995 170.955 ;
        RECT 125.165 170.625 125.495 171.125 ;
        RECT 124.825 170.285 125.490 170.455 ;
        RECT 123.795 169.905 124.550 170.075 ;
        RECT 122.835 169.565 123.975 169.735 ;
        RECT 124.145 169.395 124.550 169.905 ;
        RECT 124.740 169.465 125.090 170.115 ;
        RECT 122.900 169.225 124.550 169.395 ;
        RECT 125.260 169.295 125.490 170.285 ;
        RECT 121.975 168.745 122.275 169.075 ;
        RECT 122.445 168.575 122.720 169.055 ;
        RECT 122.900 168.835 123.195 169.225 ;
        RECT 123.365 168.575 123.620 169.055 ;
        RECT 123.795 168.835 124.055 169.225 ;
        RECT 124.825 169.125 125.490 169.295 ;
        RECT 124.225 168.575 124.505 169.055 ;
        RECT 124.825 168.835 124.995 169.125 ;
        RECT 125.165 168.575 125.495 168.955 ;
        RECT 125.665 168.835 125.890 170.955 ;
        RECT 126.105 170.625 126.435 171.125 ;
        RECT 126.605 170.455 126.775 170.955 ;
        RECT 127.010 170.740 127.840 170.910 ;
        RECT 128.080 170.745 128.460 171.125 ;
        RECT 126.080 170.285 126.775 170.455 ;
        RECT 126.080 169.315 126.250 170.285 ;
        RECT 126.420 169.495 126.830 170.115 ;
        RECT 127.000 170.065 127.500 170.445 ;
        RECT 126.080 169.125 126.775 169.315 ;
        RECT 127.000 169.195 127.220 170.065 ;
        RECT 127.670 169.895 127.840 170.740 ;
        RECT 128.640 170.575 128.810 170.865 ;
        RECT 128.980 170.745 129.310 171.125 ;
        RECT 129.780 170.655 130.410 170.905 ;
        RECT 130.590 170.745 131.010 171.125 ;
        RECT 130.240 170.575 130.410 170.655 ;
        RECT 131.210 170.575 131.450 170.865 ;
        RECT 128.010 170.325 129.380 170.575 ;
        RECT 128.010 170.065 128.260 170.325 ;
        RECT 128.770 169.895 129.020 170.055 ;
        RECT 127.670 169.725 129.020 169.895 ;
        RECT 127.670 169.685 128.090 169.725 ;
        RECT 127.400 169.135 127.750 169.505 ;
        RECT 126.105 168.575 126.435 168.955 ;
        RECT 126.605 168.795 126.775 169.125 ;
        RECT 127.920 168.955 128.090 169.685 ;
        RECT 129.190 169.555 129.380 170.325 ;
        RECT 128.260 169.225 128.670 169.555 ;
        RECT 128.960 169.215 129.380 169.555 ;
        RECT 129.550 170.145 130.070 170.455 ;
        RECT 130.240 170.405 131.450 170.575 ;
        RECT 131.680 170.435 132.010 171.125 ;
        RECT 129.550 169.385 129.720 170.145 ;
        RECT 129.890 169.555 130.070 169.965 ;
        RECT 130.240 169.895 130.410 170.405 ;
        RECT 132.180 170.255 132.350 170.865 ;
        RECT 132.620 170.405 132.950 170.915 ;
        RECT 132.180 170.235 132.500 170.255 ;
        RECT 130.580 170.065 132.500 170.235 ;
        RECT 130.240 169.725 132.140 169.895 ;
        RECT 130.470 169.385 130.800 169.505 ;
        RECT 129.550 169.215 130.800 169.385 ;
        RECT 127.075 168.755 128.090 168.955 ;
        RECT 128.260 168.575 128.670 169.015 ;
        RECT 128.960 168.785 129.210 169.215 ;
        RECT 129.410 168.575 129.730 169.035 ;
        RECT 130.970 168.965 131.140 169.725 ;
        RECT 131.810 169.665 132.140 169.725 ;
        RECT 131.330 169.495 131.660 169.555 ;
        RECT 131.330 169.225 131.990 169.495 ;
        RECT 132.310 169.170 132.500 170.065 ;
        RECT 130.290 168.795 131.140 168.965 ;
        RECT 131.340 168.575 132.000 169.055 ;
        RECT 132.180 168.840 132.500 169.170 ;
        RECT 132.700 169.815 132.950 170.405 ;
        RECT 133.130 170.325 133.415 171.125 ;
        RECT 133.595 170.785 133.850 170.815 ;
        RECT 133.595 170.615 133.935 170.785 ;
        RECT 133.595 170.145 133.850 170.615 ;
        RECT 134.400 170.455 134.655 170.955 ;
        RECT 134.825 170.625 135.155 171.125 ;
        RECT 134.400 170.285 135.150 170.455 ;
        RECT 132.700 169.485 133.500 169.815 ;
        RECT 132.700 168.835 132.950 169.485 ;
        RECT 133.670 169.285 133.850 170.145 ;
        RECT 134.400 169.465 134.750 170.115 ;
        RECT 134.920 169.295 135.150 170.285 ;
        RECT 133.130 168.575 133.415 169.035 ;
        RECT 133.595 168.755 133.850 169.285 ;
        RECT 134.400 169.125 135.150 169.295 ;
        RECT 134.400 168.835 134.655 169.125 ;
        RECT 134.825 168.575 135.155 168.955 ;
        RECT 135.325 168.835 135.495 170.955 ;
        RECT 135.665 170.155 135.990 170.940 ;
        RECT 136.160 170.665 136.410 171.125 ;
        RECT 136.580 170.625 136.830 170.955 ;
        RECT 137.045 170.625 137.725 170.955 ;
        RECT 136.580 170.495 136.750 170.625 ;
        RECT 136.355 170.325 136.750 170.495 ;
        RECT 135.725 169.105 136.185 170.155 ;
        RECT 136.355 168.965 136.525 170.325 ;
        RECT 136.920 170.065 137.385 170.455 ;
        RECT 136.695 169.255 137.045 169.875 ;
        RECT 137.215 169.475 137.385 170.065 ;
        RECT 137.555 169.845 137.725 170.625 ;
        RECT 137.895 170.525 138.065 170.865 ;
        RECT 138.300 170.695 138.630 171.125 ;
        RECT 138.800 170.525 138.970 170.865 ;
        RECT 139.265 170.665 139.635 171.125 ;
        RECT 137.895 170.355 138.970 170.525 ;
        RECT 139.805 170.495 139.975 170.955 ;
        RECT 140.210 170.615 141.080 170.955 ;
        RECT 141.250 170.665 141.500 171.125 ;
        RECT 139.415 170.325 139.975 170.495 ;
        RECT 139.415 170.185 139.585 170.325 ;
        RECT 138.085 170.015 139.585 170.185 ;
        RECT 140.280 170.155 140.740 170.445 ;
        RECT 137.555 169.675 139.245 169.845 ;
        RECT 137.215 169.255 137.570 169.475 ;
        RECT 137.740 168.965 137.910 169.675 ;
        RECT 138.115 169.255 138.905 169.505 ;
        RECT 139.075 169.495 139.245 169.675 ;
        RECT 139.415 169.325 139.585 170.015 ;
        RECT 135.855 168.575 136.185 168.935 ;
        RECT 136.355 168.795 136.850 168.965 ;
        RECT 137.055 168.795 137.910 168.965 ;
        RECT 138.785 168.575 139.115 169.035 ;
        RECT 139.325 168.935 139.585 169.325 ;
        RECT 139.775 170.145 140.740 170.155 ;
        RECT 140.910 170.235 141.080 170.615 ;
        RECT 141.670 170.575 141.840 170.865 ;
        RECT 142.020 170.745 142.350 171.125 ;
        RECT 141.670 170.405 142.470 170.575 ;
        RECT 139.775 169.985 140.450 170.145 ;
        RECT 140.910 170.065 142.130 170.235 ;
        RECT 139.775 169.195 139.985 169.985 ;
        RECT 140.910 169.975 141.080 170.065 ;
        RECT 140.155 169.195 140.505 169.815 ;
        RECT 140.675 169.805 141.080 169.975 ;
        RECT 140.675 169.025 140.845 169.805 ;
        RECT 141.015 169.355 141.235 169.635 ;
        RECT 141.415 169.525 141.955 169.895 ;
        RECT 142.300 169.815 142.470 170.405 ;
        RECT 142.690 169.985 142.995 171.125 ;
        RECT 143.165 169.935 143.415 170.815 ;
        RECT 143.585 169.985 143.835 171.125 ;
        RECT 144.515 169.960 144.805 171.125 ;
        RECT 144.975 170.690 150.320 171.125 ;
        RECT 150.495 170.690 155.840 171.125 ;
        RECT 142.300 169.785 143.040 169.815 ;
        RECT 141.015 169.185 141.545 169.355 ;
        RECT 139.325 168.765 139.675 168.935 ;
        RECT 139.895 168.745 140.845 169.025 ;
        RECT 141.015 168.575 141.205 169.015 ;
        RECT 141.375 168.955 141.545 169.185 ;
        RECT 141.715 169.125 141.955 169.525 ;
        RECT 142.125 169.485 143.040 169.785 ;
        RECT 142.125 169.310 142.450 169.485 ;
        RECT 142.125 168.955 142.445 169.310 ;
        RECT 143.210 169.285 143.415 169.935 ;
        RECT 141.375 168.785 142.445 168.955 ;
        RECT 142.690 168.575 142.995 169.035 ;
        RECT 143.165 168.755 143.415 169.285 ;
        RECT 143.585 168.575 143.835 169.330 ;
        RECT 144.515 168.575 144.805 169.300 ;
        RECT 146.560 169.120 146.900 169.950 ;
        RECT 148.380 169.440 148.730 170.690 ;
        RECT 152.080 169.120 152.420 169.950 ;
        RECT 153.900 169.440 154.250 170.690 ;
        RECT 156.935 170.035 158.145 171.125 ;
        RECT 156.935 169.495 157.455 170.035 ;
        RECT 157.625 169.325 158.145 169.865 ;
        RECT 144.975 168.575 150.320 169.120 ;
        RECT 150.495 168.575 155.840 169.120 ;
        RECT 156.935 168.575 158.145 169.325 ;
        RECT 2.750 168.405 158.230 168.575 ;
        RECT 2.835 167.655 4.045 168.405 ;
        RECT 2.835 167.115 3.355 167.655 ;
        RECT 4.215 167.635 5.885 168.405 ;
        RECT 6.055 167.730 6.315 168.235 ;
        RECT 6.495 168.025 6.825 168.405 ;
        RECT 7.005 167.855 7.175 168.235 ;
        RECT 3.525 166.945 4.045 167.485 ;
        RECT 4.215 167.115 4.965 167.635 ;
        RECT 5.135 166.945 5.885 167.465 ;
        RECT 2.835 165.855 4.045 166.945 ;
        RECT 4.215 165.855 5.885 166.945 ;
        RECT 6.055 166.930 6.225 167.730 ;
        RECT 6.510 167.685 7.175 167.855 ;
        RECT 6.510 167.430 6.680 167.685 ;
        RECT 8.360 167.665 8.615 168.235 ;
        RECT 8.785 168.005 9.115 168.405 ;
        RECT 9.540 167.870 10.070 168.235 ;
        RECT 9.540 167.835 9.715 167.870 ;
        RECT 8.785 167.665 9.715 167.835 ;
        RECT 6.395 167.100 6.680 167.430 ;
        RECT 6.915 167.135 7.245 167.505 ;
        RECT 6.510 166.955 6.680 167.100 ;
        RECT 8.360 166.995 8.530 167.665 ;
        RECT 8.785 167.495 8.955 167.665 ;
        RECT 8.700 167.165 8.955 167.495 ;
        RECT 9.180 167.165 9.375 167.495 ;
        RECT 6.055 166.025 6.325 166.930 ;
        RECT 6.510 166.785 7.175 166.955 ;
        RECT 6.495 165.855 6.825 166.615 ;
        RECT 7.005 166.025 7.175 166.785 ;
        RECT 8.360 166.025 8.695 166.995 ;
        RECT 8.865 165.855 9.035 166.995 ;
        RECT 9.205 166.195 9.375 167.165 ;
        RECT 9.545 166.535 9.715 167.665 ;
        RECT 9.885 166.875 10.055 167.675 ;
        RECT 10.260 167.385 10.535 168.235 ;
        RECT 10.255 167.215 10.535 167.385 ;
        RECT 10.260 167.075 10.535 167.215 ;
        RECT 10.705 166.875 10.895 168.235 ;
        RECT 11.075 167.870 11.585 168.405 ;
        RECT 11.805 167.595 12.050 168.200 ;
        RECT 12.495 167.665 12.880 168.235 ;
        RECT 13.050 167.945 13.375 168.405 ;
        RECT 13.895 167.775 14.175 168.235 ;
        RECT 11.095 167.425 12.325 167.595 ;
        RECT 9.885 166.705 10.895 166.875 ;
        RECT 11.065 166.860 11.815 167.050 ;
        RECT 9.545 166.365 10.670 166.535 ;
        RECT 11.065 166.195 11.235 166.860 ;
        RECT 11.985 166.615 12.325 167.425 ;
        RECT 9.205 166.025 11.235 166.195 ;
        RECT 11.405 165.855 11.575 166.615 ;
        RECT 11.810 166.205 12.325 166.615 ;
        RECT 12.495 166.995 12.775 167.665 ;
        RECT 13.050 167.605 14.175 167.775 ;
        RECT 13.050 167.495 13.500 167.605 ;
        RECT 12.945 167.165 13.500 167.495 ;
        RECT 14.365 167.435 14.765 168.235 ;
        RECT 15.165 167.945 15.435 168.405 ;
        RECT 15.605 167.775 15.890 168.235 ;
        RECT 12.495 166.025 12.880 166.995 ;
        RECT 13.050 166.705 13.500 167.165 ;
        RECT 13.670 166.875 14.765 167.435 ;
        RECT 13.050 166.485 14.175 166.705 ;
        RECT 13.050 165.855 13.375 166.315 ;
        RECT 13.895 166.025 14.175 166.485 ;
        RECT 14.365 166.025 14.765 166.875 ;
        RECT 14.935 167.605 15.890 167.775 ;
        RECT 16.180 167.665 16.435 168.235 ;
        RECT 16.605 168.005 16.935 168.405 ;
        RECT 17.360 167.870 17.890 168.235 ;
        RECT 17.360 167.835 17.535 167.870 ;
        RECT 16.605 167.665 17.535 167.835 ;
        RECT 18.080 167.725 18.355 168.235 ;
        RECT 14.935 166.705 15.145 167.605 ;
        RECT 15.315 166.875 16.005 167.435 ;
        RECT 16.180 166.995 16.350 167.665 ;
        RECT 16.605 167.495 16.775 167.665 ;
        RECT 16.520 167.165 16.775 167.495 ;
        RECT 17.000 167.165 17.195 167.495 ;
        RECT 14.935 166.485 15.890 166.705 ;
        RECT 15.165 165.855 15.435 166.315 ;
        RECT 15.605 166.025 15.890 166.485 ;
        RECT 16.180 166.025 16.515 166.995 ;
        RECT 16.685 165.855 16.855 166.995 ;
        RECT 17.025 166.195 17.195 167.165 ;
        RECT 17.365 166.535 17.535 167.665 ;
        RECT 17.705 166.875 17.875 167.675 ;
        RECT 18.075 167.555 18.355 167.725 ;
        RECT 18.080 167.075 18.355 167.555 ;
        RECT 18.525 166.875 18.715 168.235 ;
        RECT 18.895 167.870 19.405 168.405 ;
        RECT 19.625 167.595 19.870 168.200 ;
        RECT 20.315 167.635 23.825 168.405 ;
        RECT 24.085 167.755 24.255 168.235 ;
        RECT 24.425 167.925 24.755 168.405 ;
        RECT 24.980 167.985 26.515 168.235 ;
        RECT 24.980 167.755 25.150 167.985 ;
        RECT 18.915 167.425 20.145 167.595 ;
        RECT 17.705 166.705 18.715 166.875 ;
        RECT 18.885 166.860 19.635 167.050 ;
        RECT 17.365 166.365 18.490 166.535 ;
        RECT 18.885 166.195 19.055 166.860 ;
        RECT 19.805 166.615 20.145 167.425 ;
        RECT 20.315 167.115 21.965 167.635 ;
        RECT 24.085 167.585 25.150 167.755 ;
        RECT 22.135 166.945 23.825 167.465 ;
        RECT 25.330 167.415 25.610 167.815 ;
        RECT 24.000 167.205 24.350 167.415 ;
        RECT 24.520 167.215 24.965 167.415 ;
        RECT 25.135 167.215 25.610 167.415 ;
        RECT 25.880 167.415 26.165 167.815 ;
        RECT 26.345 167.755 26.515 167.985 ;
        RECT 26.685 167.925 27.015 168.405 ;
        RECT 27.230 167.905 27.485 168.235 ;
        RECT 27.300 167.825 27.485 167.905 ;
        RECT 26.345 167.585 27.145 167.755 ;
        RECT 25.880 167.215 26.210 167.415 ;
        RECT 26.380 167.215 26.745 167.415 ;
        RECT 26.975 167.035 27.145 167.585 ;
        RECT 17.025 166.025 19.055 166.195 ;
        RECT 19.225 165.855 19.395 166.615 ;
        RECT 19.630 166.205 20.145 166.615 ;
        RECT 20.315 165.855 23.825 166.945 ;
        RECT 24.085 166.865 27.145 167.035 ;
        RECT 24.085 166.025 24.255 166.865 ;
        RECT 27.315 166.705 27.485 167.825 ;
        RECT 28.595 167.680 28.885 168.405 ;
        RECT 29.060 167.855 29.315 168.145 ;
        RECT 29.485 168.025 29.815 168.405 ;
        RECT 29.060 167.685 29.810 167.855 ;
        RECT 27.275 166.695 27.485 166.705 ;
        RECT 24.425 166.195 24.755 166.695 ;
        RECT 24.925 166.455 26.560 166.695 ;
        RECT 24.925 166.365 25.155 166.455 ;
        RECT 25.265 166.195 25.595 166.235 ;
        RECT 24.425 166.025 25.595 166.195 ;
        RECT 25.785 165.855 26.140 166.275 ;
        RECT 26.310 166.025 26.560 166.455 ;
        RECT 26.730 165.855 27.060 166.615 ;
        RECT 27.230 166.025 27.485 166.695 ;
        RECT 28.595 165.855 28.885 167.020 ;
        RECT 29.060 166.865 29.410 167.515 ;
        RECT 29.580 166.695 29.810 167.685 ;
        RECT 29.060 166.525 29.810 166.695 ;
        RECT 29.060 166.025 29.315 166.525 ;
        RECT 29.485 165.855 29.815 166.355 ;
        RECT 29.985 166.025 30.155 168.145 ;
        RECT 30.515 168.045 30.845 168.405 ;
        RECT 31.015 168.015 31.510 168.185 ;
        RECT 31.715 168.015 32.570 168.185 ;
        RECT 30.385 166.825 30.845 167.875 ;
        RECT 30.325 166.040 30.650 166.825 ;
        RECT 31.015 166.655 31.185 168.015 ;
        RECT 31.355 167.105 31.705 167.725 ;
        RECT 31.875 167.505 32.230 167.725 ;
        RECT 31.875 166.915 32.045 167.505 ;
        RECT 32.400 167.305 32.570 168.015 ;
        RECT 33.445 167.945 33.775 168.405 ;
        RECT 33.985 168.045 34.335 168.215 ;
        RECT 32.775 167.475 33.565 167.725 ;
        RECT 33.985 167.655 34.245 168.045 ;
        RECT 34.555 167.955 35.505 168.235 ;
        RECT 35.675 167.965 35.865 168.405 ;
        RECT 36.035 168.025 37.105 168.195 ;
        RECT 33.735 167.305 33.905 167.485 ;
        RECT 31.015 166.485 31.410 166.655 ;
        RECT 31.580 166.525 32.045 166.915 ;
        RECT 32.215 167.135 33.905 167.305 ;
        RECT 31.240 166.355 31.410 166.485 ;
        RECT 32.215 166.355 32.385 167.135 ;
        RECT 34.075 166.965 34.245 167.655 ;
        RECT 32.745 166.795 34.245 166.965 ;
        RECT 34.435 166.995 34.645 167.785 ;
        RECT 34.815 167.165 35.165 167.785 ;
        RECT 35.335 167.175 35.505 167.955 ;
        RECT 36.035 167.795 36.205 168.025 ;
        RECT 35.675 167.625 36.205 167.795 ;
        RECT 35.675 167.345 35.895 167.625 ;
        RECT 36.375 167.455 36.615 167.855 ;
        RECT 35.335 167.005 35.740 167.175 ;
        RECT 36.075 167.085 36.615 167.455 ;
        RECT 36.785 167.670 37.105 168.025 ;
        RECT 37.350 167.945 37.655 168.405 ;
        RECT 37.825 167.695 38.080 168.225 ;
        RECT 36.785 167.495 37.110 167.670 ;
        RECT 36.785 167.195 37.700 167.495 ;
        RECT 36.960 167.165 37.700 167.195 ;
        RECT 34.435 166.835 35.110 166.995 ;
        RECT 35.570 166.915 35.740 167.005 ;
        RECT 34.435 166.825 35.400 166.835 ;
        RECT 34.075 166.655 34.245 166.795 ;
        RECT 30.820 165.855 31.070 166.315 ;
        RECT 31.240 166.025 31.490 166.355 ;
        RECT 31.705 166.025 32.385 166.355 ;
        RECT 32.555 166.455 33.630 166.625 ;
        RECT 34.075 166.485 34.635 166.655 ;
        RECT 34.940 166.535 35.400 166.825 ;
        RECT 35.570 166.745 36.790 166.915 ;
        RECT 32.555 166.115 32.725 166.455 ;
        RECT 32.960 165.855 33.290 166.285 ;
        RECT 33.460 166.115 33.630 166.455 ;
        RECT 33.925 165.855 34.295 166.315 ;
        RECT 34.465 166.025 34.635 166.485 ;
        RECT 35.570 166.365 35.740 166.745 ;
        RECT 36.960 166.575 37.130 167.165 ;
        RECT 37.870 167.045 38.080 167.695 ;
        RECT 38.345 167.755 38.515 168.235 ;
        RECT 38.685 167.925 39.015 168.405 ;
        RECT 39.240 167.985 40.775 168.235 ;
        RECT 39.240 167.755 39.410 167.985 ;
        RECT 38.345 167.585 39.410 167.755 ;
        RECT 39.590 167.415 39.870 167.815 ;
        RECT 38.260 167.205 38.610 167.415 ;
        RECT 38.780 167.215 39.225 167.415 ;
        RECT 39.395 167.215 39.870 167.415 ;
        RECT 40.140 167.415 40.425 167.815 ;
        RECT 40.605 167.755 40.775 167.985 ;
        RECT 40.945 167.925 41.275 168.405 ;
        RECT 41.490 167.905 41.745 168.235 ;
        RECT 41.560 167.825 41.745 167.905 ;
        RECT 40.605 167.585 41.405 167.755 ;
        RECT 40.140 167.215 40.470 167.415 ;
        RECT 40.640 167.215 41.005 167.415 ;
        RECT 34.870 166.025 35.740 166.365 ;
        RECT 36.330 166.405 37.130 166.575 ;
        RECT 35.910 165.855 36.160 166.315 ;
        RECT 36.330 166.115 36.500 166.405 ;
        RECT 36.680 165.855 37.010 166.235 ;
        RECT 37.350 165.855 37.655 166.995 ;
        RECT 37.825 166.165 38.080 167.045 ;
        RECT 41.235 167.035 41.405 167.585 ;
        RECT 38.345 166.865 41.405 167.035 ;
        RECT 38.345 166.025 38.515 166.865 ;
        RECT 41.575 166.695 41.745 167.825 ;
        RECT 38.685 166.195 39.015 166.695 ;
        RECT 39.185 166.455 40.820 166.695 ;
        RECT 39.185 166.365 39.415 166.455 ;
        RECT 39.525 166.195 39.855 166.235 ;
        RECT 38.685 166.025 39.855 166.195 ;
        RECT 40.045 165.855 40.400 166.275 ;
        RECT 40.570 166.025 40.820 166.455 ;
        RECT 40.990 165.855 41.320 166.615 ;
        RECT 41.490 166.025 41.745 166.695 ;
        RECT 42.395 167.755 42.655 168.235 ;
        RECT 42.825 167.865 43.075 168.405 ;
        RECT 42.395 166.725 42.565 167.755 ;
        RECT 43.245 167.700 43.465 168.185 ;
        RECT 42.735 167.105 42.965 167.500 ;
        RECT 43.135 167.275 43.465 167.700 ;
        RECT 43.635 168.025 44.525 168.195 ;
        RECT 43.635 167.300 43.805 168.025 ;
        RECT 43.975 167.470 44.525 167.855 ;
        RECT 44.695 167.585 44.955 168.405 ;
        RECT 45.125 167.585 45.455 168.005 ;
        RECT 45.635 167.920 46.425 168.185 ;
        RECT 45.205 167.495 45.455 167.585 ;
        RECT 43.635 167.230 44.525 167.300 ;
        RECT 43.630 167.205 44.525 167.230 ;
        RECT 43.620 167.190 44.525 167.205 ;
        RECT 43.615 167.175 44.525 167.190 ;
        RECT 43.605 167.170 44.525 167.175 ;
        RECT 43.600 167.160 44.525 167.170 ;
        RECT 43.595 167.150 44.525 167.160 ;
        RECT 43.585 167.145 44.525 167.150 ;
        RECT 43.575 167.135 44.525 167.145 ;
        RECT 43.565 167.130 44.525 167.135 ;
        RECT 43.565 167.125 43.900 167.130 ;
        RECT 43.550 167.120 43.900 167.125 ;
        RECT 43.535 167.110 43.900 167.120 ;
        RECT 43.510 167.105 43.900 167.110 ;
        RECT 42.735 167.100 43.900 167.105 ;
        RECT 42.735 167.065 43.870 167.100 ;
        RECT 42.735 167.040 43.835 167.065 ;
        RECT 42.735 167.010 43.805 167.040 ;
        RECT 42.735 166.980 43.785 167.010 ;
        RECT 42.735 166.950 43.765 166.980 ;
        RECT 42.735 166.940 43.695 166.950 ;
        RECT 42.735 166.930 43.670 166.940 ;
        RECT 42.735 166.915 43.650 166.930 ;
        RECT 42.735 166.900 43.630 166.915 ;
        RECT 42.840 166.890 43.625 166.900 ;
        RECT 42.840 166.855 43.610 166.890 ;
        RECT 42.395 166.025 42.670 166.725 ;
        RECT 42.840 166.605 43.595 166.855 ;
        RECT 43.765 166.535 44.095 166.780 ;
        RECT 44.265 166.680 44.525 167.130 ;
        RECT 44.695 166.535 45.035 167.415 ;
        RECT 45.205 167.245 46.000 167.495 ;
        RECT 43.910 166.510 44.095 166.535 ;
        RECT 43.910 166.410 44.525 166.510 ;
        RECT 42.840 165.855 43.095 166.400 ;
        RECT 43.265 166.025 43.745 166.365 ;
        RECT 43.920 165.855 44.525 166.410 ;
        RECT 44.695 165.855 44.955 166.365 ;
        RECT 45.205 166.025 45.375 167.245 ;
        RECT 46.170 167.065 46.425 167.920 ;
        RECT 46.595 167.765 46.795 168.185 ;
        RECT 46.985 167.945 47.315 168.405 ;
        RECT 46.595 167.245 47.005 167.765 ;
        RECT 47.485 167.755 47.745 168.235 ;
        RECT 47.175 167.065 47.405 167.495 ;
        RECT 45.615 166.895 47.405 167.065 ;
        RECT 45.615 166.530 45.865 166.895 ;
        RECT 46.035 166.535 46.365 166.725 ;
        RECT 46.585 166.600 47.300 166.895 ;
        RECT 47.575 166.725 47.745 167.755 ;
        RECT 46.035 166.360 46.230 166.535 ;
        RECT 45.615 165.855 46.230 166.360 ;
        RECT 46.400 166.025 46.875 166.365 ;
        RECT 47.045 165.855 47.260 166.400 ;
        RECT 47.470 166.025 47.745 166.725 ;
        RECT 47.915 167.945 48.475 168.235 ;
        RECT 48.645 167.945 48.895 168.405 ;
        RECT 47.915 166.575 48.165 167.945 ;
        RECT 49.515 167.775 49.845 168.135 ;
        RECT 48.455 167.585 49.845 167.775 ;
        RECT 50.305 167.755 50.475 168.235 ;
        RECT 50.645 167.925 50.975 168.405 ;
        RECT 51.200 167.985 52.735 168.235 ;
        RECT 51.200 167.755 51.370 167.985 ;
        RECT 50.305 167.585 51.370 167.755 ;
        RECT 48.455 167.495 48.625 167.585 ;
        RECT 48.335 167.165 48.625 167.495 ;
        RECT 51.550 167.415 51.830 167.815 ;
        RECT 48.795 167.165 49.135 167.415 ;
        RECT 49.355 167.165 50.030 167.415 ;
        RECT 50.220 167.205 50.570 167.415 ;
        RECT 50.740 167.215 51.185 167.415 ;
        RECT 51.355 167.215 51.830 167.415 ;
        RECT 52.100 167.415 52.385 167.815 ;
        RECT 52.565 167.755 52.735 167.985 ;
        RECT 52.905 167.925 53.235 168.405 ;
        RECT 53.450 167.905 53.705 168.235 ;
        RECT 53.520 167.825 53.705 167.905 ;
        RECT 52.565 167.585 53.365 167.755 ;
        RECT 52.100 167.215 52.430 167.415 ;
        RECT 52.600 167.215 52.965 167.415 ;
        RECT 48.455 166.915 48.625 167.165 ;
        RECT 48.455 166.745 49.395 166.915 ;
        RECT 49.765 166.805 50.030 167.165 ;
        RECT 53.195 167.035 53.365 167.585 ;
        RECT 50.305 166.865 53.365 167.035 ;
        RECT 47.915 166.025 48.375 166.575 ;
        RECT 48.565 165.855 48.895 166.575 ;
        RECT 49.095 166.195 49.395 166.745 ;
        RECT 49.565 165.855 49.845 166.525 ;
        RECT 50.305 166.025 50.475 166.865 ;
        RECT 53.535 166.705 53.705 167.825 ;
        RECT 54.355 167.680 54.645 168.405 ;
        RECT 54.815 167.685 55.155 168.195 ;
        RECT 53.495 166.695 53.705 166.705 ;
        RECT 50.645 166.195 50.975 166.695 ;
        RECT 51.145 166.455 52.780 166.695 ;
        RECT 51.145 166.365 51.375 166.455 ;
        RECT 51.485 166.195 51.815 166.235 ;
        RECT 50.645 166.025 51.815 166.195 ;
        RECT 52.005 165.855 52.360 166.275 ;
        RECT 52.530 166.025 52.780 166.455 ;
        RECT 52.950 165.855 53.280 166.615 ;
        RECT 53.450 166.025 53.705 166.695 ;
        RECT 54.355 165.855 54.645 167.020 ;
        RECT 54.815 166.285 55.075 167.685 ;
        RECT 55.325 167.605 55.595 168.405 ;
        RECT 55.250 167.165 55.580 167.415 ;
        RECT 55.775 167.165 56.055 168.135 ;
        RECT 56.235 167.165 56.535 168.135 ;
        RECT 56.715 167.165 57.065 168.130 ;
        RECT 57.285 167.905 57.780 168.235 ;
        RECT 55.265 166.995 55.580 167.165 ;
        RECT 57.285 166.995 57.455 167.905 ;
        RECT 58.585 167.855 58.755 168.235 ;
        RECT 58.935 168.025 59.265 168.405 ;
        RECT 55.265 166.825 57.455 166.995 ;
        RECT 54.815 166.025 55.155 166.285 ;
        RECT 55.325 165.855 55.655 166.655 ;
        RECT 56.120 166.025 56.370 166.825 ;
        RECT 56.555 165.855 56.885 166.575 ;
        RECT 57.105 166.025 57.355 166.825 ;
        RECT 57.625 166.415 57.865 167.725 ;
        RECT 58.585 167.685 59.250 167.855 ;
        RECT 59.445 167.730 59.705 168.235 ;
        RECT 58.515 167.135 58.845 167.505 ;
        RECT 59.080 167.430 59.250 167.685 ;
        RECT 59.080 167.100 59.365 167.430 ;
        RECT 59.080 166.955 59.250 167.100 ;
        RECT 58.585 166.785 59.250 166.955 ;
        RECT 59.535 166.930 59.705 167.730 ;
        RECT 59.880 167.855 60.135 168.145 ;
        RECT 60.305 168.025 60.635 168.405 ;
        RECT 59.880 167.685 60.630 167.855 ;
        RECT 57.525 165.855 57.860 166.235 ;
        RECT 58.585 166.025 58.755 166.785 ;
        RECT 58.935 165.855 59.265 166.615 ;
        RECT 59.435 166.025 59.705 166.930 ;
        RECT 59.880 166.865 60.230 167.515 ;
        RECT 60.400 166.695 60.630 167.685 ;
        RECT 59.880 166.525 60.630 166.695 ;
        RECT 59.880 166.025 60.135 166.525 ;
        RECT 60.305 165.855 60.635 166.355 ;
        RECT 60.805 166.025 60.975 168.145 ;
        RECT 61.335 168.045 61.665 168.405 ;
        RECT 61.835 168.015 62.330 168.185 ;
        RECT 62.535 168.015 63.390 168.185 ;
        RECT 61.205 166.825 61.665 167.875 ;
        RECT 61.145 166.040 61.470 166.825 ;
        RECT 61.835 166.655 62.005 168.015 ;
        RECT 62.175 167.105 62.525 167.725 ;
        RECT 62.695 167.505 63.050 167.725 ;
        RECT 62.695 166.915 62.865 167.505 ;
        RECT 63.220 167.305 63.390 168.015 ;
        RECT 64.265 167.945 64.595 168.405 ;
        RECT 64.805 168.045 65.155 168.215 ;
        RECT 63.595 167.475 64.385 167.725 ;
        RECT 64.805 167.655 65.065 168.045 ;
        RECT 65.375 167.955 66.325 168.235 ;
        RECT 66.495 167.965 66.685 168.405 ;
        RECT 66.855 168.025 67.925 168.195 ;
        RECT 64.555 167.305 64.725 167.485 ;
        RECT 61.835 166.485 62.230 166.655 ;
        RECT 62.400 166.525 62.865 166.915 ;
        RECT 63.035 167.135 64.725 167.305 ;
        RECT 62.060 166.355 62.230 166.485 ;
        RECT 63.035 166.355 63.205 167.135 ;
        RECT 64.895 166.965 65.065 167.655 ;
        RECT 63.565 166.795 65.065 166.965 ;
        RECT 65.255 166.995 65.465 167.785 ;
        RECT 65.635 167.165 65.985 167.785 ;
        RECT 66.155 167.175 66.325 167.955 ;
        RECT 66.855 167.795 67.025 168.025 ;
        RECT 66.495 167.625 67.025 167.795 ;
        RECT 66.495 167.345 66.715 167.625 ;
        RECT 67.195 167.455 67.435 167.855 ;
        RECT 66.155 167.005 66.560 167.175 ;
        RECT 66.895 167.085 67.435 167.455 ;
        RECT 67.605 167.670 67.925 168.025 ;
        RECT 68.170 167.945 68.475 168.405 ;
        RECT 68.645 167.695 68.900 168.225 ;
        RECT 67.605 167.495 67.930 167.670 ;
        RECT 67.605 167.195 68.520 167.495 ;
        RECT 67.780 167.165 68.520 167.195 ;
        RECT 65.255 166.835 65.930 166.995 ;
        RECT 66.390 166.915 66.560 167.005 ;
        RECT 65.255 166.825 66.220 166.835 ;
        RECT 64.895 166.655 65.065 166.795 ;
        RECT 61.640 165.855 61.890 166.315 ;
        RECT 62.060 166.025 62.310 166.355 ;
        RECT 62.525 166.025 63.205 166.355 ;
        RECT 63.375 166.455 64.450 166.625 ;
        RECT 64.895 166.485 65.455 166.655 ;
        RECT 65.760 166.535 66.220 166.825 ;
        RECT 66.390 166.745 67.610 166.915 ;
        RECT 63.375 166.115 63.545 166.455 ;
        RECT 63.780 165.855 64.110 166.285 ;
        RECT 64.280 166.115 64.450 166.455 ;
        RECT 64.745 165.855 65.115 166.315 ;
        RECT 65.285 166.025 65.455 166.485 ;
        RECT 66.390 166.365 66.560 166.745 ;
        RECT 67.780 166.575 67.950 167.165 ;
        RECT 68.690 167.045 68.900 167.695 ;
        RECT 65.690 166.025 66.560 166.365 ;
        RECT 67.150 166.405 67.950 166.575 ;
        RECT 66.730 165.855 66.980 166.315 ;
        RECT 67.150 166.115 67.320 166.405 ;
        RECT 67.500 165.855 67.830 166.235 ;
        RECT 68.170 165.855 68.475 166.995 ;
        RECT 68.645 166.165 68.900 167.045 ;
        RECT 69.535 167.755 69.795 168.235 ;
        RECT 69.965 167.865 70.215 168.405 ;
        RECT 69.535 166.725 69.705 167.755 ;
        RECT 70.385 167.700 70.605 168.185 ;
        RECT 69.875 167.105 70.105 167.500 ;
        RECT 70.275 167.275 70.605 167.700 ;
        RECT 70.775 168.025 71.665 168.195 ;
        RECT 70.775 167.300 70.945 168.025 ;
        RECT 71.115 167.470 71.665 167.855 ;
        RECT 72.110 167.595 72.355 168.200 ;
        RECT 72.575 167.870 73.085 168.405 ;
        RECT 71.835 167.425 73.065 167.595 ;
        RECT 70.775 167.230 71.665 167.300 ;
        RECT 70.770 167.205 71.665 167.230 ;
        RECT 70.760 167.190 71.665 167.205 ;
        RECT 70.755 167.175 71.665 167.190 ;
        RECT 70.745 167.170 71.665 167.175 ;
        RECT 70.740 167.160 71.665 167.170 ;
        RECT 70.735 167.150 71.665 167.160 ;
        RECT 70.725 167.145 71.665 167.150 ;
        RECT 70.715 167.135 71.665 167.145 ;
        RECT 70.705 167.130 71.665 167.135 ;
        RECT 70.705 167.125 71.040 167.130 ;
        RECT 70.690 167.120 71.040 167.125 ;
        RECT 70.675 167.110 71.040 167.120 ;
        RECT 70.650 167.105 71.040 167.110 ;
        RECT 69.875 167.100 71.040 167.105 ;
        RECT 69.875 167.065 71.010 167.100 ;
        RECT 69.875 167.040 70.975 167.065 ;
        RECT 69.875 167.010 70.945 167.040 ;
        RECT 69.875 166.980 70.925 167.010 ;
        RECT 69.875 166.950 70.905 166.980 ;
        RECT 69.875 166.940 70.835 166.950 ;
        RECT 69.875 166.930 70.810 166.940 ;
        RECT 69.875 166.915 70.790 166.930 ;
        RECT 69.875 166.900 70.770 166.915 ;
        RECT 69.980 166.890 70.765 166.900 ;
        RECT 69.980 166.855 70.750 166.890 ;
        RECT 69.535 166.025 69.810 166.725 ;
        RECT 69.980 166.605 70.735 166.855 ;
        RECT 70.905 166.535 71.235 166.780 ;
        RECT 71.405 166.680 71.665 167.130 ;
        RECT 71.050 166.510 71.235 166.535 ;
        RECT 71.835 166.615 72.175 167.425 ;
        RECT 72.345 166.860 73.095 167.050 ;
        RECT 71.050 166.410 71.665 166.510 ;
        RECT 69.980 165.855 70.235 166.400 ;
        RECT 70.405 166.025 70.885 166.365 ;
        RECT 71.060 165.855 71.665 166.410 ;
        RECT 71.835 166.205 72.350 166.615 ;
        RECT 72.585 165.855 72.755 166.615 ;
        RECT 72.925 166.195 73.095 166.860 ;
        RECT 73.265 166.875 73.455 168.235 ;
        RECT 73.625 167.385 73.900 168.235 ;
        RECT 74.090 167.870 74.620 168.235 ;
        RECT 75.045 168.005 75.375 168.405 ;
        RECT 74.445 167.835 74.620 167.870 ;
        RECT 73.625 167.215 73.905 167.385 ;
        RECT 73.625 167.075 73.900 167.215 ;
        RECT 74.105 166.875 74.275 167.675 ;
        RECT 73.265 166.705 74.275 166.875 ;
        RECT 74.445 167.665 75.375 167.835 ;
        RECT 75.545 167.665 75.800 168.235 ;
        RECT 74.445 166.535 74.615 167.665 ;
        RECT 75.205 167.495 75.375 167.665 ;
        RECT 73.490 166.365 74.615 166.535 ;
        RECT 74.785 167.165 74.980 167.495 ;
        RECT 75.205 167.165 75.460 167.495 ;
        RECT 74.785 166.195 74.955 167.165 ;
        RECT 75.630 166.995 75.800 167.665 ;
        RECT 75.975 167.570 76.265 168.405 ;
        RECT 76.435 168.005 77.390 168.175 ;
        RECT 77.805 168.015 78.135 168.405 ;
        RECT 76.435 167.125 76.605 168.005 ;
        RECT 78.305 167.835 78.475 168.155 ;
        RECT 78.645 168.015 78.975 168.405 ;
        RECT 76.775 167.665 79.025 167.835 ;
        RECT 80.115 167.680 80.405 168.405 ;
        RECT 76.775 167.165 77.005 167.665 ;
        RECT 77.175 167.245 77.550 167.415 ;
        RECT 72.925 166.025 74.955 166.195 ;
        RECT 75.125 165.855 75.295 166.995 ;
        RECT 75.465 166.025 75.800 166.995 ;
        RECT 75.975 166.955 76.605 167.125 ;
        RECT 77.380 167.045 77.550 167.245 ;
        RECT 77.720 167.215 78.270 167.415 ;
        RECT 78.440 167.045 78.685 167.495 ;
        RECT 75.975 166.025 76.295 166.955 ;
        RECT 77.380 166.875 78.685 167.045 ;
        RECT 78.855 166.705 79.025 167.665 ;
        RECT 80.575 167.585 81.260 168.225 ;
        RECT 81.430 167.585 81.600 168.405 ;
        RECT 81.770 167.755 82.100 168.220 ;
        RECT 82.270 167.935 82.440 168.405 ;
        RECT 82.700 168.015 83.885 168.185 ;
        RECT 84.055 167.845 84.385 168.235 ;
        RECT 84.880 167.895 85.120 168.405 ;
        RECT 85.300 167.895 85.580 168.225 ;
        RECT 85.810 167.895 86.025 168.405 ;
        RECT 83.085 167.755 83.470 167.845 ;
        RECT 81.770 167.585 83.470 167.755 ;
        RECT 83.875 167.665 84.385 167.845 ;
        RECT 76.475 166.535 77.715 166.705 ;
        RECT 76.475 166.025 76.875 166.535 ;
        RECT 77.045 165.855 77.215 166.365 ;
        RECT 77.385 166.025 77.715 166.535 ;
        RECT 77.885 165.855 78.055 166.705 ;
        RECT 78.645 166.025 79.025 166.705 ;
        RECT 80.115 165.855 80.405 167.020 ;
        RECT 80.575 166.615 80.825 167.585 ;
        RECT 80.995 167.205 81.330 167.415 ;
        RECT 81.500 167.205 81.950 167.415 ;
        RECT 82.140 167.385 82.625 167.415 ;
        RECT 82.140 167.215 82.645 167.385 ;
        RECT 82.140 167.205 82.625 167.215 ;
        RECT 81.160 167.035 81.330 167.205 ;
        RECT 81.160 166.865 82.080 167.035 ;
        RECT 80.575 166.025 81.240 166.615 ;
        RECT 81.410 165.855 81.740 166.695 ;
        RECT 81.910 166.615 82.080 166.865 ;
        RECT 82.250 166.785 82.625 167.205 ;
        RECT 82.815 167.165 83.195 167.415 ;
        RECT 83.375 167.205 83.705 167.415 ;
        RECT 82.815 166.785 83.135 167.165 ;
        RECT 83.875 167.035 84.045 167.665 ;
        RECT 84.215 167.205 84.545 167.495 ;
        RECT 84.775 167.165 85.130 167.725 ;
        RECT 83.305 166.865 84.390 167.035 ;
        RECT 85.300 166.995 85.470 167.895 ;
        RECT 85.640 167.165 85.905 167.725 ;
        RECT 86.195 167.665 86.810 168.235 ;
        RECT 88.265 168.005 88.595 168.405 ;
        RECT 88.765 167.835 89.095 168.175 ;
        RECT 90.145 168.005 90.475 168.405 ;
        RECT 86.155 166.995 86.325 167.495 ;
        RECT 83.305 166.615 83.475 166.865 ;
        RECT 81.910 166.445 83.475 166.615 ;
        RECT 82.250 166.025 83.055 166.445 ;
        RECT 83.645 165.855 83.895 166.695 ;
        RECT 84.090 166.025 84.390 166.865 ;
        RECT 84.900 166.825 86.325 166.995 ;
        RECT 84.900 166.650 85.290 166.825 ;
        RECT 85.775 165.855 86.105 166.655 ;
        RECT 86.495 166.645 86.810 167.665 ;
        RECT 86.275 166.025 86.810 166.645 ;
        RECT 88.110 167.665 90.475 167.835 ;
        RECT 90.645 167.680 90.975 168.190 ;
        RECT 88.110 166.665 88.280 167.665 ;
        RECT 90.305 167.495 90.475 167.665 ;
        RECT 88.450 166.835 88.695 167.495 ;
        RECT 88.910 166.835 89.175 167.495 ;
        RECT 89.370 166.835 89.655 167.495 ;
        RECT 89.830 167.165 90.135 167.495 ;
        RECT 90.305 167.165 90.615 167.495 ;
        RECT 89.830 166.835 90.045 167.165 ;
        RECT 88.110 166.495 88.565 166.665 ;
        RECT 88.235 166.065 88.565 166.495 ;
        RECT 88.745 166.495 90.035 166.665 ;
        RECT 88.745 166.075 88.995 166.495 ;
        RECT 89.225 165.855 89.555 166.325 ;
        RECT 89.785 166.075 90.035 166.495 ;
        RECT 90.225 165.855 90.475 166.995 ;
        RECT 90.785 166.915 90.975 167.680 ;
        RECT 90.645 166.065 90.975 166.915 ;
        RECT 91.165 167.680 91.495 168.190 ;
        RECT 91.665 168.005 91.995 168.405 ;
        RECT 93.045 167.835 93.375 168.175 ;
        RECT 93.545 168.005 93.875 168.405 ;
        RECT 91.165 166.915 91.355 167.680 ;
        RECT 91.665 167.665 94.030 167.835 ;
        RECT 91.665 167.495 91.835 167.665 ;
        RECT 91.525 167.165 91.835 167.495 ;
        RECT 92.005 167.165 92.310 167.495 ;
        RECT 91.165 166.065 91.495 166.915 ;
        RECT 91.665 165.855 91.915 166.995 ;
        RECT 92.095 166.835 92.310 167.165 ;
        RECT 92.485 166.835 92.770 167.495 ;
        RECT 92.965 166.835 93.230 167.495 ;
        RECT 93.445 166.835 93.690 167.495 ;
        RECT 93.860 166.665 94.030 167.665 ;
        RECT 92.105 166.495 93.395 166.665 ;
        RECT 92.105 166.075 92.355 166.495 ;
        RECT 92.585 165.855 92.915 166.325 ;
        RECT 93.145 166.075 93.395 166.495 ;
        RECT 93.575 166.495 94.030 166.665 ;
        RECT 94.835 167.665 95.220 168.235 ;
        RECT 95.390 167.945 95.715 168.405 ;
        RECT 96.235 167.775 96.515 168.235 ;
        RECT 94.835 166.995 95.115 167.665 ;
        RECT 95.390 167.605 96.515 167.775 ;
        RECT 95.390 167.495 95.840 167.605 ;
        RECT 95.285 167.165 95.840 167.495 ;
        RECT 96.705 167.435 97.105 168.235 ;
        RECT 97.505 167.945 97.775 168.405 ;
        RECT 97.945 167.775 98.230 168.235 ;
        RECT 93.575 166.065 93.905 166.495 ;
        RECT 94.835 166.025 95.220 166.995 ;
        RECT 95.390 166.705 95.840 167.165 ;
        RECT 96.010 166.875 97.105 167.435 ;
        RECT 95.390 166.485 96.515 166.705 ;
        RECT 95.390 165.855 95.715 166.315 ;
        RECT 96.235 166.025 96.515 166.485 ;
        RECT 96.705 166.025 97.105 166.875 ;
        RECT 97.275 167.605 98.230 167.775 ;
        RECT 98.550 167.665 99.165 168.235 ;
        RECT 99.335 167.895 99.550 168.405 ;
        RECT 99.780 167.895 100.060 168.225 ;
        RECT 100.240 167.895 100.480 168.405 ;
        RECT 97.275 166.705 97.485 167.605 ;
        RECT 97.655 166.875 98.345 167.435 ;
        RECT 97.275 166.485 98.230 166.705 ;
        RECT 97.505 165.855 97.775 166.315 ;
        RECT 97.945 166.025 98.230 166.485 ;
        RECT 98.550 166.645 98.865 167.665 ;
        RECT 99.035 166.995 99.205 167.495 ;
        RECT 99.455 167.165 99.720 167.725 ;
        RECT 99.890 166.995 100.060 167.895 ;
        RECT 100.230 167.165 100.585 167.725 ;
        RECT 101.735 167.605 102.075 168.235 ;
        RECT 102.365 167.945 102.535 168.405 ;
        RECT 102.805 167.775 103.135 168.220 ;
        RECT 101.735 167.035 102.005 167.605 ;
        RECT 102.385 167.585 103.135 167.775 ;
        RECT 103.305 167.755 103.475 168.075 ;
        RECT 103.700 167.945 104.030 168.405 ;
        RECT 104.230 167.755 104.560 168.235 ;
        RECT 104.775 167.945 105.105 168.405 ;
        RECT 105.275 167.755 105.605 168.235 ;
        RECT 103.305 167.585 105.605 167.755 ;
        RECT 105.875 167.680 106.165 168.405 ;
        RECT 106.395 167.585 106.605 168.405 ;
        RECT 106.775 167.605 107.105 168.235 ;
        RECT 102.385 167.415 102.755 167.585 ;
        RECT 102.175 167.205 102.755 167.415 ;
        RECT 102.925 167.205 103.345 167.415 ;
        RECT 102.495 167.035 102.755 167.205 ;
        RECT 99.035 166.825 100.460 166.995 ;
        RECT 98.550 166.025 99.085 166.645 ;
        RECT 99.255 165.855 99.585 166.655 ;
        RECT 100.070 166.650 100.460 166.825 ;
        RECT 101.735 166.025 102.260 167.035 ;
        RECT 102.495 166.745 103.245 167.035 ;
        RECT 102.495 165.855 102.825 166.575 ;
        RECT 102.995 166.025 103.245 166.745 ;
        RECT 103.515 166.100 103.845 167.415 ;
        RECT 104.055 166.100 104.385 167.415 ;
        RECT 104.555 166.100 104.925 167.415 ;
        RECT 105.135 167.165 105.645 167.415 ;
        RECT 105.255 165.855 105.585 166.975 ;
        RECT 105.875 165.855 106.165 167.020 ;
        RECT 106.775 167.005 107.025 167.605 ;
        RECT 107.275 167.585 107.505 168.405 ;
        RECT 107.715 167.895 108.020 168.405 ;
        RECT 107.195 167.165 107.525 167.415 ;
        RECT 107.715 167.165 108.030 167.725 ;
        RECT 108.200 167.415 108.450 168.225 ;
        RECT 108.620 167.880 108.880 168.405 ;
        RECT 109.060 167.415 109.310 168.225 ;
        RECT 109.480 167.845 109.740 168.405 ;
        RECT 109.910 167.755 110.170 168.210 ;
        RECT 110.340 167.925 110.600 168.405 ;
        RECT 110.770 167.755 111.030 168.210 ;
        RECT 111.200 167.925 111.460 168.405 ;
        RECT 111.630 167.755 111.890 168.210 ;
        RECT 112.060 167.925 112.305 168.405 ;
        RECT 112.475 167.755 112.750 168.210 ;
        RECT 112.920 167.925 113.165 168.405 ;
        RECT 113.335 167.755 113.595 168.210 ;
        RECT 113.775 167.925 114.025 168.405 ;
        RECT 114.195 167.755 114.455 168.210 ;
        RECT 114.635 167.925 114.885 168.405 ;
        RECT 115.055 167.755 115.315 168.210 ;
        RECT 115.495 167.925 115.755 168.405 ;
        RECT 115.925 167.755 116.185 168.210 ;
        RECT 116.355 167.925 116.655 168.405 ;
        RECT 117.225 167.935 117.395 168.405 ;
        RECT 117.565 167.755 117.895 168.235 ;
        RECT 118.065 167.935 118.235 168.405 ;
        RECT 118.405 167.755 118.735 168.235 ;
        RECT 109.910 167.585 116.655 167.755 ;
        RECT 108.200 167.165 115.320 167.415 ;
        RECT 106.395 165.855 106.605 166.995 ;
        RECT 106.775 166.025 107.105 167.005 ;
        RECT 107.275 165.855 107.505 166.995 ;
        RECT 107.725 165.855 108.020 166.665 ;
        RECT 108.200 166.025 108.445 167.165 ;
        RECT 108.620 165.855 108.880 166.665 ;
        RECT 109.060 166.030 109.310 167.165 ;
        RECT 115.490 166.995 116.655 167.585 ;
        RECT 109.910 166.770 116.655 166.995 ;
        RECT 116.970 167.585 118.735 167.755 ;
        RECT 118.905 167.595 119.075 168.405 ;
        RECT 119.275 168.025 120.345 168.195 ;
        RECT 119.275 167.670 119.595 168.025 ;
        RECT 116.970 167.035 117.380 167.585 ;
        RECT 119.270 167.415 119.595 167.670 ;
        RECT 117.565 167.205 119.595 167.415 ;
        RECT 119.250 167.195 119.595 167.205 ;
        RECT 119.765 167.455 120.005 167.855 ;
        RECT 120.175 167.795 120.345 168.025 ;
        RECT 120.515 167.965 120.705 168.405 ;
        RECT 120.875 167.955 121.825 168.235 ;
        RECT 122.045 168.045 122.395 168.215 ;
        RECT 120.175 167.625 120.705 167.795 ;
        RECT 116.970 166.865 118.695 167.035 ;
        RECT 109.910 166.755 115.315 166.770 ;
        RECT 109.480 165.860 109.740 166.655 ;
        RECT 109.910 166.030 110.170 166.755 ;
        RECT 110.340 165.860 110.600 166.585 ;
        RECT 110.770 166.030 111.030 166.755 ;
        RECT 111.200 165.860 111.460 166.585 ;
        RECT 111.630 166.030 111.890 166.755 ;
        RECT 112.060 165.860 112.320 166.585 ;
        RECT 112.490 166.030 112.750 166.755 ;
        RECT 112.920 165.860 113.165 166.585 ;
        RECT 113.335 166.030 113.595 166.755 ;
        RECT 113.780 165.860 114.025 166.585 ;
        RECT 114.195 166.030 114.455 166.755 ;
        RECT 114.640 165.860 114.885 166.585 ;
        RECT 115.055 166.030 115.315 166.755 ;
        RECT 115.500 165.860 115.755 166.585 ;
        RECT 115.925 166.030 116.215 166.770 ;
        RECT 109.480 165.855 115.755 165.860 ;
        RECT 116.385 165.855 116.655 166.600 ;
        RECT 117.225 165.855 117.395 166.695 ;
        RECT 117.605 166.025 117.855 166.865 ;
        RECT 118.065 165.855 118.235 166.695 ;
        RECT 118.405 166.025 118.695 166.865 ;
        RECT 118.905 165.855 119.075 166.915 ;
        RECT 119.250 166.575 119.420 167.195 ;
        RECT 119.765 167.085 120.305 167.455 ;
        RECT 120.485 167.345 120.705 167.625 ;
        RECT 120.875 167.175 121.045 167.955 ;
        RECT 120.640 167.005 121.045 167.175 ;
        RECT 121.215 167.165 121.565 167.785 ;
        RECT 120.640 166.915 120.810 167.005 ;
        RECT 121.735 166.995 121.945 167.785 ;
        RECT 119.590 166.745 120.810 166.915 ;
        RECT 121.270 166.835 121.945 166.995 ;
        RECT 119.250 166.405 120.050 166.575 ;
        RECT 119.370 165.855 119.700 166.235 ;
        RECT 119.880 166.115 120.050 166.405 ;
        RECT 120.640 166.365 120.810 166.745 ;
        RECT 120.980 166.825 121.945 166.835 ;
        RECT 122.135 167.655 122.395 168.045 ;
        RECT 122.605 167.945 122.935 168.405 ;
        RECT 123.810 168.015 124.665 168.185 ;
        RECT 124.870 168.015 125.365 168.185 ;
        RECT 125.535 168.045 125.865 168.405 ;
        RECT 122.135 166.965 122.305 167.655 ;
        RECT 122.475 167.305 122.645 167.485 ;
        RECT 122.815 167.475 123.605 167.725 ;
        RECT 123.810 167.305 123.980 168.015 ;
        RECT 124.150 167.505 124.505 167.725 ;
        RECT 122.475 167.135 124.165 167.305 ;
        RECT 120.980 166.535 121.440 166.825 ;
        RECT 122.135 166.795 123.635 166.965 ;
        RECT 122.135 166.655 122.305 166.795 ;
        RECT 121.745 166.485 122.305 166.655 ;
        RECT 120.220 165.855 120.470 166.315 ;
        RECT 120.640 166.025 121.510 166.365 ;
        RECT 121.745 166.025 121.915 166.485 ;
        RECT 122.750 166.455 123.825 166.625 ;
        RECT 122.085 165.855 122.455 166.315 ;
        RECT 122.750 166.115 122.920 166.455 ;
        RECT 123.090 165.855 123.420 166.285 ;
        RECT 123.655 166.115 123.825 166.455 ;
        RECT 123.995 166.355 124.165 167.135 ;
        RECT 124.335 166.915 124.505 167.505 ;
        RECT 124.675 167.105 125.025 167.725 ;
        RECT 124.335 166.525 124.800 166.915 ;
        RECT 125.195 166.655 125.365 168.015 ;
        RECT 125.535 166.825 125.995 167.875 ;
        RECT 124.970 166.485 125.365 166.655 ;
        RECT 124.970 166.355 125.140 166.485 ;
        RECT 123.995 166.025 124.675 166.355 ;
        RECT 124.890 166.025 125.140 166.355 ;
        RECT 125.310 165.855 125.560 166.315 ;
        RECT 125.730 166.040 126.055 166.825 ;
        RECT 126.225 166.025 126.395 168.145 ;
        RECT 126.565 168.025 126.895 168.405 ;
        RECT 127.065 167.855 127.320 168.145 ;
        RECT 126.570 167.685 127.320 167.855 ;
        RECT 126.570 166.695 126.800 167.685 ;
        RECT 127.495 167.635 131.005 168.405 ;
        RECT 131.635 167.680 131.925 168.405 ;
        RECT 133.230 167.935 133.515 168.405 ;
        RECT 133.685 167.765 134.015 168.235 ;
        RECT 134.185 167.935 134.355 168.405 ;
        RECT 134.525 167.765 134.855 168.235 ;
        RECT 135.025 167.935 135.195 168.405 ;
        RECT 135.365 167.765 135.695 168.235 ;
        RECT 135.865 167.935 136.035 168.405 ;
        RECT 136.205 167.765 136.535 168.235 ;
        RECT 126.970 166.865 127.320 167.515 ;
        RECT 127.495 167.115 129.145 167.635 ;
        RECT 133.015 167.585 136.535 167.765 ;
        RECT 136.705 167.585 136.980 168.405 ;
        RECT 137.245 167.755 137.415 168.235 ;
        RECT 137.595 167.925 137.835 168.405 ;
        RECT 138.085 167.755 138.255 168.235 ;
        RECT 138.425 167.925 138.755 168.405 ;
        RECT 138.925 167.755 139.095 168.235 ;
        RECT 137.245 167.585 137.880 167.755 ;
        RECT 138.085 167.585 139.095 167.755 ;
        RECT 139.265 167.605 139.595 168.405 ;
        RECT 140.065 167.605 140.395 168.405 ;
        RECT 140.565 167.755 140.735 168.235 ;
        RECT 140.905 167.925 141.235 168.405 ;
        RECT 141.405 167.755 141.575 168.235 ;
        RECT 141.825 167.925 142.065 168.405 ;
        RECT 142.245 167.755 142.415 168.235 ;
        RECT 129.315 166.945 131.005 167.465 ;
        RECT 133.015 167.045 133.415 167.585 ;
        RECT 137.710 167.415 137.880 167.585 ;
        RECT 133.585 167.215 134.950 167.415 ;
        RECT 135.270 167.215 136.930 167.415 ;
        RECT 137.160 167.175 137.540 167.415 ;
        RECT 137.710 167.245 138.210 167.415 ;
        RECT 126.570 166.525 127.320 166.695 ;
        RECT 126.565 165.855 126.895 166.355 ;
        RECT 127.065 166.025 127.320 166.525 ;
        RECT 127.495 165.855 131.005 166.945 ;
        RECT 131.635 165.855 131.925 167.020 ;
        RECT 133.015 166.745 134.775 167.045 ;
        RECT 133.180 166.195 133.595 166.575 ;
        RECT 133.765 166.365 133.935 166.745 ;
        RECT 134.105 166.195 134.435 166.555 ;
        RECT 134.605 166.365 134.775 166.745 ;
        RECT 134.945 166.825 136.980 167.035 ;
        RECT 137.710 167.005 137.880 167.245 ;
        RECT 138.600 167.045 139.095 167.585 ;
        RECT 134.945 166.195 135.275 166.825 ;
        RECT 133.180 166.025 135.275 166.195 ;
        RECT 135.445 165.855 135.695 166.655 ;
        RECT 135.865 166.025 136.035 166.825 ;
        RECT 136.205 165.855 136.535 166.655 ;
        RECT 136.705 166.025 136.980 166.825 ;
        RECT 137.165 166.835 137.880 167.005 ;
        RECT 138.085 166.875 139.095 167.045 ;
        RECT 140.565 167.585 141.575 167.755 ;
        RECT 141.780 167.585 142.415 167.755 ;
        RECT 142.675 167.635 144.345 168.405 ;
        RECT 144.630 167.775 144.915 168.235 ;
        RECT 145.085 167.945 145.355 168.405 ;
        RECT 140.565 167.045 141.060 167.585 ;
        RECT 141.780 167.415 141.950 167.585 ;
        RECT 141.450 167.245 141.950 167.415 ;
        RECT 137.165 166.025 137.495 166.835 ;
        RECT 137.665 165.855 137.905 166.655 ;
        RECT 138.085 166.025 138.255 166.875 ;
        RECT 138.425 165.855 138.755 166.655 ;
        RECT 138.925 166.025 139.095 166.875 ;
        RECT 139.265 165.855 139.595 167.005 ;
        RECT 140.065 165.855 140.395 167.005 ;
        RECT 140.565 166.875 141.575 167.045 ;
        RECT 140.565 166.025 140.735 166.875 ;
        RECT 140.905 165.855 141.235 166.655 ;
        RECT 141.405 166.025 141.575 166.875 ;
        RECT 141.780 167.005 141.950 167.245 ;
        RECT 142.120 167.175 142.500 167.415 ;
        RECT 142.675 167.115 143.425 167.635 ;
        RECT 144.630 167.605 145.585 167.775 ;
        RECT 141.780 166.835 142.495 167.005 ;
        RECT 143.595 166.945 144.345 167.465 ;
        RECT 141.755 165.855 141.995 166.655 ;
        RECT 142.165 166.025 142.495 166.835 ;
        RECT 142.675 165.855 144.345 166.945 ;
        RECT 144.515 166.875 145.205 167.435 ;
        RECT 145.375 166.705 145.585 167.605 ;
        RECT 144.630 166.485 145.585 166.705 ;
        RECT 145.755 167.435 146.155 168.235 ;
        RECT 146.345 167.775 146.625 168.235 ;
        RECT 147.145 167.945 147.470 168.405 ;
        RECT 146.345 167.605 147.470 167.775 ;
        RECT 147.640 167.665 148.025 168.235 ;
        RECT 147.020 167.495 147.470 167.605 ;
        RECT 145.755 166.875 146.850 167.435 ;
        RECT 147.020 167.165 147.575 167.495 ;
        RECT 144.630 166.025 144.915 166.485 ;
        RECT 145.085 165.855 145.355 166.315 ;
        RECT 145.755 166.025 146.155 166.875 ;
        RECT 147.020 166.705 147.470 167.165 ;
        RECT 147.745 166.995 148.025 167.665 ;
        RECT 148.200 167.565 148.460 168.405 ;
        RECT 148.635 167.660 148.890 168.235 ;
        RECT 149.060 168.025 149.390 168.405 ;
        RECT 149.605 167.855 149.775 168.235 ;
        RECT 149.060 167.685 149.775 167.855 ;
        RECT 150.125 167.855 150.295 168.235 ;
        RECT 150.510 168.025 150.840 168.405 ;
        RECT 150.125 167.685 150.840 167.855 ;
        RECT 146.345 166.485 147.470 166.705 ;
        RECT 146.345 166.025 146.625 166.485 ;
        RECT 147.145 165.855 147.470 166.315 ;
        RECT 147.640 166.025 148.025 166.995 ;
        RECT 148.200 165.855 148.460 167.005 ;
        RECT 148.635 166.930 148.805 167.660 ;
        RECT 149.060 167.495 149.230 167.685 ;
        RECT 148.975 167.165 149.230 167.495 ;
        RECT 149.060 166.955 149.230 167.165 ;
        RECT 149.510 167.135 149.865 167.505 ;
        RECT 150.035 167.135 150.390 167.505 ;
        RECT 150.670 167.495 150.840 167.685 ;
        RECT 151.010 167.660 151.265 168.235 ;
        RECT 150.670 167.165 150.925 167.495 ;
        RECT 150.670 166.955 150.840 167.165 ;
        RECT 148.635 166.025 148.890 166.930 ;
        RECT 149.060 166.785 149.775 166.955 ;
        RECT 149.060 165.855 149.390 166.615 ;
        RECT 149.605 166.025 149.775 166.785 ;
        RECT 150.125 166.785 150.840 166.955 ;
        RECT 151.095 166.930 151.265 167.660 ;
        RECT 151.440 167.565 151.700 168.405 ;
        RECT 151.875 167.635 155.385 168.405 ;
        RECT 155.555 167.655 156.765 168.405 ;
        RECT 156.935 167.655 158.145 168.405 ;
        RECT 151.875 167.115 153.525 167.635 ;
        RECT 150.125 166.025 150.295 166.785 ;
        RECT 150.510 165.855 150.840 166.615 ;
        RECT 151.010 166.025 151.265 166.930 ;
        RECT 151.440 165.855 151.700 167.005 ;
        RECT 153.695 166.945 155.385 167.465 ;
        RECT 155.555 167.115 156.075 167.655 ;
        RECT 156.245 166.945 156.765 167.485 ;
        RECT 151.875 165.855 155.385 166.945 ;
        RECT 155.555 165.855 156.765 166.945 ;
        RECT 156.935 166.945 157.455 167.485 ;
        RECT 157.625 167.115 158.145 167.655 ;
        RECT 156.935 165.855 158.145 166.945 ;
        RECT 2.750 165.685 158.230 165.855 ;
        RECT 2.835 164.595 4.045 165.685 ;
        RECT 4.305 165.015 4.475 165.515 ;
        RECT 4.645 165.185 4.975 165.685 ;
        RECT 4.305 164.845 4.970 165.015 ;
        RECT 2.835 163.885 3.355 164.425 ;
        RECT 3.525 164.055 4.045 164.595 ;
        RECT 4.220 164.025 4.570 164.675 ;
        RECT 2.835 163.135 4.045 163.885 ;
        RECT 4.740 163.855 4.970 164.845 ;
        RECT 4.305 163.685 4.970 163.855 ;
        RECT 4.305 163.395 4.475 163.685 ;
        RECT 4.645 163.135 4.975 163.515 ;
        RECT 5.145 163.395 5.370 165.515 ;
        RECT 5.585 165.185 5.915 165.685 ;
        RECT 6.085 165.015 6.255 165.515 ;
        RECT 6.490 165.300 7.320 165.470 ;
        RECT 7.560 165.305 7.940 165.685 ;
        RECT 5.560 164.845 6.255 165.015 ;
        RECT 5.560 163.875 5.730 164.845 ;
        RECT 5.900 164.055 6.310 164.675 ;
        RECT 6.480 164.625 6.980 165.005 ;
        RECT 5.560 163.685 6.255 163.875 ;
        RECT 6.480 163.755 6.700 164.625 ;
        RECT 7.150 164.455 7.320 165.300 ;
        RECT 8.120 165.135 8.290 165.425 ;
        RECT 8.460 165.305 8.790 165.685 ;
        RECT 9.260 165.215 9.890 165.465 ;
        RECT 10.070 165.305 10.490 165.685 ;
        RECT 9.720 165.135 9.890 165.215 ;
        RECT 10.690 165.135 10.930 165.425 ;
        RECT 7.490 164.885 8.860 165.135 ;
        RECT 7.490 164.625 7.740 164.885 ;
        RECT 8.250 164.455 8.500 164.615 ;
        RECT 7.150 164.285 8.500 164.455 ;
        RECT 7.150 164.245 7.570 164.285 ;
        RECT 6.880 163.695 7.230 164.065 ;
        RECT 5.585 163.135 5.915 163.515 ;
        RECT 6.085 163.355 6.255 163.685 ;
        RECT 7.400 163.515 7.570 164.245 ;
        RECT 8.670 164.115 8.860 164.885 ;
        RECT 7.740 163.785 8.150 164.115 ;
        RECT 8.440 163.775 8.860 164.115 ;
        RECT 9.030 164.705 9.550 165.015 ;
        RECT 9.720 164.965 10.930 165.135 ;
        RECT 11.160 164.995 11.490 165.685 ;
        RECT 9.030 163.945 9.200 164.705 ;
        RECT 9.370 164.115 9.550 164.525 ;
        RECT 9.720 164.455 9.890 164.965 ;
        RECT 11.660 164.815 11.830 165.425 ;
        RECT 12.100 164.965 12.430 165.475 ;
        RECT 11.660 164.795 11.980 164.815 ;
        RECT 10.060 164.625 11.980 164.795 ;
        RECT 9.720 164.285 11.620 164.455 ;
        RECT 9.950 163.945 10.280 164.065 ;
        RECT 9.030 163.775 10.280 163.945 ;
        RECT 6.555 163.315 7.570 163.515 ;
        RECT 7.740 163.135 8.150 163.575 ;
        RECT 8.440 163.345 8.690 163.775 ;
        RECT 8.890 163.135 9.210 163.595 ;
        RECT 10.450 163.525 10.620 164.285 ;
        RECT 11.290 164.225 11.620 164.285 ;
        RECT 10.810 164.055 11.140 164.115 ;
        RECT 10.810 163.785 11.470 164.055 ;
        RECT 11.790 163.730 11.980 164.625 ;
        RECT 9.770 163.355 10.620 163.525 ;
        RECT 10.820 163.135 11.480 163.615 ;
        RECT 11.660 163.400 11.980 163.730 ;
        RECT 12.180 164.375 12.430 164.965 ;
        RECT 12.610 164.885 12.895 165.685 ;
        RECT 13.075 165.345 13.330 165.375 ;
        RECT 13.075 165.175 13.415 165.345 ;
        RECT 13.075 164.705 13.330 165.175 ;
        RECT 12.180 164.045 12.980 164.375 ;
        RECT 12.180 163.395 12.430 164.045 ;
        RECT 13.150 163.845 13.330 164.705 ;
        RECT 12.610 163.135 12.895 163.595 ;
        RECT 13.075 163.315 13.330 163.845 ;
        RECT 13.875 164.610 14.145 165.515 ;
        RECT 14.315 164.925 14.645 165.685 ;
        RECT 14.825 164.755 14.995 165.515 ;
        RECT 13.875 163.810 14.045 164.610 ;
        RECT 14.330 164.585 14.995 164.755 ;
        RECT 14.330 164.440 14.500 164.585 ;
        RECT 15.715 164.520 16.005 165.685 ;
        RECT 16.180 164.545 16.515 165.515 ;
        RECT 16.685 164.545 16.855 165.685 ;
        RECT 17.025 165.345 19.055 165.515 ;
        RECT 14.215 164.110 14.500 164.440 ;
        RECT 14.330 163.855 14.500 164.110 ;
        RECT 14.735 164.035 15.065 164.405 ;
        RECT 16.180 163.875 16.350 164.545 ;
        RECT 17.025 164.375 17.195 165.345 ;
        RECT 16.520 164.045 16.775 164.375 ;
        RECT 17.000 164.045 17.195 164.375 ;
        RECT 17.365 165.005 18.490 165.175 ;
        RECT 16.605 163.875 16.775 164.045 ;
        RECT 17.365 163.875 17.535 165.005 ;
        RECT 13.875 163.305 14.135 163.810 ;
        RECT 14.330 163.685 14.995 163.855 ;
        RECT 14.315 163.135 14.645 163.515 ;
        RECT 14.825 163.305 14.995 163.685 ;
        RECT 15.715 163.135 16.005 163.860 ;
        RECT 16.180 163.305 16.435 163.875 ;
        RECT 16.605 163.705 17.535 163.875 ;
        RECT 17.705 164.665 18.715 164.835 ;
        RECT 17.705 163.865 17.875 164.665 ;
        RECT 18.080 163.985 18.355 164.465 ;
        RECT 18.075 163.815 18.355 163.985 ;
        RECT 17.360 163.670 17.535 163.705 ;
        RECT 16.605 163.135 16.935 163.535 ;
        RECT 17.360 163.305 17.890 163.670 ;
        RECT 18.080 163.305 18.355 163.815 ;
        RECT 18.525 163.305 18.715 164.665 ;
        RECT 18.885 164.680 19.055 165.345 ;
        RECT 19.225 164.925 19.395 165.685 ;
        RECT 19.630 164.925 20.145 165.335 ;
        RECT 18.885 164.490 19.635 164.680 ;
        RECT 19.805 164.115 20.145 164.925 ;
        RECT 20.315 164.595 21.985 165.685 ;
        RECT 18.915 163.945 20.145 164.115 ;
        RECT 18.895 163.135 19.405 163.670 ;
        RECT 19.625 163.340 19.870 163.945 ;
        RECT 20.315 163.905 21.065 164.425 ;
        RECT 21.235 164.075 21.985 164.595 ;
        RECT 22.245 164.675 22.415 165.515 ;
        RECT 22.585 165.345 23.755 165.515 ;
        RECT 22.585 164.845 22.915 165.345 ;
        RECT 23.425 165.305 23.755 165.345 ;
        RECT 23.945 165.265 24.300 165.685 ;
        RECT 23.085 165.085 23.315 165.175 ;
        RECT 24.470 165.085 24.720 165.515 ;
        RECT 23.085 164.845 24.720 165.085 ;
        RECT 24.890 164.925 25.220 165.685 ;
        RECT 25.390 164.845 25.645 165.515 ;
        RECT 22.245 164.505 25.305 164.675 ;
        RECT 22.160 164.125 22.510 164.335 ;
        RECT 22.680 164.125 23.125 164.325 ;
        RECT 23.295 164.125 23.770 164.325 ;
        RECT 20.315 163.135 21.985 163.905 ;
        RECT 22.245 163.785 23.310 163.955 ;
        RECT 22.245 163.305 22.415 163.785 ;
        RECT 22.585 163.135 22.915 163.615 ;
        RECT 23.140 163.555 23.310 163.785 ;
        RECT 23.490 163.725 23.770 164.125 ;
        RECT 24.040 164.125 24.370 164.325 ;
        RECT 24.540 164.125 24.905 164.325 ;
        RECT 24.040 163.725 24.325 164.125 ;
        RECT 25.135 163.955 25.305 164.505 ;
        RECT 24.505 163.785 25.305 163.955 ;
        RECT 24.505 163.555 24.675 163.785 ;
        RECT 25.475 163.715 25.645 164.845 ;
        RECT 26.845 164.755 27.015 165.515 ;
        RECT 27.195 164.925 27.525 165.685 ;
        RECT 26.845 164.585 27.510 164.755 ;
        RECT 27.695 164.610 27.965 165.515 ;
        RECT 27.340 164.440 27.510 164.585 ;
        RECT 26.775 164.035 27.105 164.405 ;
        RECT 27.340 164.110 27.625 164.440 ;
        RECT 27.340 163.855 27.510 164.110 ;
        RECT 25.460 163.645 25.645 163.715 ;
        RECT 25.435 163.635 25.645 163.645 ;
        RECT 23.140 163.305 24.675 163.555 ;
        RECT 24.845 163.135 25.175 163.615 ;
        RECT 25.390 163.305 25.645 163.635 ;
        RECT 26.845 163.685 27.510 163.855 ;
        RECT 27.795 163.810 27.965 164.610 ;
        RECT 26.845 163.305 27.015 163.685 ;
        RECT 27.195 163.135 27.525 163.515 ;
        RECT 27.705 163.305 27.965 163.810 ;
        RECT 28.140 164.545 28.475 165.515 ;
        RECT 28.645 164.545 28.815 165.685 ;
        RECT 28.985 165.345 31.015 165.515 ;
        RECT 28.140 163.875 28.310 164.545 ;
        RECT 28.985 164.375 29.155 165.345 ;
        RECT 28.480 164.045 28.735 164.375 ;
        RECT 28.960 164.045 29.155 164.375 ;
        RECT 29.325 165.005 30.450 165.175 ;
        RECT 28.565 163.875 28.735 164.045 ;
        RECT 29.325 163.875 29.495 165.005 ;
        RECT 28.140 163.305 28.395 163.875 ;
        RECT 28.565 163.705 29.495 163.875 ;
        RECT 29.665 164.665 30.675 164.835 ;
        RECT 29.665 163.865 29.835 164.665 ;
        RECT 30.040 164.325 30.315 164.465 ;
        RECT 30.035 164.155 30.315 164.325 ;
        RECT 29.320 163.670 29.495 163.705 ;
        RECT 28.565 163.135 28.895 163.535 ;
        RECT 29.320 163.305 29.850 163.670 ;
        RECT 30.040 163.305 30.315 164.155 ;
        RECT 30.485 163.305 30.675 164.665 ;
        RECT 30.845 164.680 31.015 165.345 ;
        RECT 31.185 164.925 31.355 165.685 ;
        RECT 31.590 164.925 32.105 165.335 ;
        RECT 32.365 164.940 32.635 165.685 ;
        RECT 33.265 165.680 39.540 165.685 ;
        RECT 30.845 164.490 31.595 164.680 ;
        RECT 31.765 164.115 32.105 164.925 ;
        RECT 32.805 164.770 33.095 165.510 ;
        RECT 33.265 164.955 33.520 165.680 ;
        RECT 33.705 164.785 33.965 165.510 ;
        RECT 34.135 164.955 34.380 165.680 ;
        RECT 34.565 164.785 34.825 165.510 ;
        RECT 34.995 164.955 35.240 165.680 ;
        RECT 35.425 164.785 35.685 165.510 ;
        RECT 35.855 164.955 36.100 165.680 ;
        RECT 36.270 164.785 36.530 165.510 ;
        RECT 36.700 164.955 36.960 165.680 ;
        RECT 37.130 164.785 37.390 165.510 ;
        RECT 37.560 164.955 37.820 165.680 ;
        RECT 37.990 164.785 38.250 165.510 ;
        RECT 38.420 164.955 38.680 165.680 ;
        RECT 38.850 164.785 39.110 165.510 ;
        RECT 39.280 164.885 39.540 165.680 ;
        RECT 33.705 164.770 39.110 164.785 ;
        RECT 30.875 163.945 32.105 164.115 ;
        RECT 32.365 164.545 39.110 164.770 ;
        RECT 32.365 163.955 33.530 164.545 ;
        RECT 39.710 164.375 39.960 165.510 ;
        RECT 40.140 164.875 40.400 165.685 ;
        RECT 40.575 164.375 40.820 165.515 ;
        RECT 41.000 164.875 41.295 165.685 ;
        RECT 41.475 164.520 41.765 165.685 ;
        RECT 42.025 164.675 42.195 165.515 ;
        RECT 42.365 165.345 43.535 165.515 ;
        RECT 42.365 164.845 42.695 165.345 ;
        RECT 43.205 165.305 43.535 165.345 ;
        RECT 43.725 165.265 44.080 165.685 ;
        RECT 42.865 165.085 43.095 165.175 ;
        RECT 44.250 165.085 44.500 165.515 ;
        RECT 42.865 164.845 44.500 165.085 ;
        RECT 44.670 164.925 45.000 165.685 ;
        RECT 45.170 164.845 45.425 165.515 ;
        RECT 42.025 164.505 45.085 164.675 ;
        RECT 33.700 164.125 40.820 164.375 ;
        RECT 30.855 163.135 31.365 163.670 ;
        RECT 31.585 163.340 31.830 163.945 ;
        RECT 32.365 163.785 39.110 163.955 ;
        RECT 32.365 163.135 32.665 163.615 ;
        RECT 32.835 163.330 33.095 163.785 ;
        RECT 33.265 163.135 33.525 163.615 ;
        RECT 33.705 163.330 33.965 163.785 ;
        RECT 34.135 163.135 34.385 163.615 ;
        RECT 34.565 163.330 34.825 163.785 ;
        RECT 34.995 163.135 35.245 163.615 ;
        RECT 35.425 163.330 35.685 163.785 ;
        RECT 35.855 163.135 36.100 163.615 ;
        RECT 36.270 163.330 36.545 163.785 ;
        RECT 36.715 163.135 36.960 163.615 ;
        RECT 37.130 163.330 37.390 163.785 ;
        RECT 37.560 163.135 37.820 163.615 ;
        RECT 37.990 163.330 38.250 163.785 ;
        RECT 38.420 163.135 38.680 163.615 ;
        RECT 38.850 163.330 39.110 163.785 ;
        RECT 39.280 163.135 39.540 163.695 ;
        RECT 39.710 163.315 39.960 164.125 ;
        RECT 40.140 163.135 40.400 163.660 ;
        RECT 40.570 163.315 40.820 164.125 ;
        RECT 40.990 163.815 41.305 164.375 ;
        RECT 41.940 164.125 42.290 164.335 ;
        RECT 42.460 164.125 42.905 164.325 ;
        RECT 43.075 164.125 43.550 164.325 ;
        RECT 41.000 163.135 41.305 163.645 ;
        RECT 41.475 163.135 41.765 163.860 ;
        RECT 42.025 163.785 43.090 163.955 ;
        RECT 42.025 163.305 42.195 163.785 ;
        RECT 42.365 163.135 42.695 163.615 ;
        RECT 42.920 163.555 43.090 163.785 ;
        RECT 43.270 163.725 43.550 164.125 ;
        RECT 43.820 164.125 44.150 164.325 ;
        RECT 44.320 164.155 44.695 164.325 ;
        RECT 44.320 164.125 44.685 164.155 ;
        RECT 43.820 163.725 44.105 164.125 ;
        RECT 44.915 163.955 45.085 164.505 ;
        RECT 44.285 163.785 45.085 163.955 ;
        RECT 44.285 163.555 44.455 163.785 ;
        RECT 45.255 163.715 45.425 164.845 ;
        RECT 46.130 164.815 46.415 165.685 ;
        RECT 46.585 165.055 46.845 165.515 ;
        RECT 47.020 165.225 47.275 165.685 ;
        RECT 47.445 165.055 47.705 165.515 ;
        RECT 46.585 164.885 47.705 165.055 ;
        RECT 47.875 164.885 48.185 165.685 ;
        RECT 46.585 164.635 46.845 164.885 ;
        RECT 47.055 164.835 47.225 164.885 ;
        RECT 48.355 164.715 48.665 165.515 ;
        RECT 46.090 164.465 46.845 164.635 ;
        RECT 47.635 164.545 48.665 164.715 ;
        RECT 46.090 163.955 46.495 164.465 ;
        RECT 47.635 164.295 47.805 164.545 ;
        RECT 46.665 164.125 47.805 164.295 ;
        RECT 46.090 163.785 47.740 163.955 ;
        RECT 47.975 163.805 48.325 164.375 ;
        RECT 45.240 163.645 45.425 163.715 ;
        RECT 45.215 163.635 45.425 163.645 ;
        RECT 42.920 163.305 44.455 163.555 ;
        RECT 44.625 163.135 44.955 163.615 ;
        RECT 45.170 163.305 45.425 163.635 ;
        RECT 46.135 163.135 46.415 163.615 ;
        RECT 46.585 163.395 46.845 163.785 ;
        RECT 47.020 163.135 47.275 163.615 ;
        RECT 47.445 163.395 47.740 163.785 ;
        RECT 48.495 163.635 48.665 164.545 ;
        RECT 47.920 163.135 48.195 163.615 ;
        RECT 48.365 163.305 48.665 163.635 ;
        RECT 48.840 164.545 49.175 165.515 ;
        RECT 49.345 164.545 49.515 165.685 ;
        RECT 49.685 165.345 51.715 165.515 ;
        RECT 48.840 163.875 49.010 164.545 ;
        RECT 49.685 164.375 49.855 165.345 ;
        RECT 49.180 164.045 49.435 164.375 ;
        RECT 49.660 164.045 49.855 164.375 ;
        RECT 50.025 165.005 51.150 165.175 ;
        RECT 49.265 163.875 49.435 164.045 ;
        RECT 50.025 163.875 50.195 165.005 ;
        RECT 48.840 163.305 49.095 163.875 ;
        RECT 49.265 163.705 50.195 163.875 ;
        RECT 50.365 164.665 51.375 164.835 ;
        RECT 50.365 163.865 50.535 164.665 ;
        RECT 50.740 164.325 51.015 164.465 ;
        RECT 50.735 164.155 51.015 164.325 ;
        RECT 50.020 163.670 50.195 163.705 ;
        RECT 49.265 163.135 49.595 163.535 ;
        RECT 50.020 163.305 50.550 163.670 ;
        RECT 50.740 163.305 51.015 164.155 ;
        RECT 51.185 163.305 51.375 164.665 ;
        RECT 51.545 164.680 51.715 165.345 ;
        RECT 51.885 164.925 52.055 165.685 ;
        RECT 52.290 164.925 52.805 165.335 ;
        RECT 51.545 164.490 52.295 164.680 ;
        RECT 52.465 164.115 52.805 164.925 ;
        RECT 52.980 165.015 53.235 165.515 ;
        RECT 53.405 165.185 53.735 165.685 ;
        RECT 52.980 164.845 53.730 165.015 ;
        RECT 51.575 163.945 52.805 164.115 ;
        RECT 52.980 164.025 53.330 164.675 ;
        RECT 51.555 163.135 52.065 163.670 ;
        RECT 52.285 163.340 52.530 163.945 ;
        RECT 53.500 163.855 53.730 164.845 ;
        RECT 52.980 163.685 53.730 163.855 ;
        RECT 52.980 163.395 53.235 163.685 ;
        RECT 53.405 163.135 53.735 163.515 ;
        RECT 53.905 163.395 54.075 165.515 ;
        RECT 54.245 164.715 54.570 165.500 ;
        RECT 54.740 165.225 54.990 165.685 ;
        RECT 55.160 165.185 55.410 165.515 ;
        RECT 55.625 165.185 56.305 165.515 ;
        RECT 55.160 165.055 55.330 165.185 ;
        RECT 54.935 164.885 55.330 165.055 ;
        RECT 54.305 163.665 54.765 164.715 ;
        RECT 54.935 163.525 55.105 164.885 ;
        RECT 55.500 164.625 55.965 165.015 ;
        RECT 55.275 163.815 55.625 164.435 ;
        RECT 55.795 164.035 55.965 164.625 ;
        RECT 56.135 164.405 56.305 165.185 ;
        RECT 56.475 165.085 56.645 165.425 ;
        RECT 56.880 165.255 57.210 165.685 ;
        RECT 57.380 165.085 57.550 165.425 ;
        RECT 57.845 165.225 58.215 165.685 ;
        RECT 56.475 164.915 57.550 165.085 ;
        RECT 58.385 165.055 58.555 165.515 ;
        RECT 58.790 165.175 59.660 165.515 ;
        RECT 59.830 165.225 60.080 165.685 ;
        RECT 57.995 164.885 58.555 165.055 ;
        RECT 57.995 164.745 58.165 164.885 ;
        RECT 56.665 164.575 58.165 164.745 ;
        RECT 58.860 164.715 59.320 165.005 ;
        RECT 56.135 164.235 57.825 164.405 ;
        RECT 55.795 163.815 56.150 164.035 ;
        RECT 56.320 163.525 56.490 164.235 ;
        RECT 56.695 163.815 57.485 164.065 ;
        RECT 57.655 164.055 57.825 164.235 ;
        RECT 57.995 163.885 58.165 164.575 ;
        RECT 54.435 163.135 54.765 163.495 ;
        RECT 54.935 163.355 55.430 163.525 ;
        RECT 55.635 163.355 56.490 163.525 ;
        RECT 57.365 163.135 57.695 163.595 ;
        RECT 57.905 163.495 58.165 163.885 ;
        RECT 58.355 164.705 59.320 164.715 ;
        RECT 59.490 164.795 59.660 165.175 ;
        RECT 60.250 165.135 60.420 165.425 ;
        RECT 60.600 165.305 60.930 165.685 ;
        RECT 60.250 164.965 61.050 165.135 ;
        RECT 58.355 164.545 59.030 164.705 ;
        RECT 59.490 164.625 60.710 164.795 ;
        RECT 58.355 163.755 58.565 164.545 ;
        RECT 59.490 164.535 59.660 164.625 ;
        RECT 58.735 163.755 59.085 164.375 ;
        RECT 59.255 164.365 59.660 164.535 ;
        RECT 59.255 163.585 59.425 164.365 ;
        RECT 59.595 163.915 59.815 164.195 ;
        RECT 59.995 164.085 60.535 164.455 ;
        RECT 60.880 164.375 61.050 164.965 ;
        RECT 61.270 164.545 61.575 165.685 ;
        RECT 61.745 164.495 62.000 165.375 ;
        RECT 60.880 164.345 61.620 164.375 ;
        RECT 59.595 163.745 60.125 163.915 ;
        RECT 57.905 163.325 58.255 163.495 ;
        RECT 58.475 163.305 59.425 163.585 ;
        RECT 59.595 163.135 59.785 163.575 ;
        RECT 59.955 163.515 60.125 163.745 ;
        RECT 60.295 163.685 60.535 164.085 ;
        RECT 60.705 164.045 61.620 164.345 ;
        RECT 60.705 163.870 61.030 164.045 ;
        RECT 60.705 163.515 61.025 163.870 ;
        RECT 61.790 163.845 62.000 164.495 ;
        RECT 62.175 164.925 62.690 165.335 ;
        RECT 62.925 164.925 63.095 165.685 ;
        RECT 63.265 165.345 65.295 165.515 ;
        RECT 62.175 164.115 62.515 164.925 ;
        RECT 63.265 164.680 63.435 165.345 ;
        RECT 63.830 165.005 64.955 165.175 ;
        RECT 62.685 164.490 63.435 164.680 ;
        RECT 63.605 164.665 64.615 164.835 ;
        RECT 62.175 163.945 63.405 164.115 ;
        RECT 59.955 163.345 61.025 163.515 ;
        RECT 61.270 163.135 61.575 163.595 ;
        RECT 61.745 163.315 62.000 163.845 ;
        RECT 62.450 163.340 62.695 163.945 ;
        RECT 62.915 163.135 63.425 163.670 ;
        RECT 63.605 163.305 63.795 164.665 ;
        RECT 63.965 163.645 64.240 164.465 ;
        RECT 64.445 163.865 64.615 164.665 ;
        RECT 64.785 163.875 64.955 165.005 ;
        RECT 65.125 164.375 65.295 165.345 ;
        RECT 65.465 164.545 65.635 165.685 ;
        RECT 65.805 164.545 66.140 165.515 ;
        RECT 65.125 164.045 65.320 164.375 ;
        RECT 65.545 164.045 65.800 164.375 ;
        RECT 65.545 163.875 65.715 164.045 ;
        RECT 65.970 163.875 66.140 164.545 ;
        RECT 67.235 164.520 67.525 165.685 ;
        RECT 67.705 164.875 68.000 165.685 ;
        RECT 68.180 164.375 68.425 165.515 ;
        RECT 68.600 164.875 68.860 165.685 ;
        RECT 69.460 165.680 75.735 165.685 ;
        RECT 69.040 164.375 69.290 165.510 ;
        RECT 69.460 164.885 69.720 165.680 ;
        RECT 69.890 164.785 70.150 165.510 ;
        RECT 70.320 164.955 70.580 165.680 ;
        RECT 70.750 164.785 71.010 165.510 ;
        RECT 71.180 164.955 71.440 165.680 ;
        RECT 71.610 164.785 71.870 165.510 ;
        RECT 72.040 164.955 72.300 165.680 ;
        RECT 72.470 164.785 72.730 165.510 ;
        RECT 72.900 164.955 73.145 165.680 ;
        RECT 73.315 164.785 73.575 165.510 ;
        RECT 73.760 164.955 74.005 165.680 ;
        RECT 74.175 164.785 74.435 165.510 ;
        RECT 74.620 164.955 74.865 165.680 ;
        RECT 75.035 164.785 75.295 165.510 ;
        RECT 75.480 164.955 75.735 165.680 ;
        RECT 69.890 164.770 75.295 164.785 ;
        RECT 75.905 164.770 76.195 165.510 ;
        RECT 76.365 164.940 76.635 165.685 ;
        RECT 69.890 164.545 76.635 164.770 ;
        RECT 76.895 164.595 78.565 165.685 ;
        RECT 64.785 163.705 65.715 163.875 ;
        RECT 64.785 163.670 64.960 163.705 ;
        RECT 63.965 163.475 64.245 163.645 ;
        RECT 63.965 163.305 64.240 163.475 ;
        RECT 64.430 163.305 64.960 163.670 ;
        RECT 65.385 163.135 65.715 163.535 ;
        RECT 65.885 163.305 66.140 163.875 ;
        RECT 67.235 163.135 67.525 163.860 ;
        RECT 67.695 163.815 68.010 164.375 ;
        RECT 68.180 164.125 75.300 164.375 ;
        RECT 67.695 163.135 68.000 163.645 ;
        RECT 68.180 163.315 68.430 164.125 ;
        RECT 68.600 163.135 68.860 163.660 ;
        RECT 69.040 163.315 69.290 164.125 ;
        RECT 75.470 163.955 76.635 164.545 ;
        RECT 69.890 163.785 76.635 163.955 ;
        RECT 76.895 163.905 77.645 164.425 ;
        RECT 77.815 164.075 78.565 164.595 ;
        RECT 78.735 164.925 79.250 165.335 ;
        RECT 79.485 164.925 79.655 165.685 ;
        RECT 79.825 165.345 81.855 165.515 ;
        RECT 78.735 164.115 79.075 164.925 ;
        RECT 79.825 164.680 79.995 165.345 ;
        RECT 80.390 165.005 81.515 165.175 ;
        RECT 79.245 164.490 79.995 164.680 ;
        RECT 80.165 164.665 81.175 164.835 ;
        RECT 78.735 163.945 79.965 164.115 ;
        RECT 69.460 163.135 69.720 163.695 ;
        RECT 69.890 163.330 70.150 163.785 ;
        RECT 70.320 163.135 70.580 163.615 ;
        RECT 70.750 163.330 71.010 163.785 ;
        RECT 71.180 163.135 71.440 163.615 ;
        RECT 71.610 163.330 71.870 163.785 ;
        RECT 72.040 163.135 72.285 163.615 ;
        RECT 72.455 163.330 72.730 163.785 ;
        RECT 72.900 163.135 73.145 163.615 ;
        RECT 73.315 163.330 73.575 163.785 ;
        RECT 73.755 163.135 74.005 163.615 ;
        RECT 74.175 163.330 74.435 163.785 ;
        RECT 74.615 163.135 74.865 163.615 ;
        RECT 75.035 163.330 75.295 163.785 ;
        RECT 75.475 163.135 75.735 163.615 ;
        RECT 75.905 163.330 76.165 163.785 ;
        RECT 76.335 163.135 76.635 163.615 ;
        RECT 76.895 163.135 78.565 163.905 ;
        RECT 79.010 163.340 79.255 163.945 ;
        RECT 79.475 163.135 79.985 163.670 ;
        RECT 80.165 163.305 80.355 164.665 ;
        RECT 80.525 164.325 80.800 164.465 ;
        RECT 80.525 164.155 80.805 164.325 ;
        RECT 80.525 163.305 80.800 164.155 ;
        RECT 81.005 163.865 81.175 164.665 ;
        RECT 81.345 163.875 81.515 165.005 ;
        RECT 81.685 164.375 81.855 165.345 ;
        RECT 82.025 164.545 82.195 165.685 ;
        RECT 82.365 164.545 82.700 165.515 ;
        RECT 81.685 164.045 81.880 164.375 ;
        RECT 82.105 164.045 82.360 164.375 ;
        RECT 82.105 163.875 82.275 164.045 ;
        RECT 82.530 163.875 82.700 164.545 ;
        RECT 81.345 163.705 82.275 163.875 ;
        RECT 81.345 163.670 81.520 163.705 ;
        RECT 80.990 163.305 81.520 163.670 ;
        RECT 81.945 163.135 82.275 163.535 ;
        RECT 82.445 163.305 82.700 163.875 ;
        RECT 82.875 164.715 83.185 165.515 ;
        RECT 83.355 164.885 83.665 165.685 ;
        RECT 83.835 165.055 84.095 165.515 ;
        RECT 84.265 165.225 84.520 165.685 ;
        RECT 84.695 165.055 84.955 165.515 ;
        RECT 83.835 164.885 84.955 165.055 ;
        RECT 82.875 164.545 83.905 164.715 ;
        RECT 82.875 163.635 83.045 164.545 ;
        RECT 83.215 163.805 83.565 164.375 ;
        RECT 83.735 164.295 83.905 164.545 ;
        RECT 84.695 164.635 84.955 164.885 ;
        RECT 85.125 164.815 85.410 165.685 ;
        RECT 84.695 164.465 85.450 164.635 ;
        RECT 85.640 164.535 85.900 165.685 ;
        RECT 86.075 164.610 86.330 165.515 ;
        RECT 86.500 164.925 86.830 165.685 ;
        RECT 87.045 164.755 87.215 165.515 ;
        RECT 83.735 164.125 84.875 164.295 ;
        RECT 85.045 163.955 85.450 164.465 ;
        RECT 83.800 163.785 85.450 163.955 ;
        RECT 82.875 163.305 83.175 163.635 ;
        RECT 83.345 163.135 83.620 163.615 ;
        RECT 83.800 163.395 84.095 163.785 ;
        RECT 84.265 163.135 84.520 163.615 ;
        RECT 84.695 163.395 84.955 163.785 ;
        RECT 85.125 163.135 85.405 163.615 ;
        RECT 85.640 163.135 85.900 163.975 ;
        RECT 86.075 163.880 86.245 164.610 ;
        RECT 86.500 164.585 87.215 164.755 ;
        RECT 86.500 164.375 86.670 164.585 ;
        RECT 88.455 164.545 88.665 165.685 ;
        RECT 88.835 164.535 89.165 165.515 ;
        RECT 89.335 164.545 89.565 165.685 ;
        RECT 90.275 164.545 90.505 165.685 ;
        RECT 90.675 164.535 91.005 165.515 ;
        RECT 91.175 164.545 91.385 165.685 ;
        RECT 91.625 164.545 91.955 165.685 ;
        RECT 92.485 164.715 92.815 165.500 ;
        RECT 92.135 164.545 92.815 164.715 ;
        RECT 86.415 164.045 86.670 164.375 ;
        RECT 86.075 163.305 86.330 163.880 ;
        RECT 86.500 163.855 86.670 164.045 ;
        RECT 86.950 164.035 87.305 164.405 ;
        RECT 86.500 163.685 87.215 163.855 ;
        RECT 86.500 163.135 86.830 163.515 ;
        RECT 87.045 163.305 87.215 163.685 ;
        RECT 88.455 163.135 88.665 163.955 ;
        RECT 88.835 163.935 89.085 164.535 ;
        RECT 89.255 164.125 89.585 164.375 ;
        RECT 90.255 164.125 90.585 164.375 ;
        RECT 88.835 163.305 89.165 163.935 ;
        RECT 89.335 163.135 89.565 163.955 ;
        RECT 90.275 163.135 90.505 163.955 ;
        RECT 90.755 163.935 91.005 164.535 ;
        RECT 91.615 164.125 91.965 164.375 ;
        RECT 90.675 163.305 91.005 163.935 ;
        RECT 91.175 163.135 91.385 163.955 ;
        RECT 92.135 163.945 92.305 164.545 ;
        RECT 92.995 164.520 93.285 165.685 ;
        RECT 93.765 164.845 93.935 165.685 ;
        RECT 94.145 164.675 94.395 165.515 ;
        RECT 94.605 164.845 94.775 165.685 ;
        RECT 94.945 164.675 95.235 165.515 ;
        RECT 93.510 164.505 95.235 164.675 ;
        RECT 95.445 164.625 95.615 165.685 ;
        RECT 95.910 165.305 96.240 165.685 ;
        RECT 96.420 165.135 96.590 165.425 ;
        RECT 96.760 165.225 97.010 165.685 ;
        RECT 95.790 164.965 96.590 165.135 ;
        RECT 97.180 165.175 98.050 165.515 ;
        RECT 92.475 164.125 92.825 164.375 ;
        RECT 93.510 163.955 93.920 164.505 ;
        RECT 95.790 164.345 95.960 164.965 ;
        RECT 97.180 164.795 97.350 165.175 ;
        RECT 98.285 165.055 98.455 165.515 ;
        RECT 98.625 165.225 98.995 165.685 ;
        RECT 99.290 165.085 99.460 165.425 ;
        RECT 99.630 165.255 99.960 165.685 ;
        RECT 100.195 165.085 100.365 165.425 ;
        RECT 96.130 164.625 97.350 164.795 ;
        RECT 97.520 164.715 97.980 165.005 ;
        RECT 98.285 164.885 98.845 165.055 ;
        RECT 99.290 164.915 100.365 165.085 ;
        RECT 100.535 165.185 101.215 165.515 ;
        RECT 101.430 165.185 101.680 165.515 ;
        RECT 101.850 165.225 102.100 165.685 ;
        RECT 98.675 164.745 98.845 164.885 ;
        RECT 97.520 164.705 98.485 164.715 ;
        RECT 97.180 164.535 97.350 164.625 ;
        RECT 97.810 164.545 98.485 164.705 ;
        RECT 95.790 164.335 96.135 164.345 ;
        RECT 94.105 164.125 96.135 164.335 ;
        RECT 91.625 163.135 91.895 163.945 ;
        RECT 92.065 163.305 92.395 163.945 ;
        RECT 92.565 163.135 92.805 163.945 ;
        RECT 92.995 163.135 93.285 163.860 ;
        RECT 93.510 163.785 95.275 163.955 ;
        RECT 93.765 163.135 93.935 163.605 ;
        RECT 94.105 163.305 94.435 163.785 ;
        RECT 94.605 163.135 94.775 163.605 ;
        RECT 94.945 163.305 95.275 163.785 ;
        RECT 95.445 163.135 95.615 163.945 ;
        RECT 95.810 163.870 96.135 164.125 ;
        RECT 95.815 163.515 96.135 163.870 ;
        RECT 96.305 164.085 96.845 164.455 ;
        RECT 97.180 164.365 97.585 164.535 ;
        RECT 96.305 163.685 96.545 164.085 ;
        RECT 97.025 163.915 97.245 164.195 ;
        RECT 96.715 163.745 97.245 163.915 ;
        RECT 96.715 163.515 96.885 163.745 ;
        RECT 97.415 163.585 97.585 164.365 ;
        RECT 97.755 163.755 98.105 164.375 ;
        RECT 98.275 163.755 98.485 164.545 ;
        RECT 98.675 164.575 100.175 164.745 ;
        RECT 98.675 163.885 98.845 164.575 ;
        RECT 100.535 164.405 100.705 165.185 ;
        RECT 101.510 165.055 101.680 165.185 ;
        RECT 99.015 164.235 100.705 164.405 ;
        RECT 100.875 164.625 101.340 165.015 ;
        RECT 101.510 164.885 101.905 165.055 ;
        RECT 99.015 164.055 99.185 164.235 ;
        RECT 95.815 163.345 96.885 163.515 ;
        RECT 97.055 163.135 97.245 163.575 ;
        RECT 97.415 163.305 98.365 163.585 ;
        RECT 98.675 163.495 98.935 163.885 ;
        RECT 99.355 163.815 100.145 164.065 ;
        RECT 98.585 163.325 98.935 163.495 ;
        RECT 99.145 163.135 99.475 163.595 ;
        RECT 100.350 163.525 100.520 164.235 ;
        RECT 100.875 164.035 101.045 164.625 ;
        RECT 100.690 163.815 101.045 164.035 ;
        RECT 101.215 163.815 101.565 164.435 ;
        RECT 101.735 163.525 101.905 164.885 ;
        RECT 102.270 164.715 102.595 165.500 ;
        RECT 102.075 163.665 102.535 164.715 ;
        RECT 100.350 163.355 101.205 163.525 ;
        RECT 101.410 163.355 101.905 163.525 ;
        RECT 102.075 163.135 102.405 163.495 ;
        RECT 102.765 163.395 102.935 165.515 ;
        RECT 103.105 165.185 103.435 165.685 ;
        RECT 103.605 165.015 103.860 165.515 ;
        RECT 103.110 164.845 103.860 165.015 ;
        RECT 103.110 163.855 103.340 164.845 ;
        RECT 103.510 164.025 103.860 164.675 ;
        RECT 104.495 164.545 104.880 165.515 ;
        RECT 105.050 165.225 105.375 165.685 ;
        RECT 105.895 165.055 106.175 165.515 ;
        RECT 105.050 164.835 106.175 165.055 ;
        RECT 104.495 163.875 104.775 164.545 ;
        RECT 105.050 164.375 105.500 164.835 ;
        RECT 106.365 164.665 106.765 165.515 ;
        RECT 107.165 165.225 107.435 165.685 ;
        RECT 107.605 165.055 107.890 165.515 ;
        RECT 104.945 164.045 105.500 164.375 ;
        RECT 105.670 164.105 106.765 164.665 ;
        RECT 105.050 163.935 105.500 164.045 ;
        RECT 103.110 163.685 103.860 163.855 ;
        RECT 103.105 163.135 103.435 163.515 ;
        RECT 103.605 163.395 103.860 163.685 ;
        RECT 104.495 163.305 104.880 163.875 ;
        RECT 105.050 163.765 106.175 163.935 ;
        RECT 105.050 163.135 105.375 163.595 ;
        RECT 105.895 163.305 106.175 163.765 ;
        RECT 106.365 163.305 106.765 164.105 ;
        RECT 106.935 164.835 107.890 165.055 ;
        RECT 108.485 164.845 108.655 165.685 ;
        RECT 106.935 163.935 107.145 164.835 ;
        RECT 108.865 164.675 109.115 165.515 ;
        RECT 109.325 164.845 109.495 165.685 ;
        RECT 109.665 164.675 109.955 165.515 ;
        RECT 107.315 164.105 108.005 164.665 ;
        RECT 108.230 164.505 109.955 164.675 ;
        RECT 110.165 164.625 110.335 165.685 ;
        RECT 110.630 165.305 110.960 165.685 ;
        RECT 111.140 165.135 111.310 165.425 ;
        RECT 111.480 165.225 111.730 165.685 ;
        RECT 110.510 164.965 111.310 165.135 ;
        RECT 111.900 165.175 112.770 165.515 ;
        RECT 108.230 163.955 108.640 164.505 ;
        RECT 110.510 164.345 110.680 164.965 ;
        RECT 111.900 164.795 112.070 165.175 ;
        RECT 113.005 165.055 113.175 165.515 ;
        RECT 113.345 165.225 113.715 165.685 ;
        RECT 114.010 165.085 114.180 165.425 ;
        RECT 114.350 165.255 114.680 165.685 ;
        RECT 114.915 165.085 115.085 165.425 ;
        RECT 110.850 164.625 112.070 164.795 ;
        RECT 112.240 164.715 112.700 165.005 ;
        RECT 113.005 164.885 113.565 165.055 ;
        RECT 114.010 164.915 115.085 165.085 ;
        RECT 115.255 165.185 115.935 165.515 ;
        RECT 116.150 165.185 116.400 165.515 ;
        RECT 116.570 165.225 116.820 165.685 ;
        RECT 113.395 164.745 113.565 164.885 ;
        RECT 112.240 164.705 113.205 164.715 ;
        RECT 111.900 164.535 112.070 164.625 ;
        RECT 112.530 164.545 113.205 164.705 ;
        RECT 110.510 164.335 110.855 164.345 ;
        RECT 108.825 164.125 110.855 164.335 ;
        RECT 106.935 163.765 107.890 163.935 ;
        RECT 108.230 163.785 109.995 163.955 ;
        RECT 107.165 163.135 107.435 163.595 ;
        RECT 107.605 163.305 107.890 163.765 ;
        RECT 108.485 163.135 108.655 163.605 ;
        RECT 108.825 163.305 109.155 163.785 ;
        RECT 109.325 163.135 109.495 163.605 ;
        RECT 109.665 163.305 109.995 163.785 ;
        RECT 110.165 163.135 110.335 163.945 ;
        RECT 110.530 163.870 110.855 164.125 ;
        RECT 110.535 163.515 110.855 163.870 ;
        RECT 111.025 164.085 111.565 164.455 ;
        RECT 111.900 164.365 112.305 164.535 ;
        RECT 111.025 163.685 111.265 164.085 ;
        RECT 111.745 163.915 111.965 164.195 ;
        RECT 111.435 163.745 111.965 163.915 ;
        RECT 111.435 163.515 111.605 163.745 ;
        RECT 112.135 163.585 112.305 164.365 ;
        RECT 112.475 163.755 112.825 164.375 ;
        RECT 112.995 163.755 113.205 164.545 ;
        RECT 113.395 164.575 114.895 164.745 ;
        RECT 113.395 163.885 113.565 164.575 ;
        RECT 115.255 164.405 115.425 165.185 ;
        RECT 116.230 165.055 116.400 165.185 ;
        RECT 113.735 164.235 115.425 164.405 ;
        RECT 115.595 164.625 116.060 165.015 ;
        RECT 116.230 164.885 116.625 165.055 ;
        RECT 113.735 164.055 113.905 164.235 ;
        RECT 110.535 163.345 111.605 163.515 ;
        RECT 111.775 163.135 111.965 163.575 ;
        RECT 112.135 163.305 113.085 163.585 ;
        RECT 113.395 163.495 113.655 163.885 ;
        RECT 114.075 163.815 114.865 164.065 ;
        RECT 113.305 163.325 113.655 163.495 ;
        RECT 113.865 163.135 114.195 163.595 ;
        RECT 115.070 163.525 115.240 164.235 ;
        RECT 115.595 164.035 115.765 164.625 ;
        RECT 115.410 163.815 115.765 164.035 ;
        RECT 115.935 163.815 116.285 164.435 ;
        RECT 116.455 163.525 116.625 164.885 ;
        RECT 116.990 164.715 117.315 165.500 ;
        RECT 116.795 163.665 117.255 164.715 ;
        RECT 115.070 163.355 115.925 163.525 ;
        RECT 116.130 163.355 116.625 163.525 ;
        RECT 116.795 163.135 117.125 163.495 ;
        RECT 117.485 163.395 117.655 165.515 ;
        RECT 117.825 165.185 118.155 165.685 ;
        RECT 118.325 165.015 118.580 165.515 ;
        RECT 117.830 164.845 118.580 165.015 ;
        RECT 117.830 163.855 118.060 164.845 ;
        RECT 118.230 164.025 118.580 164.675 ;
        RECT 118.755 164.520 119.045 165.685 ;
        RECT 119.215 164.715 119.525 165.515 ;
        RECT 119.695 164.885 120.005 165.685 ;
        RECT 120.175 165.055 120.435 165.515 ;
        RECT 120.605 165.225 120.860 165.685 ;
        RECT 121.035 165.055 121.295 165.515 ;
        RECT 120.175 164.885 121.295 165.055 ;
        RECT 119.215 164.545 120.245 164.715 ;
        RECT 117.830 163.685 118.580 163.855 ;
        RECT 117.825 163.135 118.155 163.515 ;
        RECT 118.325 163.395 118.580 163.685 ;
        RECT 118.755 163.135 119.045 163.860 ;
        RECT 119.215 163.635 119.385 164.545 ;
        RECT 119.555 163.805 119.905 164.375 ;
        RECT 120.075 164.295 120.245 164.545 ;
        RECT 121.035 164.635 121.295 164.885 ;
        RECT 121.465 164.815 121.750 165.685 ;
        RECT 121.035 164.465 121.790 164.635 ;
        RECT 122.485 164.545 122.735 165.685 ;
        RECT 120.075 164.125 121.215 164.295 ;
        RECT 121.385 163.955 121.790 164.465 ;
        RECT 120.140 163.785 121.790 163.955 ;
        RECT 122.905 164.495 123.155 165.375 ;
        RECT 123.325 164.545 123.630 165.685 ;
        RECT 123.970 165.305 124.300 165.685 ;
        RECT 124.480 165.135 124.650 165.425 ;
        RECT 124.820 165.225 125.070 165.685 ;
        RECT 123.850 164.965 124.650 165.135 ;
        RECT 125.240 165.175 126.110 165.515 ;
        RECT 119.215 163.305 119.515 163.635 ;
        RECT 119.685 163.135 119.960 163.615 ;
        RECT 120.140 163.395 120.435 163.785 ;
        RECT 120.605 163.135 120.860 163.615 ;
        RECT 121.035 163.395 121.295 163.785 ;
        RECT 121.465 163.135 121.745 163.615 ;
        RECT 122.485 163.135 122.735 163.890 ;
        RECT 122.905 163.845 123.110 164.495 ;
        RECT 123.850 164.375 124.020 164.965 ;
        RECT 125.240 164.795 125.410 165.175 ;
        RECT 126.345 165.055 126.515 165.515 ;
        RECT 126.685 165.225 127.055 165.685 ;
        RECT 127.350 165.085 127.520 165.425 ;
        RECT 127.690 165.255 128.020 165.685 ;
        RECT 128.255 165.085 128.425 165.425 ;
        RECT 124.190 164.625 125.410 164.795 ;
        RECT 125.580 164.715 126.040 165.005 ;
        RECT 126.345 164.885 126.905 165.055 ;
        RECT 127.350 164.915 128.425 165.085 ;
        RECT 128.595 165.185 129.275 165.515 ;
        RECT 129.490 165.185 129.740 165.515 ;
        RECT 129.910 165.225 130.160 165.685 ;
        RECT 126.735 164.745 126.905 164.885 ;
        RECT 125.580 164.705 126.545 164.715 ;
        RECT 125.240 164.535 125.410 164.625 ;
        RECT 125.870 164.545 126.545 164.705 ;
        RECT 123.280 164.345 124.020 164.375 ;
        RECT 123.280 164.045 124.195 164.345 ;
        RECT 123.870 163.870 124.195 164.045 ;
        RECT 122.905 163.315 123.155 163.845 ;
        RECT 123.325 163.135 123.630 163.595 ;
        RECT 123.875 163.515 124.195 163.870 ;
        RECT 124.365 164.085 124.905 164.455 ;
        RECT 125.240 164.365 125.645 164.535 ;
        RECT 124.365 163.685 124.605 164.085 ;
        RECT 125.085 163.915 125.305 164.195 ;
        RECT 124.775 163.745 125.305 163.915 ;
        RECT 124.775 163.515 124.945 163.745 ;
        RECT 125.475 163.585 125.645 164.365 ;
        RECT 125.815 163.755 126.165 164.375 ;
        RECT 126.335 163.755 126.545 164.545 ;
        RECT 126.735 164.575 128.235 164.745 ;
        RECT 126.735 163.885 126.905 164.575 ;
        RECT 128.595 164.405 128.765 165.185 ;
        RECT 129.570 165.055 129.740 165.185 ;
        RECT 127.075 164.235 128.765 164.405 ;
        RECT 128.935 164.625 129.400 165.015 ;
        RECT 129.570 164.885 129.965 165.055 ;
        RECT 127.075 164.055 127.245 164.235 ;
        RECT 123.875 163.345 124.945 163.515 ;
        RECT 125.115 163.135 125.305 163.575 ;
        RECT 125.475 163.305 126.425 163.585 ;
        RECT 126.735 163.495 126.995 163.885 ;
        RECT 127.415 163.815 128.205 164.065 ;
        RECT 126.645 163.325 126.995 163.495 ;
        RECT 127.205 163.135 127.535 163.595 ;
        RECT 128.410 163.525 128.580 164.235 ;
        RECT 128.935 164.035 129.105 164.625 ;
        RECT 128.750 163.815 129.105 164.035 ;
        RECT 129.275 163.815 129.625 164.435 ;
        RECT 129.795 163.525 129.965 164.885 ;
        RECT 130.330 164.715 130.655 165.500 ;
        RECT 130.135 163.665 130.595 164.715 ;
        RECT 128.410 163.355 129.265 163.525 ;
        RECT 129.470 163.355 129.965 163.525 ;
        RECT 130.135 163.135 130.465 163.495 ;
        RECT 130.825 163.395 130.995 165.515 ;
        RECT 131.165 165.185 131.495 165.685 ;
        RECT 131.665 165.015 131.920 165.515 ;
        RECT 131.170 164.845 131.920 165.015 ;
        RECT 131.170 163.855 131.400 164.845 ;
        RECT 131.570 164.025 131.920 164.675 ;
        RECT 132.145 164.545 132.395 165.685 ;
        RECT 132.565 164.495 132.815 165.375 ;
        RECT 132.985 164.545 133.290 165.685 ;
        RECT 133.630 165.305 133.960 165.685 ;
        RECT 134.140 165.135 134.310 165.425 ;
        RECT 134.480 165.225 134.730 165.685 ;
        RECT 133.510 164.965 134.310 165.135 ;
        RECT 134.900 165.175 135.770 165.515 ;
        RECT 131.170 163.685 131.920 163.855 ;
        RECT 131.165 163.135 131.495 163.515 ;
        RECT 131.665 163.395 131.920 163.685 ;
        RECT 132.145 163.135 132.395 163.890 ;
        RECT 132.565 163.845 132.770 164.495 ;
        RECT 133.510 164.375 133.680 164.965 ;
        RECT 134.900 164.795 135.070 165.175 ;
        RECT 136.005 165.055 136.175 165.515 ;
        RECT 136.345 165.225 136.715 165.685 ;
        RECT 137.010 165.085 137.180 165.425 ;
        RECT 137.350 165.255 137.680 165.685 ;
        RECT 137.915 165.085 138.085 165.425 ;
        RECT 133.850 164.625 135.070 164.795 ;
        RECT 135.240 164.715 135.700 165.005 ;
        RECT 136.005 164.885 136.565 165.055 ;
        RECT 137.010 164.915 138.085 165.085 ;
        RECT 138.255 165.185 138.935 165.515 ;
        RECT 139.150 165.185 139.400 165.515 ;
        RECT 139.570 165.225 139.820 165.685 ;
        RECT 136.395 164.745 136.565 164.885 ;
        RECT 135.240 164.705 136.205 164.715 ;
        RECT 134.900 164.535 135.070 164.625 ;
        RECT 135.530 164.545 136.205 164.705 ;
        RECT 132.940 164.345 133.680 164.375 ;
        RECT 132.940 164.045 133.855 164.345 ;
        RECT 133.530 163.870 133.855 164.045 ;
        RECT 132.565 163.315 132.815 163.845 ;
        RECT 132.985 163.135 133.290 163.595 ;
        RECT 133.535 163.515 133.855 163.870 ;
        RECT 134.025 164.085 134.565 164.455 ;
        RECT 134.900 164.365 135.305 164.535 ;
        RECT 134.025 163.685 134.265 164.085 ;
        RECT 134.745 163.915 134.965 164.195 ;
        RECT 134.435 163.745 134.965 163.915 ;
        RECT 134.435 163.515 134.605 163.745 ;
        RECT 135.135 163.585 135.305 164.365 ;
        RECT 135.475 163.755 135.825 164.375 ;
        RECT 135.995 163.755 136.205 164.545 ;
        RECT 136.395 164.575 137.895 164.745 ;
        RECT 136.395 163.885 136.565 164.575 ;
        RECT 138.255 164.405 138.425 165.185 ;
        RECT 139.230 165.055 139.400 165.185 ;
        RECT 136.735 164.235 138.425 164.405 ;
        RECT 138.595 164.625 139.060 165.015 ;
        RECT 139.230 164.885 139.625 165.055 ;
        RECT 136.735 164.055 136.905 164.235 ;
        RECT 133.535 163.345 134.605 163.515 ;
        RECT 134.775 163.135 134.965 163.575 ;
        RECT 135.135 163.305 136.085 163.585 ;
        RECT 136.395 163.495 136.655 163.885 ;
        RECT 137.075 163.815 137.865 164.065 ;
        RECT 136.305 163.325 136.655 163.495 ;
        RECT 136.865 163.135 137.195 163.595 ;
        RECT 138.070 163.525 138.240 164.235 ;
        RECT 138.595 164.035 138.765 164.625 ;
        RECT 138.410 163.815 138.765 164.035 ;
        RECT 138.935 163.815 139.285 164.435 ;
        RECT 139.455 163.525 139.625 164.885 ;
        RECT 139.990 164.715 140.315 165.500 ;
        RECT 139.795 163.665 140.255 164.715 ;
        RECT 138.070 163.355 138.925 163.525 ;
        RECT 139.130 163.355 139.625 163.525 ;
        RECT 139.795 163.135 140.125 163.495 ;
        RECT 140.485 163.395 140.655 165.515 ;
        RECT 140.825 165.185 141.155 165.685 ;
        RECT 141.325 165.015 141.580 165.515 ;
        RECT 140.830 164.845 141.580 165.015 ;
        RECT 140.830 163.855 141.060 164.845 ;
        RECT 141.230 164.025 141.580 164.675 ;
        RECT 141.755 164.595 144.345 165.685 ;
        RECT 141.755 163.905 142.965 164.425 ;
        RECT 143.135 164.075 144.345 164.595 ;
        RECT 144.515 164.520 144.805 165.685 ;
        RECT 145.030 164.815 145.315 165.685 ;
        RECT 145.485 165.055 145.745 165.515 ;
        RECT 145.920 165.225 146.175 165.685 ;
        RECT 146.345 165.055 146.605 165.515 ;
        RECT 145.485 164.885 146.605 165.055 ;
        RECT 146.775 164.885 147.085 165.685 ;
        RECT 145.485 164.635 145.745 164.885 ;
        RECT 147.255 164.715 147.565 165.515 ;
        RECT 144.990 164.465 145.745 164.635 ;
        RECT 146.535 164.545 147.565 164.715 ;
        RECT 144.990 163.955 145.395 164.465 ;
        RECT 146.535 164.295 146.705 164.545 ;
        RECT 145.565 164.125 146.705 164.295 ;
        RECT 140.830 163.685 141.580 163.855 ;
        RECT 140.825 163.135 141.155 163.515 ;
        RECT 141.325 163.395 141.580 163.685 ;
        RECT 141.755 163.135 144.345 163.905 ;
        RECT 144.515 163.135 144.805 163.860 ;
        RECT 144.990 163.785 146.640 163.955 ;
        RECT 146.875 163.805 147.225 164.375 ;
        RECT 145.035 163.135 145.315 163.615 ;
        RECT 145.485 163.395 145.745 163.785 ;
        RECT 145.920 163.135 146.175 163.615 ;
        RECT 146.345 163.395 146.640 163.785 ;
        RECT 147.395 163.635 147.565 164.545 ;
        RECT 147.740 164.535 148.000 165.685 ;
        RECT 148.175 164.610 148.430 165.515 ;
        RECT 148.600 164.925 148.930 165.685 ;
        RECT 149.145 164.755 149.315 165.515 ;
        RECT 149.575 165.250 154.920 165.685 ;
        RECT 146.820 163.135 147.095 163.615 ;
        RECT 147.265 163.305 147.565 163.635 ;
        RECT 147.740 163.135 148.000 163.975 ;
        RECT 148.175 163.880 148.345 164.610 ;
        RECT 148.600 164.585 149.315 164.755 ;
        RECT 148.600 164.375 148.770 164.585 ;
        RECT 148.515 164.045 148.770 164.375 ;
        RECT 148.175 163.305 148.430 163.880 ;
        RECT 148.600 163.855 148.770 164.045 ;
        RECT 149.050 164.035 149.405 164.405 ;
        RECT 148.600 163.685 149.315 163.855 ;
        RECT 148.600 163.135 148.930 163.515 ;
        RECT 149.145 163.305 149.315 163.685 ;
        RECT 151.160 163.680 151.500 164.510 ;
        RECT 152.980 164.000 153.330 165.250 ;
        RECT 155.095 164.595 156.765 165.685 ;
        RECT 155.095 163.905 155.845 164.425 ;
        RECT 156.015 164.075 156.765 164.595 ;
        RECT 156.935 164.595 158.145 165.685 ;
        RECT 156.935 164.055 157.455 164.595 ;
        RECT 149.575 163.135 154.920 163.680 ;
        RECT 155.095 163.135 156.765 163.905 ;
        RECT 157.625 163.885 158.145 164.425 ;
        RECT 156.935 163.135 158.145 163.885 ;
        RECT 2.750 162.965 158.230 163.135 ;
        RECT 2.835 162.215 4.045 162.965 ;
        RECT 5.135 162.290 5.395 162.795 ;
        RECT 5.575 162.585 5.905 162.965 ;
        RECT 6.085 162.415 6.255 162.795 ;
        RECT 2.835 161.675 3.355 162.215 ;
        RECT 3.525 161.505 4.045 162.045 ;
        RECT 2.835 160.415 4.045 161.505 ;
        RECT 5.135 161.490 5.305 162.290 ;
        RECT 5.590 162.245 6.255 162.415 ;
        RECT 5.590 161.990 5.760 162.245 ;
        RECT 6.520 162.225 6.775 162.795 ;
        RECT 6.945 162.565 7.275 162.965 ;
        RECT 7.700 162.430 8.230 162.795 ;
        RECT 7.700 162.395 7.875 162.430 ;
        RECT 6.945 162.225 7.875 162.395 ;
        RECT 5.475 161.660 5.760 161.990 ;
        RECT 5.995 161.695 6.325 162.065 ;
        RECT 5.590 161.515 5.760 161.660 ;
        RECT 6.520 161.555 6.690 162.225 ;
        RECT 6.945 162.055 7.115 162.225 ;
        RECT 6.860 161.725 7.115 162.055 ;
        RECT 7.340 161.725 7.535 162.055 ;
        RECT 5.135 160.585 5.405 161.490 ;
        RECT 5.590 161.345 6.255 161.515 ;
        RECT 5.575 160.415 5.905 161.175 ;
        RECT 6.085 160.585 6.255 161.345 ;
        RECT 6.520 160.585 6.855 161.555 ;
        RECT 7.025 160.415 7.195 161.555 ;
        RECT 7.365 160.755 7.535 161.725 ;
        RECT 7.705 161.095 7.875 162.225 ;
        RECT 8.045 161.435 8.215 162.235 ;
        RECT 8.420 161.945 8.695 162.795 ;
        RECT 8.415 161.775 8.695 161.945 ;
        RECT 8.420 161.635 8.695 161.775 ;
        RECT 8.865 161.435 9.055 162.795 ;
        RECT 9.235 162.430 9.745 162.965 ;
        RECT 9.965 162.155 10.210 162.760 ;
        RECT 10.660 162.415 10.915 162.705 ;
        RECT 11.085 162.585 11.415 162.965 ;
        RECT 10.660 162.245 11.410 162.415 ;
        RECT 9.255 161.985 10.485 162.155 ;
        RECT 8.045 161.265 9.055 161.435 ;
        RECT 9.225 161.420 9.975 161.610 ;
        RECT 7.705 160.925 8.830 161.095 ;
        RECT 9.225 160.755 9.395 161.420 ;
        RECT 10.145 161.175 10.485 161.985 ;
        RECT 10.660 161.425 11.010 162.075 ;
        RECT 11.180 161.255 11.410 162.245 ;
        RECT 7.365 160.585 9.395 160.755 ;
        RECT 9.565 160.415 9.735 161.175 ;
        RECT 9.970 160.765 10.485 161.175 ;
        RECT 10.660 161.085 11.410 161.255 ;
        RECT 10.660 160.585 10.915 161.085 ;
        RECT 11.085 160.415 11.415 160.915 ;
        RECT 11.585 160.585 11.755 162.705 ;
        RECT 12.115 162.605 12.445 162.965 ;
        RECT 12.615 162.575 13.110 162.745 ;
        RECT 13.315 162.575 14.170 162.745 ;
        RECT 11.985 161.385 12.445 162.435 ;
        RECT 11.925 160.600 12.250 161.385 ;
        RECT 12.615 161.215 12.785 162.575 ;
        RECT 12.955 161.665 13.305 162.285 ;
        RECT 13.475 162.065 13.830 162.285 ;
        RECT 13.475 161.475 13.645 162.065 ;
        RECT 14.000 161.865 14.170 162.575 ;
        RECT 15.045 162.505 15.375 162.965 ;
        RECT 15.585 162.605 15.935 162.775 ;
        RECT 14.375 162.035 15.165 162.285 ;
        RECT 15.585 162.215 15.845 162.605 ;
        RECT 16.155 162.515 17.105 162.795 ;
        RECT 17.275 162.525 17.465 162.965 ;
        RECT 17.635 162.585 18.705 162.755 ;
        RECT 15.335 161.865 15.505 162.045 ;
        RECT 12.615 161.045 13.010 161.215 ;
        RECT 13.180 161.085 13.645 161.475 ;
        RECT 13.815 161.695 15.505 161.865 ;
        RECT 12.840 160.915 13.010 161.045 ;
        RECT 13.815 160.915 13.985 161.695 ;
        RECT 15.675 161.525 15.845 162.215 ;
        RECT 14.345 161.355 15.845 161.525 ;
        RECT 16.035 161.555 16.245 162.345 ;
        RECT 16.415 161.725 16.765 162.345 ;
        RECT 16.935 161.735 17.105 162.515 ;
        RECT 17.635 162.355 17.805 162.585 ;
        RECT 17.275 162.185 17.805 162.355 ;
        RECT 17.275 161.905 17.495 162.185 ;
        RECT 17.975 162.015 18.215 162.415 ;
        RECT 16.935 161.565 17.340 161.735 ;
        RECT 17.675 161.645 18.215 162.015 ;
        RECT 18.385 162.230 18.705 162.585 ;
        RECT 18.950 162.505 19.255 162.965 ;
        RECT 19.425 162.255 19.680 162.785 ;
        RECT 18.385 162.055 18.710 162.230 ;
        RECT 18.385 161.755 19.300 162.055 ;
        RECT 18.560 161.725 19.300 161.755 ;
        RECT 16.035 161.395 16.710 161.555 ;
        RECT 17.170 161.475 17.340 161.565 ;
        RECT 16.035 161.385 17.000 161.395 ;
        RECT 15.675 161.215 15.845 161.355 ;
        RECT 12.420 160.415 12.670 160.875 ;
        RECT 12.840 160.585 13.090 160.915 ;
        RECT 13.305 160.585 13.985 160.915 ;
        RECT 14.155 161.015 15.230 161.185 ;
        RECT 15.675 161.045 16.235 161.215 ;
        RECT 16.540 161.095 17.000 161.385 ;
        RECT 17.170 161.305 18.390 161.475 ;
        RECT 14.155 160.675 14.325 161.015 ;
        RECT 14.560 160.415 14.890 160.845 ;
        RECT 15.060 160.675 15.230 161.015 ;
        RECT 15.525 160.415 15.895 160.875 ;
        RECT 16.065 160.585 16.235 161.045 ;
        RECT 17.170 160.925 17.340 161.305 ;
        RECT 18.560 161.135 18.730 161.725 ;
        RECT 19.470 161.605 19.680 162.255 ;
        RECT 16.470 160.585 17.340 160.925 ;
        RECT 17.930 160.965 18.730 161.135 ;
        RECT 17.510 160.415 17.760 160.875 ;
        RECT 17.930 160.675 18.100 160.965 ;
        RECT 18.280 160.415 18.610 160.795 ;
        RECT 18.950 160.415 19.255 161.555 ;
        RECT 19.425 160.725 19.680 161.605 ;
        RECT 19.855 162.225 20.240 162.795 ;
        RECT 20.410 162.505 20.735 162.965 ;
        RECT 21.255 162.335 21.535 162.795 ;
        RECT 19.855 161.555 20.135 162.225 ;
        RECT 20.410 162.165 21.535 162.335 ;
        RECT 20.410 162.055 20.860 162.165 ;
        RECT 20.305 161.725 20.860 162.055 ;
        RECT 21.725 161.995 22.125 162.795 ;
        RECT 22.525 162.505 22.795 162.965 ;
        RECT 22.965 162.335 23.250 162.795 ;
        RECT 19.855 160.585 20.240 161.555 ;
        RECT 20.410 161.265 20.860 161.725 ;
        RECT 21.030 161.435 22.125 161.995 ;
        RECT 20.410 161.045 21.535 161.265 ;
        RECT 20.410 160.415 20.735 160.875 ;
        RECT 21.255 160.585 21.535 161.045 ;
        RECT 21.725 160.585 22.125 161.435 ;
        RECT 22.295 162.165 23.250 162.335 ;
        RECT 23.540 162.200 23.995 162.965 ;
        RECT 24.270 162.585 25.570 162.795 ;
        RECT 25.825 162.605 26.155 162.965 ;
        RECT 25.400 162.435 25.570 162.585 ;
        RECT 26.325 162.465 26.585 162.795 ;
        RECT 26.355 162.455 26.585 162.465 ;
        RECT 22.295 161.265 22.505 162.165 ;
        RECT 22.675 161.435 23.365 161.995 ;
        RECT 24.470 161.975 24.690 162.375 ;
        RECT 23.535 161.775 24.025 161.975 ;
        RECT 24.215 161.765 24.690 161.975 ;
        RECT 24.935 161.975 25.145 162.375 ;
        RECT 25.400 162.310 26.155 162.435 ;
        RECT 25.400 162.265 26.245 162.310 ;
        RECT 25.975 162.145 26.245 162.265 ;
        RECT 24.935 161.765 25.265 161.975 ;
        RECT 25.435 161.705 25.845 162.010 ;
        RECT 23.540 161.535 24.715 161.595 ;
        RECT 26.075 161.570 26.245 162.145 ;
        RECT 26.045 161.535 26.245 161.570 ;
        RECT 23.540 161.425 26.245 161.535 ;
        RECT 22.295 161.045 23.250 161.265 ;
        RECT 22.525 160.415 22.795 160.875 ;
        RECT 22.965 160.585 23.250 161.045 ;
        RECT 23.540 160.805 23.795 161.425 ;
        RECT 24.385 161.365 26.185 161.425 ;
        RECT 24.385 161.335 24.715 161.365 ;
        RECT 26.415 161.265 26.585 162.455 ;
        RECT 26.755 162.195 28.425 162.965 ;
        RECT 28.595 162.240 28.885 162.965 ;
        RECT 29.975 162.505 30.535 162.795 ;
        RECT 30.705 162.505 30.955 162.965 ;
        RECT 26.755 161.675 27.505 162.195 ;
        RECT 27.675 161.505 28.425 162.025 ;
        RECT 24.045 161.165 24.230 161.255 ;
        RECT 24.820 161.165 25.655 161.175 ;
        RECT 24.045 160.965 25.655 161.165 ;
        RECT 24.045 160.925 24.275 160.965 ;
        RECT 23.540 160.585 23.875 160.805 ;
        RECT 24.880 160.415 25.235 160.795 ;
        RECT 25.405 160.585 25.655 160.965 ;
        RECT 25.905 160.415 26.155 161.195 ;
        RECT 26.325 160.585 26.585 161.265 ;
        RECT 26.755 160.415 28.425 161.505 ;
        RECT 28.595 160.415 28.885 161.580 ;
        RECT 29.975 161.135 30.225 162.505 ;
        RECT 31.575 162.335 31.905 162.695 ;
        RECT 32.365 162.485 32.665 162.965 ;
        RECT 30.515 162.145 31.905 162.335 ;
        RECT 32.835 162.315 33.095 162.770 ;
        RECT 33.265 162.485 33.525 162.965 ;
        RECT 33.705 162.315 33.965 162.770 ;
        RECT 34.135 162.485 34.385 162.965 ;
        RECT 34.565 162.315 34.825 162.770 ;
        RECT 34.995 162.485 35.245 162.965 ;
        RECT 35.425 162.315 35.685 162.770 ;
        RECT 35.855 162.485 36.100 162.965 ;
        RECT 36.270 162.315 36.545 162.770 ;
        RECT 36.715 162.485 36.960 162.965 ;
        RECT 37.130 162.315 37.390 162.770 ;
        RECT 37.560 162.485 37.820 162.965 ;
        RECT 37.990 162.315 38.250 162.770 ;
        RECT 38.420 162.485 38.680 162.965 ;
        RECT 38.850 162.315 39.110 162.770 ;
        RECT 39.280 162.405 39.540 162.965 ;
        RECT 32.365 162.145 39.110 162.315 ;
        RECT 30.515 162.055 30.685 162.145 ;
        RECT 30.395 161.725 30.685 162.055 ;
        RECT 30.855 161.725 31.195 161.975 ;
        RECT 31.415 161.725 32.090 161.975 ;
        RECT 30.515 161.475 30.685 161.725 ;
        RECT 30.515 161.305 31.455 161.475 ;
        RECT 31.825 161.365 32.090 161.725 ;
        RECT 32.365 161.555 33.530 162.145 ;
        RECT 39.710 161.975 39.960 162.785 ;
        RECT 40.140 162.440 40.400 162.965 ;
        RECT 40.570 161.975 40.820 162.785 ;
        RECT 41.000 162.455 41.305 162.965 ;
        RECT 33.700 161.725 40.820 161.975 ;
        RECT 40.990 161.725 41.305 162.285 ;
        RECT 41.480 162.255 41.735 162.785 ;
        RECT 41.905 162.505 42.210 162.965 ;
        RECT 42.455 162.585 43.525 162.755 ;
        RECT 32.365 161.330 39.110 161.555 ;
        RECT 29.975 160.585 30.435 161.135 ;
        RECT 30.625 160.415 30.955 161.135 ;
        RECT 31.155 160.755 31.455 161.305 ;
        RECT 31.625 160.415 31.905 161.085 ;
        RECT 32.365 160.415 32.635 161.160 ;
        RECT 32.805 160.590 33.095 161.330 ;
        RECT 33.705 161.315 39.110 161.330 ;
        RECT 33.265 160.420 33.520 161.145 ;
        RECT 33.705 160.590 33.965 161.315 ;
        RECT 34.135 160.420 34.380 161.145 ;
        RECT 34.565 160.590 34.825 161.315 ;
        RECT 34.995 160.420 35.240 161.145 ;
        RECT 35.425 160.590 35.685 161.315 ;
        RECT 35.855 160.420 36.100 161.145 ;
        RECT 36.270 160.590 36.530 161.315 ;
        RECT 36.700 160.420 36.960 161.145 ;
        RECT 37.130 160.590 37.390 161.315 ;
        RECT 37.560 160.420 37.820 161.145 ;
        RECT 37.990 160.590 38.250 161.315 ;
        RECT 38.420 160.420 38.680 161.145 ;
        RECT 38.850 160.590 39.110 161.315 ;
        RECT 39.280 160.420 39.540 161.215 ;
        RECT 39.710 160.590 39.960 161.725 ;
        RECT 33.265 160.415 39.540 160.420 ;
        RECT 40.140 160.415 40.400 161.225 ;
        RECT 40.575 160.585 40.820 161.725 ;
        RECT 41.480 161.605 41.690 162.255 ;
        RECT 42.455 162.230 42.775 162.585 ;
        RECT 42.450 162.055 42.775 162.230 ;
        RECT 41.860 161.755 42.775 162.055 ;
        RECT 42.945 162.015 43.185 162.415 ;
        RECT 43.355 162.355 43.525 162.585 ;
        RECT 43.695 162.525 43.885 162.965 ;
        RECT 44.055 162.515 45.005 162.795 ;
        RECT 45.225 162.605 45.575 162.775 ;
        RECT 43.355 162.185 43.885 162.355 ;
        RECT 41.860 161.725 42.600 161.755 ;
        RECT 41.000 160.415 41.295 161.225 ;
        RECT 41.480 160.725 41.735 161.605 ;
        RECT 41.905 160.415 42.210 161.555 ;
        RECT 42.430 161.135 42.600 161.725 ;
        RECT 42.945 161.645 43.485 162.015 ;
        RECT 43.665 161.905 43.885 162.185 ;
        RECT 44.055 161.735 44.225 162.515 ;
        RECT 43.820 161.565 44.225 161.735 ;
        RECT 44.395 161.725 44.745 162.345 ;
        RECT 43.820 161.475 43.990 161.565 ;
        RECT 44.915 161.555 45.125 162.345 ;
        RECT 42.770 161.305 43.990 161.475 ;
        RECT 44.450 161.395 45.125 161.555 ;
        RECT 42.430 160.965 43.230 161.135 ;
        RECT 42.550 160.415 42.880 160.795 ;
        RECT 43.060 160.675 43.230 160.965 ;
        RECT 43.820 160.925 43.990 161.305 ;
        RECT 44.160 161.385 45.125 161.395 ;
        RECT 45.315 162.215 45.575 162.605 ;
        RECT 45.785 162.505 46.115 162.965 ;
        RECT 46.990 162.575 47.845 162.745 ;
        RECT 48.050 162.575 48.545 162.745 ;
        RECT 48.715 162.605 49.045 162.965 ;
        RECT 45.315 161.525 45.485 162.215 ;
        RECT 45.655 161.865 45.825 162.045 ;
        RECT 45.995 162.035 46.785 162.285 ;
        RECT 46.990 161.865 47.160 162.575 ;
        RECT 47.330 162.065 47.685 162.285 ;
        RECT 45.655 161.695 47.345 161.865 ;
        RECT 44.160 161.095 44.620 161.385 ;
        RECT 45.315 161.355 46.815 161.525 ;
        RECT 45.315 161.215 45.485 161.355 ;
        RECT 44.925 161.045 45.485 161.215 ;
        RECT 43.400 160.415 43.650 160.875 ;
        RECT 43.820 160.585 44.690 160.925 ;
        RECT 44.925 160.585 45.095 161.045 ;
        RECT 45.930 161.015 47.005 161.185 ;
        RECT 45.265 160.415 45.635 160.875 ;
        RECT 45.930 160.675 46.100 161.015 ;
        RECT 46.270 160.415 46.600 160.845 ;
        RECT 46.835 160.675 47.005 161.015 ;
        RECT 47.175 160.915 47.345 161.695 ;
        RECT 47.515 161.475 47.685 162.065 ;
        RECT 47.855 161.665 48.205 162.285 ;
        RECT 47.515 161.085 47.980 161.475 ;
        RECT 48.375 161.215 48.545 162.575 ;
        RECT 48.715 161.385 49.175 162.435 ;
        RECT 48.150 161.045 48.545 161.215 ;
        RECT 48.150 160.915 48.320 161.045 ;
        RECT 47.175 160.585 47.855 160.915 ;
        RECT 48.070 160.585 48.320 160.915 ;
        RECT 48.490 160.415 48.740 160.875 ;
        RECT 48.910 160.600 49.235 161.385 ;
        RECT 49.405 160.585 49.575 162.705 ;
        RECT 49.745 162.585 50.075 162.965 ;
        RECT 50.245 162.415 50.500 162.705 ;
        RECT 49.750 162.245 50.500 162.415 ;
        RECT 49.750 161.255 49.980 162.245 ;
        RECT 51.145 162.240 51.475 162.750 ;
        RECT 51.645 162.565 51.975 162.965 ;
        RECT 53.025 162.395 53.355 162.735 ;
        RECT 53.525 162.565 53.855 162.965 ;
        RECT 50.150 161.425 50.500 162.075 ;
        RECT 51.145 161.475 51.335 162.240 ;
        RECT 51.645 162.225 54.010 162.395 ;
        RECT 54.355 162.240 54.645 162.965 ;
        RECT 54.825 162.240 55.155 162.750 ;
        RECT 55.325 162.565 55.655 162.965 ;
        RECT 56.705 162.395 57.035 162.735 ;
        RECT 57.205 162.565 57.535 162.965 ;
        RECT 51.645 162.055 51.815 162.225 ;
        RECT 51.505 161.725 51.815 162.055 ;
        RECT 51.985 161.725 52.290 162.055 ;
        RECT 49.750 161.085 50.500 161.255 ;
        RECT 49.745 160.415 50.075 160.915 ;
        RECT 50.245 160.585 50.500 161.085 ;
        RECT 51.145 160.625 51.475 161.475 ;
        RECT 51.645 160.415 51.895 161.555 ;
        RECT 52.075 161.395 52.290 161.725 ;
        RECT 52.465 161.395 52.750 162.055 ;
        RECT 52.945 161.395 53.210 162.055 ;
        RECT 53.425 161.395 53.670 162.055 ;
        RECT 53.840 161.225 54.010 162.225 ;
        RECT 52.085 161.055 53.375 161.225 ;
        RECT 52.085 160.635 52.335 161.055 ;
        RECT 52.565 160.415 52.895 160.885 ;
        RECT 53.125 160.635 53.375 161.055 ;
        RECT 53.555 161.055 54.010 161.225 ;
        RECT 53.555 160.625 53.885 161.055 ;
        RECT 54.355 160.415 54.645 161.580 ;
        RECT 54.825 161.475 55.015 162.240 ;
        RECT 55.325 162.225 57.690 162.395 ;
        RECT 55.325 162.055 55.495 162.225 ;
        RECT 55.185 161.725 55.495 162.055 ;
        RECT 55.665 161.725 55.970 162.055 ;
        RECT 54.825 160.625 55.155 161.475 ;
        RECT 55.325 160.415 55.575 161.555 ;
        RECT 55.755 161.395 55.970 161.725 ;
        RECT 56.145 161.395 56.430 162.055 ;
        RECT 56.625 161.395 56.890 162.055 ;
        RECT 57.105 161.395 57.350 162.055 ;
        RECT 57.520 161.225 57.690 162.225 ;
        RECT 55.765 161.055 57.055 161.225 ;
        RECT 55.765 160.635 56.015 161.055 ;
        RECT 56.245 160.415 56.575 160.885 ;
        RECT 56.805 160.635 57.055 161.055 ;
        RECT 57.235 161.055 57.690 161.225 ;
        RECT 58.035 162.290 58.295 162.795 ;
        RECT 58.475 162.585 58.805 162.965 ;
        RECT 58.985 162.415 59.155 162.795 ;
        RECT 58.035 161.490 58.205 162.290 ;
        RECT 58.490 162.245 59.155 162.415 ;
        RECT 58.490 161.990 58.660 162.245 ;
        RECT 58.375 161.660 58.660 161.990 ;
        RECT 58.895 161.695 59.225 162.065 ;
        RECT 58.490 161.515 58.660 161.660 ;
        RECT 57.235 160.625 57.565 161.055 ;
        RECT 58.035 160.585 58.305 161.490 ;
        RECT 58.490 161.345 59.155 161.515 ;
        RECT 58.475 160.415 58.805 161.175 ;
        RECT 58.985 160.585 59.155 161.345 ;
        RECT 59.880 161.215 60.210 162.795 ;
        RECT 60.380 162.465 60.580 162.965 ;
        RECT 60.840 162.315 61.030 162.630 ;
        RECT 61.200 162.585 62.495 162.755 ;
        RECT 62.665 162.585 62.995 162.965 ;
        RECT 62.325 162.415 62.495 162.585 ;
        RECT 60.380 161.425 60.570 162.295 ;
        RECT 60.840 162.025 61.305 162.315 ;
        RECT 61.485 161.770 62.115 162.285 ;
        RECT 62.325 162.245 62.935 162.415 ;
        RECT 63.165 162.300 63.415 162.795 ;
        RECT 62.765 162.055 62.935 162.245 ;
        RECT 61.485 161.735 61.655 161.770 ;
        RECT 60.840 161.425 61.655 161.735 ;
        RECT 62.425 161.555 62.595 162.055 ;
        RECT 61.935 161.385 62.595 161.555 ;
        RECT 62.765 161.725 63.075 162.055 ;
        RECT 61.935 161.215 62.105 161.385 ;
        RECT 62.765 161.215 62.935 161.725 ;
        RECT 63.245 161.455 63.415 162.300 ;
        RECT 63.585 162.165 63.840 162.965 ;
        RECT 64.020 162.415 64.275 162.705 ;
        RECT 64.445 162.585 64.775 162.965 ;
        RECT 64.020 162.245 64.770 162.415 ;
        RECT 59.880 161.045 62.105 161.215 ;
        RECT 62.275 161.045 62.935 161.215 ;
        RECT 59.880 160.585 60.215 161.045 ;
        RECT 60.385 160.415 60.605 160.875 ;
        RECT 62.275 160.795 62.445 161.045 ;
        RECT 61.135 160.625 62.445 160.795 ;
        RECT 62.615 160.415 62.905 160.875 ;
        RECT 63.105 160.585 63.415 161.455 ;
        RECT 63.585 160.415 63.840 161.555 ;
        RECT 64.020 161.425 64.370 162.075 ;
        RECT 64.540 161.255 64.770 162.245 ;
        RECT 64.020 161.085 64.770 161.255 ;
        RECT 64.020 160.585 64.275 161.085 ;
        RECT 64.445 160.415 64.775 160.915 ;
        RECT 64.945 160.585 65.115 162.705 ;
        RECT 65.475 162.605 65.805 162.965 ;
        RECT 65.975 162.575 66.470 162.745 ;
        RECT 66.675 162.575 67.530 162.745 ;
        RECT 65.345 161.385 65.805 162.435 ;
        RECT 65.285 160.600 65.610 161.385 ;
        RECT 65.975 161.215 66.145 162.575 ;
        RECT 66.315 161.665 66.665 162.285 ;
        RECT 66.835 162.065 67.190 162.285 ;
        RECT 66.835 161.475 67.005 162.065 ;
        RECT 67.360 161.865 67.530 162.575 ;
        RECT 68.405 162.505 68.735 162.965 ;
        RECT 68.945 162.605 69.295 162.775 ;
        RECT 67.735 162.035 68.525 162.285 ;
        RECT 68.945 162.215 69.205 162.605 ;
        RECT 69.515 162.515 70.465 162.795 ;
        RECT 70.635 162.525 70.825 162.965 ;
        RECT 70.995 162.585 72.065 162.755 ;
        RECT 68.695 161.865 68.865 162.045 ;
        RECT 65.975 161.045 66.370 161.215 ;
        RECT 66.540 161.085 67.005 161.475 ;
        RECT 67.175 161.695 68.865 161.865 ;
        RECT 66.200 160.915 66.370 161.045 ;
        RECT 67.175 160.915 67.345 161.695 ;
        RECT 69.035 161.525 69.205 162.215 ;
        RECT 67.705 161.355 69.205 161.525 ;
        RECT 69.395 161.555 69.605 162.345 ;
        RECT 69.775 161.725 70.125 162.345 ;
        RECT 70.295 161.735 70.465 162.515 ;
        RECT 70.995 162.355 71.165 162.585 ;
        RECT 70.635 162.185 71.165 162.355 ;
        RECT 70.635 161.905 70.855 162.185 ;
        RECT 71.335 162.015 71.575 162.415 ;
        RECT 70.295 161.565 70.700 161.735 ;
        RECT 71.035 161.645 71.575 162.015 ;
        RECT 71.745 162.230 72.065 162.585 ;
        RECT 72.310 162.505 72.615 162.965 ;
        RECT 72.785 162.255 73.040 162.785 ;
        RECT 71.745 162.055 72.070 162.230 ;
        RECT 71.745 161.755 72.660 162.055 ;
        RECT 71.920 161.725 72.660 161.755 ;
        RECT 69.395 161.395 70.070 161.555 ;
        RECT 70.530 161.475 70.700 161.565 ;
        RECT 69.395 161.385 70.360 161.395 ;
        RECT 69.035 161.215 69.205 161.355 ;
        RECT 65.780 160.415 66.030 160.875 ;
        RECT 66.200 160.585 66.450 160.915 ;
        RECT 66.665 160.585 67.345 160.915 ;
        RECT 67.515 161.015 68.590 161.185 ;
        RECT 69.035 161.045 69.595 161.215 ;
        RECT 69.900 161.095 70.360 161.385 ;
        RECT 70.530 161.305 71.750 161.475 ;
        RECT 67.515 160.675 67.685 161.015 ;
        RECT 67.920 160.415 68.250 160.845 ;
        RECT 68.420 160.675 68.590 161.015 ;
        RECT 68.885 160.415 69.255 160.875 ;
        RECT 69.425 160.585 69.595 161.045 ;
        RECT 70.530 160.925 70.700 161.305 ;
        RECT 71.920 161.135 72.090 161.725 ;
        RECT 72.830 161.605 73.040 162.255 ;
        RECT 73.490 162.155 73.735 162.760 ;
        RECT 73.955 162.430 74.465 162.965 ;
        RECT 69.830 160.585 70.700 160.925 ;
        RECT 71.290 160.965 72.090 161.135 ;
        RECT 70.870 160.415 71.120 160.875 ;
        RECT 71.290 160.675 71.460 160.965 ;
        RECT 71.640 160.415 71.970 160.795 ;
        RECT 72.310 160.415 72.615 161.555 ;
        RECT 72.785 160.725 73.040 161.605 ;
        RECT 73.215 161.985 74.445 162.155 ;
        RECT 73.215 161.175 73.555 161.985 ;
        RECT 73.725 161.420 74.475 161.610 ;
        RECT 73.215 160.765 73.730 161.175 ;
        RECT 73.965 160.415 74.135 161.175 ;
        RECT 74.305 160.755 74.475 161.420 ;
        RECT 74.645 161.435 74.835 162.795 ;
        RECT 75.005 162.625 75.280 162.795 ;
        RECT 75.005 162.455 75.285 162.625 ;
        RECT 75.005 161.635 75.280 162.455 ;
        RECT 75.470 162.430 76.000 162.795 ;
        RECT 76.425 162.565 76.755 162.965 ;
        RECT 75.825 162.395 76.000 162.430 ;
        RECT 75.485 161.435 75.655 162.235 ;
        RECT 74.645 161.265 75.655 161.435 ;
        RECT 75.825 162.225 76.755 162.395 ;
        RECT 76.925 162.225 77.180 162.795 ;
        RECT 77.415 162.485 77.695 162.965 ;
        RECT 77.865 162.315 78.125 162.705 ;
        RECT 78.300 162.485 78.555 162.965 ;
        RECT 78.725 162.315 79.020 162.705 ;
        RECT 79.200 162.485 79.475 162.965 ;
        RECT 79.645 162.465 79.945 162.795 ;
        RECT 75.825 161.095 75.995 162.225 ;
        RECT 76.585 162.055 76.755 162.225 ;
        RECT 74.870 160.925 75.995 161.095 ;
        RECT 76.165 161.725 76.360 162.055 ;
        RECT 76.585 161.725 76.840 162.055 ;
        RECT 76.165 160.755 76.335 161.725 ;
        RECT 77.010 161.555 77.180 162.225 ;
        RECT 74.305 160.585 76.335 160.755 ;
        RECT 76.505 160.415 76.675 161.555 ;
        RECT 76.845 160.585 77.180 161.555 ;
        RECT 77.370 162.145 79.020 162.315 ;
        RECT 77.370 161.635 77.775 162.145 ;
        RECT 77.945 161.805 79.085 161.975 ;
        RECT 77.370 161.465 78.125 161.635 ;
        RECT 77.410 160.415 77.695 161.285 ;
        RECT 77.865 161.215 78.125 161.465 ;
        RECT 78.915 161.555 79.085 161.805 ;
        RECT 79.255 161.725 79.605 162.295 ;
        RECT 79.775 161.555 79.945 162.465 ;
        RECT 80.115 162.240 80.405 162.965 ;
        RECT 80.850 162.155 81.095 162.760 ;
        RECT 81.315 162.430 81.825 162.965 ;
        RECT 80.575 161.985 81.805 162.155 ;
        RECT 78.915 161.385 79.945 161.555 ;
        RECT 77.865 161.045 78.985 161.215 ;
        RECT 77.865 160.585 78.125 161.045 ;
        RECT 78.300 160.415 78.555 160.875 ;
        RECT 78.725 160.585 78.985 161.045 ;
        RECT 79.155 160.415 79.465 161.215 ;
        RECT 79.635 160.585 79.945 161.385 ;
        RECT 80.115 160.415 80.405 161.580 ;
        RECT 80.575 161.175 80.915 161.985 ;
        RECT 81.085 161.420 81.835 161.610 ;
        RECT 80.575 160.765 81.090 161.175 ;
        RECT 81.325 160.415 81.495 161.175 ;
        RECT 81.665 160.755 81.835 161.420 ;
        RECT 82.005 161.435 82.195 162.795 ;
        RECT 82.365 161.945 82.640 162.795 ;
        RECT 82.830 162.430 83.360 162.795 ;
        RECT 83.785 162.565 84.115 162.965 ;
        RECT 83.185 162.395 83.360 162.430 ;
        RECT 82.365 161.775 82.645 161.945 ;
        RECT 82.365 161.635 82.640 161.775 ;
        RECT 82.845 161.435 83.015 162.235 ;
        RECT 82.005 161.265 83.015 161.435 ;
        RECT 83.185 162.225 84.115 162.395 ;
        RECT 84.285 162.225 84.540 162.795 ;
        RECT 83.185 161.095 83.355 162.225 ;
        RECT 83.945 162.055 84.115 162.225 ;
        RECT 82.230 160.925 83.355 161.095 ;
        RECT 83.525 161.725 83.720 162.055 ;
        RECT 83.945 161.725 84.200 162.055 ;
        RECT 83.525 160.755 83.695 161.725 ;
        RECT 84.370 161.555 84.540 162.225 ;
        RECT 81.665 160.585 83.695 160.755 ;
        RECT 83.865 160.415 84.035 161.555 ;
        RECT 84.205 160.585 84.540 161.555 ;
        RECT 85.635 162.245 85.975 162.755 ;
        RECT 85.635 160.845 85.895 162.245 ;
        RECT 86.145 162.165 86.415 162.965 ;
        RECT 86.070 161.725 86.400 161.975 ;
        RECT 86.595 161.725 86.875 162.695 ;
        RECT 87.055 161.725 87.355 162.695 ;
        RECT 87.535 161.725 87.885 162.690 ;
        RECT 88.105 162.465 88.600 162.795 ;
        RECT 88.965 162.585 90.135 162.795 ;
        RECT 88.965 162.565 89.295 162.585 ;
        RECT 86.085 161.555 86.400 161.725 ;
        RECT 88.105 161.555 88.275 162.465 ;
        RECT 86.085 161.385 88.275 161.555 ;
        RECT 85.635 160.585 85.975 160.845 ;
        RECT 86.145 160.415 86.475 161.215 ;
        RECT 86.940 160.585 87.190 161.385 ;
        RECT 87.375 160.415 87.705 161.135 ;
        RECT 87.925 160.585 88.175 161.385 ;
        RECT 88.445 160.975 88.685 162.285 ;
        RECT 88.855 162.145 89.715 162.395 ;
        RECT 89.885 162.335 90.135 162.585 ;
        RECT 90.305 162.505 90.475 162.965 ;
        RECT 90.645 162.335 90.985 162.795 ;
        RECT 89.885 162.165 90.985 162.335 ;
        RECT 91.155 162.165 91.850 162.795 ;
        RECT 92.055 162.165 92.365 162.965 ;
        RECT 93.545 162.415 93.715 162.795 ;
        RECT 93.930 162.585 94.260 162.965 ;
        RECT 93.545 162.245 94.260 162.415 ;
        RECT 88.855 161.555 89.135 162.145 ;
        RECT 89.305 161.725 90.055 161.975 ;
        RECT 90.225 161.725 90.985 161.975 ;
        RECT 91.175 161.725 91.510 161.975 ;
        RECT 91.680 161.565 91.850 162.165 ;
        RECT 92.020 161.725 92.355 161.995 ;
        RECT 93.455 161.695 93.810 162.065 ;
        RECT 94.090 162.055 94.260 162.245 ;
        RECT 94.430 162.220 94.685 162.795 ;
        RECT 94.090 161.725 94.345 162.055 ;
        RECT 88.855 161.385 90.555 161.555 ;
        RECT 88.345 160.415 88.680 160.795 ;
        RECT 88.960 160.415 89.215 161.215 ;
        RECT 89.385 160.585 89.715 161.385 ;
        RECT 89.885 160.415 90.055 161.215 ;
        RECT 90.225 160.585 90.555 161.385 ;
        RECT 90.725 160.415 90.985 161.555 ;
        RECT 91.155 160.415 91.415 161.555 ;
        RECT 91.585 160.585 91.915 161.565 ;
        RECT 92.085 160.415 92.365 161.555 ;
        RECT 94.090 161.515 94.260 161.725 ;
        RECT 93.545 161.345 94.260 161.515 ;
        RECT 94.515 161.490 94.685 162.220 ;
        RECT 94.860 162.125 95.120 162.965 ;
        RECT 95.295 162.225 95.680 162.795 ;
        RECT 95.850 162.505 96.175 162.965 ;
        RECT 96.695 162.335 96.975 162.795 ;
        RECT 93.545 160.585 93.715 161.345 ;
        RECT 93.930 160.415 94.260 161.175 ;
        RECT 94.430 160.585 94.685 161.490 ;
        RECT 94.860 160.415 95.120 161.565 ;
        RECT 95.295 161.555 95.575 162.225 ;
        RECT 95.850 162.165 96.975 162.335 ;
        RECT 95.850 162.055 96.300 162.165 ;
        RECT 95.745 161.725 96.300 162.055 ;
        RECT 97.165 161.995 97.565 162.795 ;
        RECT 97.965 162.505 98.235 162.965 ;
        RECT 98.405 162.335 98.690 162.795 ;
        RECT 95.295 160.585 95.680 161.555 ;
        RECT 95.850 161.265 96.300 161.725 ;
        RECT 96.470 161.435 97.565 161.995 ;
        RECT 95.850 161.045 96.975 161.265 ;
        RECT 95.850 160.415 96.175 160.875 ;
        RECT 96.695 160.585 96.975 161.045 ;
        RECT 97.165 160.585 97.565 161.435 ;
        RECT 97.735 162.165 98.690 162.335 ;
        RECT 98.975 162.465 99.275 162.795 ;
        RECT 99.445 162.485 99.720 162.965 ;
        RECT 97.735 161.265 97.945 162.165 ;
        RECT 98.115 161.435 98.805 161.995 ;
        RECT 98.975 161.555 99.145 162.465 ;
        RECT 99.900 162.315 100.195 162.705 ;
        RECT 100.365 162.485 100.620 162.965 ;
        RECT 100.795 162.315 101.055 162.705 ;
        RECT 101.225 162.485 101.505 162.965 ;
        RECT 99.315 161.725 99.665 162.295 ;
        RECT 99.900 162.145 101.550 162.315 ;
        RECT 102.010 162.155 102.255 162.760 ;
        RECT 102.475 162.430 102.985 162.965 ;
        RECT 99.835 161.805 100.975 161.975 ;
        RECT 99.835 161.555 100.005 161.805 ;
        RECT 101.145 161.635 101.550 162.145 ;
        RECT 98.975 161.385 100.005 161.555 ;
        RECT 100.795 161.465 101.550 161.635 ;
        RECT 101.735 161.985 102.965 162.155 ;
        RECT 97.735 161.045 98.690 161.265 ;
        RECT 97.965 160.415 98.235 160.875 ;
        RECT 98.405 160.585 98.690 161.045 ;
        RECT 98.975 160.585 99.285 161.385 ;
        RECT 100.795 161.215 101.055 161.465 ;
        RECT 99.455 160.415 99.765 161.215 ;
        RECT 99.935 161.045 101.055 161.215 ;
        RECT 99.935 160.585 100.195 161.045 ;
        RECT 100.365 160.415 100.620 160.875 ;
        RECT 100.795 160.585 101.055 161.045 ;
        RECT 101.225 160.415 101.510 161.285 ;
        RECT 101.735 161.175 102.075 161.985 ;
        RECT 102.245 161.420 102.995 161.610 ;
        RECT 101.735 160.765 102.250 161.175 ;
        RECT 102.485 160.415 102.655 161.175 ;
        RECT 102.825 160.755 102.995 161.420 ;
        RECT 103.165 161.435 103.355 162.795 ;
        RECT 103.525 161.945 103.800 162.795 ;
        RECT 103.990 162.430 104.520 162.795 ;
        RECT 104.945 162.565 105.275 162.965 ;
        RECT 104.345 162.395 104.520 162.430 ;
        RECT 103.525 161.775 103.805 161.945 ;
        RECT 103.525 161.635 103.800 161.775 ;
        RECT 104.005 161.435 104.175 162.235 ;
        RECT 103.165 161.265 104.175 161.435 ;
        RECT 104.345 162.225 105.275 162.395 ;
        RECT 105.445 162.225 105.700 162.795 ;
        RECT 105.875 162.240 106.165 162.965 ;
        RECT 106.645 162.495 106.815 162.965 ;
        RECT 106.985 162.315 107.315 162.795 ;
        RECT 107.485 162.495 107.655 162.965 ;
        RECT 107.825 162.315 108.155 162.795 ;
        RECT 104.345 161.095 104.515 162.225 ;
        RECT 105.105 162.055 105.275 162.225 ;
        RECT 103.390 160.925 104.515 161.095 ;
        RECT 104.685 161.725 104.880 162.055 ;
        RECT 105.105 161.725 105.360 162.055 ;
        RECT 104.685 160.755 104.855 161.725 ;
        RECT 105.530 161.555 105.700 162.225 ;
        RECT 106.390 162.145 108.155 162.315 ;
        RECT 108.325 162.155 108.495 162.965 ;
        RECT 108.695 162.585 109.765 162.755 ;
        RECT 108.695 162.230 109.015 162.585 ;
        RECT 106.390 161.595 106.800 162.145 ;
        RECT 108.690 161.975 109.015 162.230 ;
        RECT 106.985 161.765 109.015 161.975 ;
        RECT 108.670 161.755 109.015 161.765 ;
        RECT 109.185 162.015 109.425 162.415 ;
        RECT 109.595 162.355 109.765 162.585 ;
        RECT 109.935 162.525 110.125 162.965 ;
        RECT 110.295 162.515 111.245 162.795 ;
        RECT 111.465 162.605 111.815 162.775 ;
        RECT 109.595 162.185 110.125 162.355 ;
        RECT 102.825 160.585 104.855 160.755 ;
        RECT 105.025 160.415 105.195 161.555 ;
        RECT 105.365 160.585 105.700 161.555 ;
        RECT 105.875 160.415 106.165 161.580 ;
        RECT 106.390 161.425 108.115 161.595 ;
        RECT 106.645 160.415 106.815 161.255 ;
        RECT 107.025 160.585 107.275 161.425 ;
        RECT 107.485 160.415 107.655 161.255 ;
        RECT 107.825 160.585 108.115 161.425 ;
        RECT 108.325 160.415 108.495 161.475 ;
        RECT 108.670 161.135 108.840 161.755 ;
        RECT 109.185 161.645 109.725 162.015 ;
        RECT 109.905 161.905 110.125 162.185 ;
        RECT 110.295 161.735 110.465 162.515 ;
        RECT 110.060 161.565 110.465 161.735 ;
        RECT 110.635 161.725 110.985 162.345 ;
        RECT 110.060 161.475 110.230 161.565 ;
        RECT 111.155 161.555 111.365 162.345 ;
        RECT 109.010 161.305 110.230 161.475 ;
        RECT 110.690 161.395 111.365 161.555 ;
        RECT 108.670 160.965 109.470 161.135 ;
        RECT 108.790 160.415 109.120 160.795 ;
        RECT 109.300 160.675 109.470 160.965 ;
        RECT 110.060 160.925 110.230 161.305 ;
        RECT 110.400 161.385 111.365 161.395 ;
        RECT 111.555 162.215 111.815 162.605 ;
        RECT 112.025 162.505 112.355 162.965 ;
        RECT 113.230 162.575 114.085 162.745 ;
        RECT 114.290 162.575 114.785 162.745 ;
        RECT 114.955 162.605 115.285 162.965 ;
        RECT 111.555 161.525 111.725 162.215 ;
        RECT 111.895 161.865 112.065 162.045 ;
        RECT 112.235 162.035 113.025 162.285 ;
        RECT 113.230 161.865 113.400 162.575 ;
        RECT 113.570 162.065 113.925 162.285 ;
        RECT 111.895 161.695 113.585 161.865 ;
        RECT 110.400 161.095 110.860 161.385 ;
        RECT 111.555 161.355 113.055 161.525 ;
        RECT 111.555 161.215 111.725 161.355 ;
        RECT 111.165 161.045 111.725 161.215 ;
        RECT 109.640 160.415 109.890 160.875 ;
        RECT 110.060 160.585 110.930 160.925 ;
        RECT 111.165 160.585 111.335 161.045 ;
        RECT 112.170 161.015 113.245 161.185 ;
        RECT 111.505 160.415 111.875 160.875 ;
        RECT 112.170 160.675 112.340 161.015 ;
        RECT 112.510 160.415 112.840 160.845 ;
        RECT 113.075 160.675 113.245 161.015 ;
        RECT 113.415 160.915 113.585 161.695 ;
        RECT 113.755 161.475 113.925 162.065 ;
        RECT 114.095 161.665 114.445 162.285 ;
        RECT 113.755 161.085 114.220 161.475 ;
        RECT 114.615 161.215 114.785 162.575 ;
        RECT 114.955 161.385 115.415 162.435 ;
        RECT 114.390 161.045 114.785 161.215 ;
        RECT 114.390 160.915 114.560 161.045 ;
        RECT 113.415 160.585 114.095 160.915 ;
        RECT 114.310 160.585 114.560 160.915 ;
        RECT 114.730 160.415 114.980 160.875 ;
        RECT 115.150 160.600 115.475 161.385 ;
        RECT 115.645 160.585 115.815 162.705 ;
        RECT 115.985 162.585 116.315 162.965 ;
        RECT 116.485 162.415 116.740 162.705 ;
        RECT 115.990 162.245 116.740 162.415 ;
        RECT 115.990 161.255 116.220 162.245 ;
        RECT 117.190 162.155 117.435 162.760 ;
        RECT 117.655 162.430 118.165 162.965 ;
        RECT 116.390 161.425 116.740 162.075 ;
        RECT 116.915 161.985 118.145 162.155 ;
        RECT 115.990 161.085 116.740 161.255 ;
        RECT 115.985 160.415 116.315 160.915 ;
        RECT 116.485 160.585 116.740 161.085 ;
        RECT 116.915 161.175 117.255 161.985 ;
        RECT 117.425 161.420 118.175 161.610 ;
        RECT 116.915 160.765 117.430 161.175 ;
        RECT 117.665 160.415 117.835 161.175 ;
        RECT 118.005 160.755 118.175 161.420 ;
        RECT 118.345 161.435 118.535 162.795 ;
        RECT 118.705 161.945 118.980 162.795 ;
        RECT 119.170 162.430 119.700 162.795 ;
        RECT 120.125 162.565 120.455 162.965 ;
        RECT 119.525 162.395 119.700 162.430 ;
        RECT 118.705 161.775 118.985 161.945 ;
        RECT 118.705 161.635 118.980 161.775 ;
        RECT 119.185 161.435 119.355 162.235 ;
        RECT 118.345 161.265 119.355 161.435 ;
        RECT 119.525 162.225 120.455 162.395 ;
        RECT 120.625 162.225 120.880 162.795 ;
        RECT 119.525 161.095 119.695 162.225 ;
        RECT 120.285 162.055 120.455 162.225 ;
        RECT 118.570 160.925 119.695 161.095 ;
        RECT 119.865 161.725 120.060 162.055 ;
        RECT 120.285 161.725 120.540 162.055 ;
        RECT 119.865 160.755 120.035 161.725 ;
        RECT 120.710 161.555 120.880 162.225 ;
        RECT 118.005 160.585 120.035 160.755 ;
        RECT 120.205 160.415 120.375 161.555 ;
        RECT 120.545 160.585 120.880 161.555 ;
        RECT 121.055 162.290 121.315 162.795 ;
        RECT 121.495 162.585 121.825 162.965 ;
        RECT 122.005 162.415 122.175 162.795 ;
        RECT 121.055 161.490 121.225 162.290 ;
        RECT 121.510 162.245 122.175 162.415 ;
        RECT 121.510 161.990 121.680 162.245 ;
        RECT 122.455 162.155 122.695 162.965 ;
        RECT 122.865 162.155 123.195 162.795 ;
        RECT 123.365 162.155 123.635 162.965 ;
        RECT 124.550 162.155 124.795 162.760 ;
        RECT 125.015 162.430 125.525 162.965 ;
        RECT 121.395 161.660 121.680 161.990 ;
        RECT 121.915 161.695 122.245 162.065 ;
        RECT 122.435 161.725 122.785 161.975 ;
        RECT 121.510 161.515 121.680 161.660 ;
        RECT 122.955 161.555 123.125 162.155 ;
        RECT 124.275 161.985 125.505 162.155 ;
        RECT 123.295 161.725 123.645 161.975 ;
        RECT 121.055 160.585 121.325 161.490 ;
        RECT 121.510 161.345 122.175 161.515 ;
        RECT 121.495 160.415 121.825 161.175 ;
        RECT 122.005 160.585 122.175 161.345 ;
        RECT 122.445 161.385 123.125 161.555 ;
        RECT 122.445 160.600 122.775 161.385 ;
        RECT 123.305 160.415 123.635 161.555 ;
        RECT 124.275 161.175 124.615 161.985 ;
        RECT 124.785 161.420 125.535 161.610 ;
        RECT 124.275 160.765 124.790 161.175 ;
        RECT 125.025 160.415 125.195 161.175 ;
        RECT 125.365 160.755 125.535 161.420 ;
        RECT 125.705 161.435 125.895 162.795 ;
        RECT 126.065 162.625 126.340 162.795 ;
        RECT 126.065 162.455 126.345 162.625 ;
        RECT 126.065 161.635 126.340 162.455 ;
        RECT 126.530 162.430 127.060 162.795 ;
        RECT 127.485 162.565 127.815 162.965 ;
        RECT 126.885 162.395 127.060 162.430 ;
        RECT 126.545 161.435 126.715 162.235 ;
        RECT 125.705 161.265 126.715 161.435 ;
        RECT 126.885 162.225 127.815 162.395 ;
        RECT 127.985 162.225 128.240 162.795 ;
        RECT 126.885 161.095 127.055 162.225 ;
        RECT 127.645 162.055 127.815 162.225 ;
        RECT 125.930 160.925 127.055 161.095 ;
        RECT 127.225 161.725 127.420 162.055 ;
        RECT 127.645 161.725 127.900 162.055 ;
        RECT 127.225 160.755 127.395 161.725 ;
        RECT 128.070 161.555 128.240 162.225 ;
        RECT 125.365 160.585 127.395 160.755 ;
        RECT 127.565 160.415 127.735 161.555 ;
        RECT 127.905 160.585 128.240 161.555 ;
        RECT 128.415 162.290 128.675 162.795 ;
        RECT 128.855 162.585 129.185 162.965 ;
        RECT 129.365 162.415 129.535 162.795 ;
        RECT 128.415 161.490 128.585 162.290 ;
        RECT 128.870 162.245 129.535 162.415 ;
        RECT 129.885 162.415 130.055 162.795 ;
        RECT 130.235 162.585 130.565 162.965 ;
        RECT 129.885 162.245 130.550 162.415 ;
        RECT 130.745 162.290 131.005 162.795 ;
        RECT 128.870 161.990 129.040 162.245 ;
        RECT 128.755 161.660 129.040 161.990 ;
        RECT 129.275 161.695 129.605 162.065 ;
        RECT 129.815 161.695 130.145 162.065 ;
        RECT 130.380 161.990 130.550 162.245 ;
        RECT 128.870 161.515 129.040 161.660 ;
        RECT 130.380 161.660 130.665 161.990 ;
        RECT 130.380 161.515 130.550 161.660 ;
        RECT 128.415 160.585 128.685 161.490 ;
        RECT 128.870 161.345 129.535 161.515 ;
        RECT 128.855 160.415 129.185 161.175 ;
        RECT 129.365 160.585 129.535 161.345 ;
        RECT 129.885 161.345 130.550 161.515 ;
        RECT 130.835 161.490 131.005 162.290 ;
        RECT 131.635 162.240 131.925 162.965 ;
        RECT 132.370 162.155 132.615 162.760 ;
        RECT 132.835 162.430 133.345 162.965 ;
        RECT 132.095 161.985 133.325 162.155 ;
        RECT 129.885 160.585 130.055 161.345 ;
        RECT 130.235 160.415 130.565 161.175 ;
        RECT 130.735 160.585 131.005 161.490 ;
        RECT 131.635 160.415 131.925 161.580 ;
        RECT 132.095 161.175 132.435 161.985 ;
        RECT 132.605 161.420 133.355 161.610 ;
        RECT 132.095 160.765 132.610 161.175 ;
        RECT 132.845 160.415 133.015 161.175 ;
        RECT 133.185 160.755 133.355 161.420 ;
        RECT 133.525 161.435 133.715 162.795 ;
        RECT 133.885 162.625 134.160 162.795 ;
        RECT 133.885 162.455 134.165 162.625 ;
        RECT 133.885 161.635 134.160 162.455 ;
        RECT 134.350 162.430 134.880 162.795 ;
        RECT 135.305 162.565 135.635 162.965 ;
        RECT 134.705 162.395 134.880 162.430 ;
        RECT 134.365 161.435 134.535 162.235 ;
        RECT 133.525 161.265 134.535 161.435 ;
        RECT 134.705 162.225 135.635 162.395 ;
        RECT 135.805 162.225 136.060 162.795 ;
        RECT 136.325 162.415 136.495 162.795 ;
        RECT 136.675 162.585 137.005 162.965 ;
        RECT 136.325 162.245 136.990 162.415 ;
        RECT 137.185 162.290 137.445 162.795 ;
        RECT 134.705 161.095 134.875 162.225 ;
        RECT 135.465 162.055 135.635 162.225 ;
        RECT 133.750 160.925 134.875 161.095 ;
        RECT 135.045 161.725 135.240 162.055 ;
        RECT 135.465 161.725 135.720 162.055 ;
        RECT 135.045 160.755 135.215 161.725 ;
        RECT 135.890 161.555 136.060 162.225 ;
        RECT 136.255 161.695 136.585 162.065 ;
        RECT 136.820 161.990 136.990 162.245 ;
        RECT 133.185 160.585 135.215 160.755 ;
        RECT 135.385 160.415 135.555 161.555 ;
        RECT 135.725 160.585 136.060 161.555 ;
        RECT 136.820 161.660 137.105 161.990 ;
        RECT 136.820 161.515 136.990 161.660 ;
        RECT 136.325 161.345 136.990 161.515 ;
        RECT 137.275 161.490 137.445 162.290 ;
        RECT 137.665 162.210 137.915 162.965 ;
        RECT 138.085 162.255 138.335 162.785 ;
        RECT 138.505 162.505 138.810 162.965 ;
        RECT 139.055 162.585 140.125 162.755 ;
        RECT 138.085 161.605 138.290 162.255 ;
        RECT 139.055 162.230 139.375 162.585 ;
        RECT 139.050 162.055 139.375 162.230 ;
        RECT 138.460 161.755 139.375 162.055 ;
        RECT 139.545 162.015 139.785 162.415 ;
        RECT 139.955 162.355 140.125 162.585 ;
        RECT 140.295 162.525 140.485 162.965 ;
        RECT 140.655 162.515 141.605 162.795 ;
        RECT 141.825 162.605 142.175 162.775 ;
        RECT 139.955 162.185 140.485 162.355 ;
        RECT 138.460 161.725 139.200 161.755 ;
        RECT 136.325 160.585 136.495 161.345 ;
        RECT 136.675 160.415 137.005 161.175 ;
        RECT 137.175 160.585 137.445 161.490 ;
        RECT 137.665 160.415 137.915 161.555 ;
        RECT 138.085 160.725 138.335 161.605 ;
        RECT 138.505 160.415 138.810 161.555 ;
        RECT 139.030 161.135 139.200 161.725 ;
        RECT 139.545 161.645 140.085 162.015 ;
        RECT 140.265 161.905 140.485 162.185 ;
        RECT 140.655 161.735 140.825 162.515 ;
        RECT 140.420 161.565 140.825 161.735 ;
        RECT 140.995 161.725 141.345 162.345 ;
        RECT 140.420 161.475 140.590 161.565 ;
        RECT 141.515 161.555 141.725 162.345 ;
        RECT 139.370 161.305 140.590 161.475 ;
        RECT 141.050 161.395 141.725 161.555 ;
        RECT 139.030 160.965 139.830 161.135 ;
        RECT 139.150 160.415 139.480 160.795 ;
        RECT 139.660 160.675 139.830 160.965 ;
        RECT 140.420 160.925 140.590 161.305 ;
        RECT 140.760 161.385 141.725 161.395 ;
        RECT 141.915 162.215 142.175 162.605 ;
        RECT 142.385 162.505 142.715 162.965 ;
        RECT 143.590 162.575 144.445 162.745 ;
        RECT 144.650 162.575 145.145 162.745 ;
        RECT 145.315 162.605 145.645 162.965 ;
        RECT 141.915 161.525 142.085 162.215 ;
        RECT 142.255 161.865 142.425 162.045 ;
        RECT 142.595 162.035 143.385 162.285 ;
        RECT 143.590 161.865 143.760 162.575 ;
        RECT 143.930 162.065 144.285 162.285 ;
        RECT 142.255 161.695 143.945 161.865 ;
        RECT 140.760 161.095 141.220 161.385 ;
        RECT 141.915 161.355 143.415 161.525 ;
        RECT 141.915 161.215 142.085 161.355 ;
        RECT 141.525 161.045 142.085 161.215 ;
        RECT 140.000 160.415 140.250 160.875 ;
        RECT 140.420 160.585 141.290 160.925 ;
        RECT 141.525 160.585 141.695 161.045 ;
        RECT 142.530 161.015 143.605 161.185 ;
        RECT 141.865 160.415 142.235 160.875 ;
        RECT 142.530 160.675 142.700 161.015 ;
        RECT 142.870 160.415 143.200 160.845 ;
        RECT 143.435 160.675 143.605 161.015 ;
        RECT 143.775 160.915 143.945 161.695 ;
        RECT 144.115 161.475 144.285 162.065 ;
        RECT 144.455 161.665 144.805 162.285 ;
        RECT 144.115 161.085 144.580 161.475 ;
        RECT 144.975 161.215 145.145 162.575 ;
        RECT 145.315 161.385 145.775 162.435 ;
        RECT 144.750 161.045 145.145 161.215 ;
        RECT 144.750 160.915 144.920 161.045 ;
        RECT 143.775 160.585 144.455 160.915 ;
        RECT 144.670 160.585 144.920 160.915 ;
        RECT 145.090 160.415 145.340 160.875 ;
        RECT 145.510 160.600 145.835 161.385 ;
        RECT 146.005 160.585 146.175 162.705 ;
        RECT 146.345 162.585 146.675 162.965 ;
        RECT 146.845 162.415 147.100 162.705 ;
        RECT 147.275 162.420 152.620 162.965 ;
        RECT 146.350 162.245 147.100 162.415 ;
        RECT 146.350 161.255 146.580 162.245 ;
        RECT 146.750 161.425 147.100 162.075 ;
        RECT 148.860 161.590 149.200 162.420 ;
        RECT 152.795 162.195 156.305 162.965 ;
        RECT 156.935 162.215 158.145 162.965 ;
        RECT 146.350 161.085 147.100 161.255 ;
        RECT 146.345 160.415 146.675 160.915 ;
        RECT 146.845 160.585 147.100 161.085 ;
        RECT 150.680 160.850 151.030 162.100 ;
        RECT 152.795 161.675 154.445 162.195 ;
        RECT 154.615 161.505 156.305 162.025 ;
        RECT 147.275 160.415 152.620 160.850 ;
        RECT 152.795 160.415 156.305 161.505 ;
        RECT 156.935 161.505 157.455 162.045 ;
        RECT 157.625 161.675 158.145 162.215 ;
        RECT 156.935 160.415 158.145 161.505 ;
        RECT 2.750 160.245 158.230 160.415 ;
        RECT 2.835 159.155 4.045 160.245 ;
        RECT 4.220 159.575 4.475 160.075 ;
        RECT 4.645 159.745 4.975 160.245 ;
        RECT 4.220 159.405 4.970 159.575 ;
        RECT 2.835 158.445 3.355 158.985 ;
        RECT 3.525 158.615 4.045 159.155 ;
        RECT 4.220 158.585 4.570 159.235 ;
        RECT 2.835 157.695 4.045 158.445 ;
        RECT 4.740 158.415 4.970 159.405 ;
        RECT 4.220 158.245 4.970 158.415 ;
        RECT 4.220 157.955 4.475 158.245 ;
        RECT 4.645 157.695 4.975 158.075 ;
        RECT 5.145 157.955 5.315 160.075 ;
        RECT 5.485 159.275 5.810 160.060 ;
        RECT 5.980 159.785 6.230 160.245 ;
        RECT 6.400 159.745 6.650 160.075 ;
        RECT 6.865 159.745 7.545 160.075 ;
        RECT 6.400 159.615 6.570 159.745 ;
        RECT 6.175 159.445 6.570 159.615 ;
        RECT 5.545 158.225 6.005 159.275 ;
        RECT 6.175 158.085 6.345 159.445 ;
        RECT 6.740 159.185 7.205 159.575 ;
        RECT 6.515 158.375 6.865 158.995 ;
        RECT 7.035 158.595 7.205 159.185 ;
        RECT 7.375 158.965 7.545 159.745 ;
        RECT 7.715 159.645 7.885 159.985 ;
        RECT 8.120 159.815 8.450 160.245 ;
        RECT 8.620 159.645 8.790 159.985 ;
        RECT 9.085 159.785 9.455 160.245 ;
        RECT 7.715 159.475 8.790 159.645 ;
        RECT 9.625 159.615 9.795 160.075 ;
        RECT 10.030 159.735 10.900 160.075 ;
        RECT 11.070 159.785 11.320 160.245 ;
        RECT 9.235 159.445 9.795 159.615 ;
        RECT 9.235 159.305 9.405 159.445 ;
        RECT 7.905 159.135 9.405 159.305 ;
        RECT 10.100 159.275 10.560 159.565 ;
        RECT 7.375 158.795 9.065 158.965 ;
        RECT 7.035 158.375 7.390 158.595 ;
        RECT 7.560 158.085 7.730 158.795 ;
        RECT 7.935 158.375 8.725 158.625 ;
        RECT 8.895 158.615 9.065 158.795 ;
        RECT 9.235 158.445 9.405 159.135 ;
        RECT 5.675 157.695 6.005 158.055 ;
        RECT 6.175 157.915 6.670 158.085 ;
        RECT 6.875 157.915 7.730 158.085 ;
        RECT 8.605 157.695 8.935 158.155 ;
        RECT 9.145 158.055 9.405 158.445 ;
        RECT 9.595 159.265 10.560 159.275 ;
        RECT 10.730 159.355 10.900 159.735 ;
        RECT 11.490 159.695 11.660 159.985 ;
        RECT 11.840 159.865 12.170 160.245 ;
        RECT 11.490 159.525 12.290 159.695 ;
        RECT 9.595 159.105 10.270 159.265 ;
        RECT 10.730 159.185 11.950 159.355 ;
        RECT 9.595 158.315 9.805 159.105 ;
        RECT 10.730 159.095 10.900 159.185 ;
        RECT 9.975 158.315 10.325 158.935 ;
        RECT 10.495 158.925 10.900 159.095 ;
        RECT 10.495 158.145 10.665 158.925 ;
        RECT 10.835 158.475 11.055 158.755 ;
        RECT 11.235 158.645 11.775 159.015 ;
        RECT 12.120 158.935 12.290 159.525 ;
        RECT 12.510 159.105 12.815 160.245 ;
        RECT 12.985 159.055 13.240 159.935 ;
        RECT 12.120 158.905 12.860 158.935 ;
        RECT 10.835 158.305 11.365 158.475 ;
        RECT 9.145 157.885 9.495 158.055 ;
        RECT 9.715 157.865 10.665 158.145 ;
        RECT 10.835 157.695 11.025 158.135 ;
        RECT 11.195 158.075 11.365 158.305 ;
        RECT 11.535 158.245 11.775 158.645 ;
        RECT 11.945 158.605 12.860 158.905 ;
        RECT 11.945 158.430 12.270 158.605 ;
        RECT 11.945 158.075 12.265 158.430 ;
        RECT 13.030 158.405 13.240 159.055 ;
        RECT 11.195 157.905 12.265 158.075 ;
        RECT 12.510 157.695 12.815 158.155 ;
        RECT 12.985 157.875 13.240 158.405 ;
        RECT 13.415 159.170 13.685 160.075 ;
        RECT 13.855 159.485 14.185 160.245 ;
        RECT 14.365 159.315 14.535 160.075 ;
        RECT 13.415 158.370 13.585 159.170 ;
        RECT 13.870 159.145 14.535 159.315 ;
        RECT 13.870 159.000 14.040 159.145 ;
        RECT 15.715 159.080 16.005 160.245 ;
        RECT 16.180 159.105 16.515 160.075 ;
        RECT 16.685 159.105 16.855 160.245 ;
        RECT 17.025 159.905 19.055 160.075 ;
        RECT 13.755 158.670 14.040 159.000 ;
        RECT 13.870 158.415 14.040 158.670 ;
        RECT 14.275 158.595 14.605 158.965 ;
        RECT 16.180 158.435 16.350 159.105 ;
        RECT 17.025 158.935 17.195 159.905 ;
        RECT 16.520 158.605 16.775 158.935 ;
        RECT 17.000 158.605 17.195 158.935 ;
        RECT 17.365 159.565 18.490 159.735 ;
        RECT 16.605 158.435 16.775 158.605 ;
        RECT 17.365 158.435 17.535 159.565 ;
        RECT 13.415 157.865 13.675 158.370 ;
        RECT 13.870 158.245 14.535 158.415 ;
        RECT 13.855 157.695 14.185 158.075 ;
        RECT 14.365 157.865 14.535 158.245 ;
        RECT 15.715 157.695 16.005 158.420 ;
        RECT 16.180 157.865 16.435 158.435 ;
        RECT 16.605 158.265 17.535 158.435 ;
        RECT 17.705 159.225 18.715 159.395 ;
        RECT 17.705 158.425 17.875 159.225 ;
        RECT 18.080 158.885 18.355 159.025 ;
        RECT 18.075 158.715 18.355 158.885 ;
        RECT 17.360 158.230 17.535 158.265 ;
        RECT 16.605 157.695 16.935 158.095 ;
        RECT 17.360 157.865 17.890 158.230 ;
        RECT 18.080 157.865 18.355 158.715 ;
        RECT 18.525 157.865 18.715 159.225 ;
        RECT 18.885 159.240 19.055 159.905 ;
        RECT 19.225 159.485 19.395 160.245 ;
        RECT 19.630 159.485 20.145 159.895 ;
        RECT 18.885 159.050 19.635 159.240 ;
        RECT 19.805 158.675 20.145 159.485 ;
        RECT 20.315 159.155 21.985 160.245 ;
        RECT 18.915 158.505 20.145 158.675 ;
        RECT 18.895 157.695 19.405 158.230 ;
        RECT 19.625 157.900 19.870 158.505 ;
        RECT 20.315 158.465 21.065 158.985 ;
        RECT 21.235 158.635 21.985 159.155 ;
        RECT 22.705 159.235 22.875 160.075 ;
        RECT 23.045 159.905 24.215 160.075 ;
        RECT 23.045 159.405 23.375 159.905 ;
        RECT 23.885 159.865 24.215 159.905 ;
        RECT 24.405 159.825 24.760 160.245 ;
        RECT 23.545 159.645 23.775 159.735 ;
        RECT 24.930 159.645 25.180 160.075 ;
        RECT 23.545 159.405 25.180 159.645 ;
        RECT 25.350 159.485 25.680 160.245 ;
        RECT 25.850 159.405 26.105 160.075 ;
        RECT 22.705 159.065 25.765 159.235 ;
        RECT 22.620 158.685 22.970 158.895 ;
        RECT 23.140 158.685 23.585 158.885 ;
        RECT 23.755 158.685 24.230 158.885 ;
        RECT 20.315 157.695 21.985 158.465 ;
        RECT 22.705 158.345 23.770 158.515 ;
        RECT 22.705 157.865 22.875 158.345 ;
        RECT 23.045 157.695 23.375 158.175 ;
        RECT 23.600 158.115 23.770 158.345 ;
        RECT 23.950 158.285 24.230 158.685 ;
        RECT 24.500 158.685 24.830 158.885 ;
        RECT 25.000 158.715 25.375 158.885 ;
        RECT 25.000 158.685 25.365 158.715 ;
        RECT 24.500 158.285 24.785 158.685 ;
        RECT 25.595 158.515 25.765 159.065 ;
        RECT 24.965 158.345 25.765 158.515 ;
        RECT 24.965 158.115 25.135 158.345 ;
        RECT 25.935 158.275 26.105 159.405 ;
        RECT 26.295 159.155 28.885 160.245 ;
        RECT 25.920 158.205 26.105 158.275 ;
        RECT 25.895 158.195 26.105 158.205 ;
        RECT 23.600 157.865 25.135 158.115 ;
        RECT 25.305 157.695 25.635 158.175 ;
        RECT 25.850 157.865 26.105 158.195 ;
        RECT 26.295 158.465 27.505 158.985 ;
        RECT 27.675 158.635 28.885 159.155 ;
        RECT 29.055 159.485 29.570 159.895 ;
        RECT 29.805 159.485 29.975 160.245 ;
        RECT 30.145 159.905 32.175 160.075 ;
        RECT 29.055 158.675 29.395 159.485 ;
        RECT 30.145 159.240 30.315 159.905 ;
        RECT 30.710 159.565 31.835 159.735 ;
        RECT 29.565 159.050 30.315 159.240 ;
        RECT 30.485 159.225 31.495 159.395 ;
        RECT 29.055 158.505 30.285 158.675 ;
        RECT 26.295 157.695 28.885 158.465 ;
        RECT 29.330 157.900 29.575 158.505 ;
        RECT 29.795 157.695 30.305 158.230 ;
        RECT 30.485 157.865 30.675 159.225 ;
        RECT 30.845 158.545 31.120 159.025 ;
        RECT 30.845 158.375 31.125 158.545 ;
        RECT 31.325 158.425 31.495 159.225 ;
        RECT 31.665 158.435 31.835 159.565 ;
        RECT 32.005 158.935 32.175 159.905 ;
        RECT 32.345 159.105 32.515 160.245 ;
        RECT 32.685 159.105 33.020 160.075 ;
        RECT 32.005 158.605 32.200 158.935 ;
        RECT 32.425 158.605 32.680 158.935 ;
        RECT 32.425 158.435 32.595 158.605 ;
        RECT 32.850 158.435 33.020 159.105 ;
        RECT 34.205 159.235 34.375 160.075 ;
        RECT 34.545 159.905 35.715 160.075 ;
        RECT 34.545 159.405 34.875 159.905 ;
        RECT 35.385 159.865 35.715 159.905 ;
        RECT 35.905 159.825 36.260 160.245 ;
        RECT 35.045 159.645 35.275 159.735 ;
        RECT 36.430 159.645 36.680 160.075 ;
        RECT 35.045 159.405 36.680 159.645 ;
        RECT 36.850 159.485 37.180 160.245 ;
        RECT 37.350 159.405 37.605 160.075 ;
        RECT 34.205 159.065 37.265 159.235 ;
        RECT 34.120 158.685 34.470 158.895 ;
        RECT 34.640 158.685 35.085 158.885 ;
        RECT 35.255 158.685 35.730 158.885 ;
        RECT 30.845 157.865 31.120 158.375 ;
        RECT 31.665 158.265 32.595 158.435 ;
        RECT 31.665 158.230 31.840 158.265 ;
        RECT 31.310 157.865 31.840 158.230 ;
        RECT 32.265 157.695 32.595 158.095 ;
        RECT 32.765 157.865 33.020 158.435 ;
        RECT 34.205 158.345 35.270 158.515 ;
        RECT 34.205 157.865 34.375 158.345 ;
        RECT 34.545 157.695 34.875 158.175 ;
        RECT 35.100 158.115 35.270 158.345 ;
        RECT 35.450 158.285 35.730 158.685 ;
        RECT 36.000 158.685 36.330 158.885 ;
        RECT 36.500 158.715 36.875 158.885 ;
        RECT 36.500 158.685 36.865 158.715 ;
        RECT 36.000 158.285 36.285 158.685 ;
        RECT 37.095 158.515 37.265 159.065 ;
        RECT 36.465 158.345 37.265 158.515 ;
        RECT 36.465 158.115 36.635 158.345 ;
        RECT 37.435 158.275 37.605 159.405 ;
        RECT 37.885 159.235 38.055 160.075 ;
        RECT 38.225 159.905 39.395 160.075 ;
        RECT 38.225 159.405 38.555 159.905 ;
        RECT 39.065 159.865 39.395 159.905 ;
        RECT 39.585 159.825 39.940 160.245 ;
        RECT 38.725 159.645 38.955 159.735 ;
        RECT 40.110 159.645 40.360 160.075 ;
        RECT 38.725 159.405 40.360 159.645 ;
        RECT 40.530 159.485 40.860 160.245 ;
        RECT 41.030 159.405 41.285 160.075 ;
        RECT 37.885 159.065 40.945 159.235 ;
        RECT 37.800 158.685 38.150 158.895 ;
        RECT 38.320 158.685 38.765 158.885 ;
        RECT 38.935 158.685 39.410 158.885 ;
        RECT 37.420 158.205 37.605 158.275 ;
        RECT 37.395 158.195 37.605 158.205 ;
        RECT 35.100 157.865 36.635 158.115 ;
        RECT 36.805 157.695 37.135 158.175 ;
        RECT 37.350 157.865 37.605 158.195 ;
        RECT 37.885 158.345 38.950 158.515 ;
        RECT 37.885 157.865 38.055 158.345 ;
        RECT 38.225 157.695 38.555 158.175 ;
        RECT 38.780 158.115 38.950 158.345 ;
        RECT 39.130 158.285 39.410 158.685 ;
        RECT 39.680 158.685 40.010 158.885 ;
        RECT 40.180 158.685 40.545 158.885 ;
        RECT 39.680 158.285 39.965 158.685 ;
        RECT 40.775 158.515 40.945 159.065 ;
        RECT 40.145 158.345 40.945 158.515 ;
        RECT 40.145 158.115 40.315 158.345 ;
        RECT 41.115 158.275 41.285 159.405 ;
        RECT 41.475 159.080 41.765 160.245 ;
        RECT 41.940 159.105 42.275 160.075 ;
        RECT 42.445 159.105 42.615 160.245 ;
        RECT 42.785 159.905 44.815 160.075 ;
        RECT 41.940 158.435 42.110 159.105 ;
        RECT 42.785 158.935 42.955 159.905 ;
        RECT 42.280 158.605 42.535 158.935 ;
        RECT 42.760 158.605 42.955 158.935 ;
        RECT 43.125 159.565 44.250 159.735 ;
        RECT 42.365 158.435 42.535 158.605 ;
        RECT 43.125 158.435 43.295 159.565 ;
        RECT 41.100 158.205 41.285 158.275 ;
        RECT 41.075 158.195 41.285 158.205 ;
        RECT 38.780 157.865 40.315 158.115 ;
        RECT 40.485 157.695 40.815 158.175 ;
        RECT 41.030 157.865 41.285 158.195 ;
        RECT 41.475 157.695 41.765 158.420 ;
        RECT 41.940 157.865 42.195 158.435 ;
        RECT 42.365 158.265 43.295 158.435 ;
        RECT 43.465 159.225 44.475 159.395 ;
        RECT 43.465 158.425 43.635 159.225 ;
        RECT 43.840 158.885 44.115 159.025 ;
        RECT 43.835 158.715 44.115 158.885 ;
        RECT 43.120 158.230 43.295 158.265 ;
        RECT 42.365 157.695 42.695 158.095 ;
        RECT 43.120 157.865 43.650 158.230 ;
        RECT 43.840 157.865 44.115 158.715 ;
        RECT 44.285 157.865 44.475 159.225 ;
        RECT 44.645 159.240 44.815 159.905 ;
        RECT 44.985 159.485 45.155 160.245 ;
        RECT 45.390 159.485 45.905 159.895 ;
        RECT 44.645 159.050 45.395 159.240 ;
        RECT 45.565 158.675 45.905 159.485 ;
        RECT 44.675 158.505 45.905 158.675 ;
        RECT 46.110 159.455 46.645 160.075 ;
        RECT 44.655 157.695 45.165 158.230 ;
        RECT 45.385 157.900 45.630 158.505 ;
        RECT 46.110 158.435 46.425 159.455 ;
        RECT 46.815 159.445 47.145 160.245 ;
        RECT 48.375 159.485 48.890 159.895 ;
        RECT 49.125 159.485 49.295 160.245 ;
        RECT 49.465 159.905 51.495 160.075 ;
        RECT 47.630 159.275 48.020 159.450 ;
        RECT 46.595 159.105 48.020 159.275 ;
        RECT 46.595 158.605 46.765 159.105 ;
        RECT 46.110 157.865 46.725 158.435 ;
        RECT 47.015 158.375 47.280 158.935 ;
        RECT 47.450 158.205 47.620 159.105 ;
        RECT 47.790 158.375 48.145 158.935 ;
        RECT 48.375 158.675 48.715 159.485 ;
        RECT 49.465 159.240 49.635 159.905 ;
        RECT 50.030 159.565 51.155 159.735 ;
        RECT 48.885 159.050 49.635 159.240 ;
        RECT 49.805 159.225 50.815 159.395 ;
        RECT 48.375 158.505 49.605 158.675 ;
        RECT 46.895 157.695 47.110 158.205 ;
        RECT 47.340 157.875 47.620 158.205 ;
        RECT 47.800 157.695 48.040 158.205 ;
        RECT 48.650 157.900 48.895 158.505 ;
        RECT 49.115 157.695 49.625 158.230 ;
        RECT 49.805 157.865 49.995 159.225 ;
        RECT 50.165 158.885 50.440 159.025 ;
        RECT 50.165 158.715 50.445 158.885 ;
        RECT 50.165 157.865 50.440 158.715 ;
        RECT 50.645 158.425 50.815 159.225 ;
        RECT 50.985 158.435 51.155 159.565 ;
        RECT 51.325 158.935 51.495 159.905 ;
        RECT 51.665 159.105 51.835 160.245 ;
        RECT 52.005 159.105 52.340 160.075 ;
        RECT 51.325 158.605 51.520 158.935 ;
        RECT 51.745 158.605 52.000 158.935 ;
        RECT 51.745 158.435 51.915 158.605 ;
        RECT 52.170 158.435 52.340 159.105 ;
        RECT 50.985 158.265 51.915 158.435 ;
        RECT 50.985 158.230 51.160 158.265 ;
        RECT 50.630 157.865 51.160 158.230 ;
        RECT 51.585 157.695 51.915 158.095 ;
        RECT 52.085 157.865 52.340 158.435 ;
        RECT 52.520 159.055 52.775 159.935 ;
        RECT 52.945 159.105 53.250 160.245 ;
        RECT 53.590 159.865 53.920 160.245 ;
        RECT 54.100 159.695 54.270 159.985 ;
        RECT 54.440 159.785 54.690 160.245 ;
        RECT 53.470 159.525 54.270 159.695 ;
        RECT 54.860 159.735 55.730 160.075 ;
        RECT 52.520 158.405 52.730 159.055 ;
        RECT 53.470 158.935 53.640 159.525 ;
        RECT 54.860 159.355 55.030 159.735 ;
        RECT 55.965 159.615 56.135 160.075 ;
        RECT 56.305 159.785 56.675 160.245 ;
        RECT 56.970 159.645 57.140 159.985 ;
        RECT 57.310 159.815 57.640 160.245 ;
        RECT 57.875 159.645 58.045 159.985 ;
        RECT 53.810 159.185 55.030 159.355 ;
        RECT 55.200 159.275 55.660 159.565 ;
        RECT 55.965 159.445 56.525 159.615 ;
        RECT 56.970 159.475 58.045 159.645 ;
        RECT 58.215 159.745 58.895 160.075 ;
        RECT 59.110 159.745 59.360 160.075 ;
        RECT 59.530 159.785 59.780 160.245 ;
        RECT 56.355 159.305 56.525 159.445 ;
        RECT 55.200 159.265 56.165 159.275 ;
        RECT 54.860 159.095 55.030 159.185 ;
        RECT 55.490 159.105 56.165 159.265 ;
        RECT 52.900 158.905 53.640 158.935 ;
        RECT 52.900 158.605 53.815 158.905 ;
        RECT 53.490 158.430 53.815 158.605 ;
        RECT 52.520 157.875 52.775 158.405 ;
        RECT 52.945 157.695 53.250 158.155 ;
        RECT 53.495 158.075 53.815 158.430 ;
        RECT 53.985 158.645 54.525 159.015 ;
        RECT 54.860 158.925 55.265 159.095 ;
        RECT 53.985 158.245 54.225 158.645 ;
        RECT 54.705 158.475 54.925 158.755 ;
        RECT 54.395 158.305 54.925 158.475 ;
        RECT 54.395 158.075 54.565 158.305 ;
        RECT 55.095 158.145 55.265 158.925 ;
        RECT 55.435 158.315 55.785 158.935 ;
        RECT 55.955 158.315 56.165 159.105 ;
        RECT 56.355 159.135 57.855 159.305 ;
        RECT 56.355 158.445 56.525 159.135 ;
        RECT 58.215 158.965 58.385 159.745 ;
        RECT 59.190 159.615 59.360 159.745 ;
        RECT 56.695 158.795 58.385 158.965 ;
        RECT 58.555 159.185 59.020 159.575 ;
        RECT 59.190 159.445 59.585 159.615 ;
        RECT 56.695 158.615 56.865 158.795 ;
        RECT 53.495 157.905 54.565 158.075 ;
        RECT 54.735 157.695 54.925 158.135 ;
        RECT 55.095 157.865 56.045 158.145 ;
        RECT 56.355 158.055 56.615 158.445 ;
        RECT 57.035 158.375 57.825 158.625 ;
        RECT 56.265 157.885 56.615 158.055 ;
        RECT 56.825 157.695 57.155 158.155 ;
        RECT 58.030 158.085 58.200 158.795 ;
        RECT 58.555 158.595 58.725 159.185 ;
        RECT 58.370 158.375 58.725 158.595 ;
        RECT 58.895 158.375 59.245 158.995 ;
        RECT 59.415 158.085 59.585 159.445 ;
        RECT 59.950 159.275 60.275 160.060 ;
        RECT 59.755 158.225 60.215 159.275 ;
        RECT 58.030 157.915 58.885 158.085 ;
        RECT 59.090 157.915 59.585 158.085 ;
        RECT 59.755 157.695 60.085 158.055 ;
        RECT 60.445 157.955 60.615 160.075 ;
        RECT 60.785 159.745 61.115 160.245 ;
        RECT 61.285 159.575 61.540 160.075 ;
        RECT 60.790 159.405 61.540 159.575 ;
        RECT 60.790 158.415 61.020 159.405 ;
        RECT 61.805 159.315 61.975 160.075 ;
        RECT 62.155 159.485 62.485 160.245 ;
        RECT 61.190 158.585 61.540 159.235 ;
        RECT 61.805 159.145 62.470 159.315 ;
        RECT 62.655 159.170 62.925 160.075 ;
        RECT 62.300 159.000 62.470 159.145 ;
        RECT 61.735 158.595 62.065 158.965 ;
        RECT 62.300 158.670 62.585 159.000 ;
        RECT 62.300 158.415 62.470 158.670 ;
        RECT 60.790 158.245 61.540 158.415 ;
        RECT 60.785 157.695 61.115 158.075 ;
        RECT 61.285 157.955 61.540 158.245 ;
        RECT 61.805 158.245 62.470 158.415 ;
        RECT 62.755 158.370 62.925 159.170 ;
        RECT 61.805 157.865 61.975 158.245 ;
        RECT 62.155 157.695 62.485 158.075 ;
        RECT 62.665 157.865 62.925 158.370 ;
        RECT 63.100 159.105 63.435 160.075 ;
        RECT 63.605 159.105 63.775 160.245 ;
        RECT 63.945 159.905 65.975 160.075 ;
        RECT 63.100 158.435 63.270 159.105 ;
        RECT 63.945 158.935 64.115 159.905 ;
        RECT 63.440 158.605 63.695 158.935 ;
        RECT 63.920 158.605 64.115 158.935 ;
        RECT 64.285 159.565 65.410 159.735 ;
        RECT 63.525 158.435 63.695 158.605 ;
        RECT 64.285 158.435 64.455 159.565 ;
        RECT 63.100 157.865 63.355 158.435 ;
        RECT 63.525 158.265 64.455 158.435 ;
        RECT 64.625 159.225 65.635 159.395 ;
        RECT 64.625 158.425 64.795 159.225 ;
        RECT 64.280 158.230 64.455 158.265 ;
        RECT 63.525 157.695 63.855 158.095 ;
        RECT 64.280 157.865 64.810 158.230 ;
        RECT 65.000 158.205 65.275 159.025 ;
        RECT 64.995 158.035 65.275 158.205 ;
        RECT 65.000 157.865 65.275 158.035 ;
        RECT 65.445 157.865 65.635 159.225 ;
        RECT 65.805 159.240 65.975 159.905 ;
        RECT 66.145 159.485 66.315 160.245 ;
        RECT 66.550 159.485 67.065 159.895 ;
        RECT 65.805 159.050 66.555 159.240 ;
        RECT 66.725 158.675 67.065 159.485 ;
        RECT 67.235 159.080 67.525 160.245 ;
        RECT 68.160 159.575 68.415 160.075 ;
        RECT 68.585 159.745 68.915 160.245 ;
        RECT 68.160 159.405 68.910 159.575 ;
        RECT 65.835 158.505 67.065 158.675 ;
        RECT 68.160 158.585 68.510 159.235 ;
        RECT 65.815 157.695 66.325 158.230 ;
        RECT 66.545 157.900 66.790 158.505 ;
        RECT 67.235 157.695 67.525 158.420 ;
        RECT 68.680 158.415 68.910 159.405 ;
        RECT 68.160 158.245 68.910 158.415 ;
        RECT 68.160 157.955 68.415 158.245 ;
        RECT 68.585 157.695 68.915 158.075 ;
        RECT 69.085 157.955 69.255 160.075 ;
        RECT 69.425 159.275 69.750 160.060 ;
        RECT 69.920 159.785 70.170 160.245 ;
        RECT 70.340 159.745 70.590 160.075 ;
        RECT 70.805 159.745 71.485 160.075 ;
        RECT 70.340 159.615 70.510 159.745 ;
        RECT 70.115 159.445 70.510 159.615 ;
        RECT 69.485 158.225 69.945 159.275 ;
        RECT 70.115 158.085 70.285 159.445 ;
        RECT 70.680 159.185 71.145 159.575 ;
        RECT 70.455 158.375 70.805 158.995 ;
        RECT 70.975 158.595 71.145 159.185 ;
        RECT 71.315 158.965 71.485 159.745 ;
        RECT 71.655 159.645 71.825 159.985 ;
        RECT 72.060 159.815 72.390 160.245 ;
        RECT 72.560 159.645 72.730 159.985 ;
        RECT 73.025 159.785 73.395 160.245 ;
        RECT 71.655 159.475 72.730 159.645 ;
        RECT 73.565 159.615 73.735 160.075 ;
        RECT 73.970 159.735 74.840 160.075 ;
        RECT 75.010 159.785 75.260 160.245 ;
        RECT 73.175 159.445 73.735 159.615 ;
        RECT 73.175 159.305 73.345 159.445 ;
        RECT 71.845 159.135 73.345 159.305 ;
        RECT 74.040 159.275 74.500 159.565 ;
        RECT 71.315 158.795 73.005 158.965 ;
        RECT 70.975 158.375 71.330 158.595 ;
        RECT 71.500 158.085 71.670 158.795 ;
        RECT 71.875 158.375 72.665 158.625 ;
        RECT 72.835 158.615 73.005 158.795 ;
        RECT 73.175 158.445 73.345 159.135 ;
        RECT 69.615 157.695 69.945 158.055 ;
        RECT 70.115 157.915 70.610 158.085 ;
        RECT 70.815 157.915 71.670 158.085 ;
        RECT 72.545 157.695 72.875 158.155 ;
        RECT 73.085 158.055 73.345 158.445 ;
        RECT 73.535 159.265 74.500 159.275 ;
        RECT 74.670 159.355 74.840 159.735 ;
        RECT 75.430 159.695 75.600 159.985 ;
        RECT 75.780 159.865 76.110 160.245 ;
        RECT 75.430 159.525 76.230 159.695 ;
        RECT 73.535 159.105 74.210 159.265 ;
        RECT 74.670 159.185 75.890 159.355 ;
        RECT 73.535 158.315 73.745 159.105 ;
        RECT 74.670 159.095 74.840 159.185 ;
        RECT 73.915 158.315 74.265 158.935 ;
        RECT 74.435 158.925 74.840 159.095 ;
        RECT 74.435 158.145 74.605 158.925 ;
        RECT 74.775 158.475 74.995 158.755 ;
        RECT 75.175 158.645 75.715 159.015 ;
        RECT 76.060 158.935 76.230 159.525 ;
        RECT 76.450 159.105 76.755 160.245 ;
        RECT 76.925 159.055 77.180 159.935 ;
        RECT 77.360 159.105 77.615 160.245 ;
        RECT 77.785 159.205 78.095 160.075 ;
        RECT 78.295 159.785 78.585 160.245 ;
        RECT 78.755 159.865 80.065 160.035 ;
        RECT 78.755 159.615 78.925 159.865 ;
        RECT 80.595 159.785 80.815 160.245 ;
        RECT 80.985 159.615 81.320 160.075 ;
        RECT 78.265 159.445 78.925 159.615 ;
        RECT 79.095 159.445 81.320 159.615 ;
        RECT 76.060 158.905 76.800 158.935 ;
        RECT 74.775 158.305 75.305 158.475 ;
        RECT 73.085 157.885 73.435 158.055 ;
        RECT 73.655 157.865 74.605 158.145 ;
        RECT 74.775 157.695 74.965 158.135 ;
        RECT 75.135 158.075 75.305 158.305 ;
        RECT 75.475 158.245 75.715 158.645 ;
        RECT 75.885 158.605 76.800 158.905 ;
        RECT 75.885 158.430 76.210 158.605 ;
        RECT 75.885 158.075 76.205 158.430 ;
        RECT 76.970 158.405 77.180 159.055 ;
        RECT 75.135 157.905 76.205 158.075 ;
        RECT 76.450 157.695 76.755 158.155 ;
        RECT 76.925 157.875 77.180 158.405 ;
        RECT 77.360 157.695 77.615 158.495 ;
        RECT 77.785 158.360 77.955 159.205 ;
        RECT 78.265 158.935 78.435 159.445 ;
        RECT 79.095 159.275 79.265 159.445 ;
        RECT 78.125 158.605 78.435 158.935 ;
        RECT 78.605 159.105 79.265 159.275 ;
        RECT 78.605 158.605 78.775 159.105 ;
        RECT 79.545 158.925 80.360 159.235 ;
        RECT 79.545 158.890 79.715 158.925 ;
        RECT 78.265 158.415 78.435 158.605 ;
        RECT 77.785 157.865 78.035 158.360 ;
        RECT 78.265 158.245 78.875 158.415 ;
        RECT 79.085 158.375 79.715 158.890 ;
        RECT 79.895 158.345 80.360 158.635 ;
        RECT 80.630 158.365 80.820 159.235 ;
        RECT 78.705 158.075 78.875 158.245 ;
        RECT 78.205 157.695 78.535 158.075 ;
        RECT 78.705 157.905 80.000 158.075 ;
        RECT 80.170 158.030 80.360 158.345 ;
        RECT 80.620 157.695 80.820 158.195 ;
        RECT 80.990 157.865 81.320 159.445 ;
        RECT 81.585 159.625 81.755 160.055 ;
        RECT 81.925 159.795 82.255 160.245 ;
        RECT 81.585 159.395 82.260 159.625 ;
        RECT 81.555 158.375 81.855 159.225 ;
        RECT 82.025 158.745 82.260 159.395 ;
        RECT 82.430 159.085 82.715 160.030 ;
        RECT 82.895 159.775 83.580 160.245 ;
        RECT 82.890 159.255 83.585 159.565 ;
        RECT 83.760 159.190 84.065 159.975 ;
        RECT 84.345 159.625 84.515 160.055 ;
        RECT 84.685 159.795 85.015 160.245 ;
        RECT 84.345 159.395 85.020 159.625 ;
        RECT 82.430 158.935 83.290 159.085 ;
        RECT 82.430 158.915 83.715 158.935 ;
        RECT 82.025 158.415 82.560 158.745 ;
        RECT 82.730 158.555 83.715 158.915 ;
        RECT 82.025 158.265 82.245 158.415 ;
        RECT 81.500 157.695 81.835 158.200 ;
        RECT 82.005 157.890 82.245 158.265 ;
        RECT 82.730 158.220 82.900 158.555 ;
        RECT 83.890 158.385 84.065 159.190 ;
        RECT 82.525 158.025 82.900 158.220 ;
        RECT 82.525 157.880 82.695 158.025 ;
        RECT 83.260 157.695 83.655 158.190 ;
        RECT 83.825 157.865 84.065 158.385 ;
        RECT 84.315 158.375 84.615 159.225 ;
        RECT 84.785 158.745 85.020 159.395 ;
        RECT 85.190 159.085 85.475 160.030 ;
        RECT 85.655 159.775 86.340 160.245 ;
        RECT 85.650 159.255 86.345 159.565 ;
        RECT 86.520 159.190 86.825 159.975 ;
        RECT 85.190 158.935 86.050 159.085 ;
        RECT 85.190 158.915 86.475 158.935 ;
        RECT 84.785 158.415 85.320 158.745 ;
        RECT 85.490 158.555 86.475 158.915 ;
        RECT 84.785 158.265 85.005 158.415 ;
        RECT 84.260 157.695 84.595 158.200 ;
        RECT 84.765 157.890 85.005 158.265 ;
        RECT 85.490 158.220 85.660 158.555 ;
        RECT 86.650 158.385 86.825 159.190 ;
        RECT 87.105 159.315 87.275 160.075 ;
        RECT 87.455 159.485 87.785 160.245 ;
        RECT 87.105 159.145 87.770 159.315 ;
        RECT 87.955 159.170 88.225 160.075 ;
        RECT 88.395 159.650 88.655 159.830 ;
        RECT 88.860 159.820 89.220 160.245 ;
        RECT 89.735 159.820 90.065 160.245 ;
        RECT 90.245 159.735 91.445 159.975 ;
        RECT 88.395 159.565 90.030 159.650 ;
        RECT 88.395 159.480 90.970 159.565 ;
        RECT 88.395 159.420 89.075 159.480 ;
        RECT 87.600 159.000 87.770 159.145 ;
        RECT 87.035 158.595 87.365 158.965 ;
        RECT 87.600 158.670 87.885 159.000 ;
        RECT 87.600 158.415 87.770 158.670 ;
        RECT 85.285 158.025 85.660 158.220 ;
        RECT 85.285 157.880 85.455 158.025 ;
        RECT 86.020 157.695 86.415 158.190 ;
        RECT 86.585 157.865 86.825 158.385 ;
        RECT 87.105 158.245 87.770 158.415 ;
        RECT 88.055 158.370 88.225 159.170 ;
        RECT 88.395 158.685 88.735 159.250 ;
        RECT 88.905 158.515 89.075 159.420 ;
        RECT 89.860 159.395 90.970 159.480 ;
        RECT 87.105 157.865 87.275 158.245 ;
        RECT 87.455 157.695 87.785 158.075 ;
        RECT 87.965 157.865 88.225 158.370 ;
        RECT 88.395 158.345 89.075 158.515 ;
        RECT 89.245 159.105 89.640 159.310 ;
        RECT 88.395 157.900 88.655 158.345 ;
        RECT 89.245 158.205 89.415 159.105 ;
        RECT 89.585 158.545 89.755 158.935 ;
        RECT 90.005 158.685 90.540 159.225 ;
        RECT 90.800 158.935 90.970 159.395 ;
        RECT 91.140 159.105 91.445 159.535 ;
        RECT 91.615 159.155 92.825 160.245 ;
        RECT 90.800 158.605 91.100 158.935 ;
        RECT 89.585 158.515 89.905 158.545 ;
        RECT 89.585 158.435 90.470 158.515 ;
        RECT 91.275 158.435 91.445 159.105 ;
        RECT 89.585 158.375 91.445 158.435 ;
        RECT 89.735 158.345 91.445 158.375 ;
        RECT 90.300 158.265 91.445 158.345 ;
        RECT 88.905 157.695 89.075 158.175 ;
        RECT 89.245 157.875 89.595 158.205 ;
        RECT 89.830 157.695 90.000 158.175 ;
        RECT 90.300 157.915 90.470 158.265 ;
        RECT 91.140 158.215 91.445 158.265 ;
        RECT 91.615 158.445 92.135 158.985 ;
        RECT 92.305 158.615 92.825 159.155 ;
        RECT 92.995 159.080 93.285 160.245 ;
        RECT 90.640 157.695 90.970 158.095 ;
        RECT 91.140 157.915 91.395 158.215 ;
        RECT 91.615 157.695 92.825 158.445 ;
        RECT 92.995 157.695 93.285 158.420 ;
        RECT 93.465 157.875 93.725 160.065 ;
        RECT 93.895 159.515 94.235 160.245 ;
        RECT 94.415 159.335 94.685 160.065 ;
        RECT 93.915 159.115 94.685 159.335 ;
        RECT 94.865 159.355 95.095 160.065 ;
        RECT 95.265 159.535 95.595 160.245 ;
        RECT 95.765 159.355 96.025 160.065 ;
        RECT 97.140 159.575 97.395 160.075 ;
        RECT 97.565 159.745 97.895 160.245 ;
        RECT 97.140 159.405 97.890 159.575 ;
        RECT 94.865 159.115 96.025 159.355 ;
        RECT 93.915 158.445 94.205 159.115 ;
        RECT 94.385 158.625 94.850 158.935 ;
        RECT 95.030 158.625 95.555 158.935 ;
        RECT 93.915 158.245 95.145 158.445 ;
        RECT 93.985 157.695 94.655 158.065 ;
        RECT 94.835 157.875 95.145 158.245 ;
        RECT 95.325 157.985 95.555 158.625 ;
        RECT 95.735 158.605 96.035 158.935 ;
        RECT 97.140 158.585 97.490 159.235 ;
        RECT 95.735 157.695 96.025 158.425 ;
        RECT 97.660 158.415 97.890 159.405 ;
        RECT 97.140 158.245 97.890 158.415 ;
        RECT 97.140 157.955 97.395 158.245 ;
        RECT 97.565 157.695 97.895 158.075 ;
        RECT 98.065 157.955 98.235 160.075 ;
        RECT 98.405 159.275 98.730 160.060 ;
        RECT 98.900 159.785 99.150 160.245 ;
        RECT 99.320 159.745 99.570 160.075 ;
        RECT 99.785 159.745 100.465 160.075 ;
        RECT 99.320 159.615 99.490 159.745 ;
        RECT 99.095 159.445 99.490 159.615 ;
        RECT 98.465 158.225 98.925 159.275 ;
        RECT 99.095 158.085 99.265 159.445 ;
        RECT 99.660 159.185 100.125 159.575 ;
        RECT 99.435 158.375 99.785 158.995 ;
        RECT 99.955 158.595 100.125 159.185 ;
        RECT 100.295 158.965 100.465 159.745 ;
        RECT 100.635 159.645 100.805 159.985 ;
        RECT 101.040 159.815 101.370 160.245 ;
        RECT 101.540 159.645 101.710 159.985 ;
        RECT 102.005 159.785 102.375 160.245 ;
        RECT 100.635 159.475 101.710 159.645 ;
        RECT 102.545 159.615 102.715 160.075 ;
        RECT 102.950 159.735 103.820 160.075 ;
        RECT 103.990 159.785 104.240 160.245 ;
        RECT 102.155 159.445 102.715 159.615 ;
        RECT 102.155 159.305 102.325 159.445 ;
        RECT 100.825 159.135 102.325 159.305 ;
        RECT 103.020 159.275 103.480 159.565 ;
        RECT 100.295 158.795 101.985 158.965 ;
        RECT 99.955 158.375 100.310 158.595 ;
        RECT 100.480 158.085 100.650 158.795 ;
        RECT 100.855 158.375 101.645 158.625 ;
        RECT 101.815 158.615 101.985 158.795 ;
        RECT 102.155 158.445 102.325 159.135 ;
        RECT 98.595 157.695 98.925 158.055 ;
        RECT 99.095 157.915 99.590 158.085 ;
        RECT 99.795 157.915 100.650 158.085 ;
        RECT 101.525 157.695 101.855 158.155 ;
        RECT 102.065 158.055 102.325 158.445 ;
        RECT 102.515 159.265 103.480 159.275 ;
        RECT 103.650 159.355 103.820 159.735 ;
        RECT 104.410 159.695 104.580 159.985 ;
        RECT 104.760 159.865 105.090 160.245 ;
        RECT 104.410 159.525 105.210 159.695 ;
        RECT 102.515 159.105 103.190 159.265 ;
        RECT 103.650 159.185 104.870 159.355 ;
        RECT 102.515 158.315 102.725 159.105 ;
        RECT 103.650 159.095 103.820 159.185 ;
        RECT 102.895 158.315 103.245 158.935 ;
        RECT 103.415 158.925 103.820 159.095 ;
        RECT 103.415 158.145 103.585 158.925 ;
        RECT 103.755 158.475 103.975 158.755 ;
        RECT 104.155 158.645 104.695 159.015 ;
        RECT 105.040 158.935 105.210 159.525 ;
        RECT 105.430 159.105 105.735 160.245 ;
        RECT 105.905 159.055 106.160 159.935 ;
        RECT 106.340 159.105 106.595 160.245 ;
        RECT 106.790 159.695 107.985 160.025 ;
        RECT 105.040 158.905 105.780 158.935 ;
        RECT 103.755 158.305 104.285 158.475 ;
        RECT 102.065 157.885 102.415 158.055 ;
        RECT 102.635 157.865 103.585 158.145 ;
        RECT 103.755 157.695 103.945 158.135 ;
        RECT 104.115 158.075 104.285 158.305 ;
        RECT 104.455 158.245 104.695 158.645 ;
        RECT 104.865 158.605 105.780 158.905 ;
        RECT 104.865 158.430 105.190 158.605 ;
        RECT 104.865 158.075 105.185 158.430 ;
        RECT 105.950 158.405 106.160 159.055 ;
        RECT 106.845 158.935 107.015 159.495 ;
        RECT 107.240 159.275 107.660 159.525 ;
        RECT 108.165 159.445 108.445 160.245 ;
        RECT 107.240 159.105 108.485 159.275 ;
        RECT 108.655 159.105 108.925 160.075 ;
        RECT 109.565 159.435 109.860 160.245 ;
        RECT 108.315 158.935 108.485 159.105 ;
        RECT 106.340 158.685 106.675 158.935 ;
        RECT 106.845 158.605 107.585 158.935 ;
        RECT 108.315 158.605 108.545 158.935 ;
        RECT 106.845 158.515 107.095 158.605 ;
        RECT 104.115 157.905 105.185 158.075 ;
        RECT 105.430 157.695 105.735 158.155 ;
        RECT 105.905 157.875 106.160 158.405 ;
        RECT 106.360 158.345 107.095 158.515 ;
        RECT 108.315 158.435 108.485 158.605 ;
        RECT 106.360 157.875 106.670 158.345 ;
        RECT 107.745 158.265 108.485 158.435 ;
        RECT 108.755 158.370 108.925 159.105 ;
        RECT 110.040 158.935 110.285 160.075 ;
        RECT 110.460 159.435 110.720 160.245 ;
        RECT 111.320 160.240 117.595 160.245 ;
        RECT 110.900 158.935 111.150 160.070 ;
        RECT 111.320 159.445 111.580 160.240 ;
        RECT 111.750 159.345 112.010 160.070 ;
        RECT 112.180 159.515 112.440 160.240 ;
        RECT 112.610 159.345 112.870 160.070 ;
        RECT 113.040 159.515 113.300 160.240 ;
        RECT 113.470 159.345 113.730 160.070 ;
        RECT 113.900 159.515 114.160 160.240 ;
        RECT 114.330 159.345 114.590 160.070 ;
        RECT 114.760 159.515 115.005 160.240 ;
        RECT 115.175 159.345 115.435 160.070 ;
        RECT 115.620 159.515 115.865 160.240 ;
        RECT 116.035 159.345 116.295 160.070 ;
        RECT 116.480 159.515 116.725 160.240 ;
        RECT 116.895 159.345 117.155 160.070 ;
        RECT 117.340 159.515 117.595 160.240 ;
        RECT 111.750 159.330 117.155 159.345 ;
        RECT 117.765 159.330 118.055 160.070 ;
        RECT 118.225 159.500 118.495 160.245 ;
        RECT 111.750 159.105 118.495 159.330 ;
        RECT 109.555 158.375 109.870 158.935 ;
        RECT 110.040 158.685 117.160 158.935 ;
        RECT 106.840 157.695 107.575 158.175 ;
        RECT 107.745 157.915 107.915 158.265 ;
        RECT 108.085 157.695 108.465 158.095 ;
        RECT 108.655 158.025 108.925 158.370 ;
        RECT 109.555 157.695 109.860 158.205 ;
        RECT 110.040 157.875 110.290 158.685 ;
        RECT 110.460 157.695 110.720 158.220 ;
        RECT 110.900 157.875 111.150 158.685 ;
        RECT 117.330 158.515 118.495 159.105 ;
        RECT 118.755 159.080 119.045 160.245 ;
        RECT 119.220 159.105 119.555 160.075 ;
        RECT 119.725 159.105 119.895 160.245 ;
        RECT 120.065 159.905 122.095 160.075 ;
        RECT 111.750 158.345 118.495 158.515 ;
        RECT 119.220 158.435 119.390 159.105 ;
        RECT 120.065 158.935 120.235 159.905 ;
        RECT 119.560 158.605 119.815 158.935 ;
        RECT 120.040 158.605 120.235 158.935 ;
        RECT 120.405 159.565 121.530 159.735 ;
        RECT 119.645 158.435 119.815 158.605 ;
        RECT 120.405 158.435 120.575 159.565 ;
        RECT 111.320 157.695 111.580 158.255 ;
        RECT 111.750 157.890 112.010 158.345 ;
        RECT 112.180 157.695 112.440 158.175 ;
        RECT 112.610 157.890 112.870 158.345 ;
        RECT 113.040 157.695 113.300 158.175 ;
        RECT 113.470 157.890 113.730 158.345 ;
        RECT 113.900 157.695 114.145 158.175 ;
        RECT 114.315 157.890 114.590 158.345 ;
        RECT 114.760 157.695 115.005 158.175 ;
        RECT 115.175 157.890 115.435 158.345 ;
        RECT 115.615 157.695 115.865 158.175 ;
        RECT 116.035 157.890 116.295 158.345 ;
        RECT 116.475 157.695 116.725 158.175 ;
        RECT 116.895 157.890 117.155 158.345 ;
        RECT 117.335 157.695 117.595 158.175 ;
        RECT 117.765 157.890 118.025 158.345 ;
        RECT 118.195 157.695 118.495 158.175 ;
        RECT 118.755 157.695 119.045 158.420 ;
        RECT 119.220 157.865 119.475 158.435 ;
        RECT 119.645 158.265 120.575 158.435 ;
        RECT 120.745 159.225 121.755 159.395 ;
        RECT 120.745 158.425 120.915 159.225 ;
        RECT 121.120 158.885 121.395 159.025 ;
        RECT 121.115 158.715 121.395 158.885 ;
        RECT 120.400 158.230 120.575 158.265 ;
        RECT 119.645 157.695 119.975 158.095 ;
        RECT 120.400 157.865 120.930 158.230 ;
        RECT 121.120 157.865 121.395 158.715 ;
        RECT 121.565 157.865 121.755 159.225 ;
        RECT 121.925 159.240 122.095 159.905 ;
        RECT 122.265 159.485 122.435 160.245 ;
        RECT 122.670 159.485 123.185 159.895 ;
        RECT 121.925 159.050 122.675 159.240 ;
        RECT 122.845 158.675 123.185 159.485 ;
        RECT 123.365 159.265 123.695 160.075 ;
        RECT 123.865 159.445 124.105 160.245 ;
        RECT 123.365 159.095 124.080 159.265 ;
        RECT 123.360 158.685 123.740 158.925 ;
        RECT 123.910 158.855 124.080 159.095 ;
        RECT 124.285 159.225 124.455 160.075 ;
        RECT 124.625 159.445 124.955 160.245 ;
        RECT 125.125 159.225 125.295 160.075 ;
        RECT 124.285 159.055 125.295 159.225 ;
        RECT 125.465 159.095 125.795 160.245 ;
        RECT 126.300 159.275 126.690 159.450 ;
        RECT 127.175 159.445 127.505 160.245 ;
        RECT 127.675 159.455 128.210 160.075 ;
        RECT 126.300 159.105 127.725 159.275 ;
        RECT 123.910 158.685 124.410 158.855 ;
        RECT 121.955 158.505 123.185 158.675 ;
        RECT 123.910 158.515 124.080 158.685 ;
        RECT 124.800 158.545 125.295 159.055 ;
        RECT 124.795 158.515 125.295 158.545 ;
        RECT 121.935 157.695 122.445 158.230 ;
        RECT 122.665 157.900 122.910 158.505 ;
        RECT 123.445 158.345 124.080 158.515 ;
        RECT 124.285 158.345 125.295 158.515 ;
        RECT 123.445 157.865 123.615 158.345 ;
        RECT 123.795 157.695 124.035 158.175 ;
        RECT 124.285 157.865 124.455 158.345 ;
        RECT 124.625 157.695 124.955 158.175 ;
        RECT 125.125 157.865 125.295 158.345 ;
        RECT 125.465 157.695 125.795 158.495 ;
        RECT 126.175 158.375 126.530 158.935 ;
        RECT 126.700 158.205 126.870 159.105 ;
        RECT 127.040 158.375 127.305 158.935 ;
        RECT 127.555 158.605 127.725 159.105 ;
        RECT 127.895 158.435 128.210 159.455 ;
        RECT 128.455 159.105 128.685 160.245 ;
        RECT 128.855 159.095 129.185 160.075 ;
        RECT 129.355 159.105 129.565 160.245 ;
        RECT 129.795 159.170 130.065 160.075 ;
        RECT 130.235 159.485 130.565 160.245 ;
        RECT 130.745 159.315 130.915 160.075 ;
        RECT 128.435 158.685 128.765 158.935 ;
        RECT 126.280 157.695 126.520 158.205 ;
        RECT 126.700 157.875 126.980 158.205 ;
        RECT 127.210 157.695 127.425 158.205 ;
        RECT 127.595 157.865 128.210 158.435 ;
        RECT 128.455 157.695 128.685 158.515 ;
        RECT 128.935 158.495 129.185 159.095 ;
        RECT 128.855 157.865 129.185 158.495 ;
        RECT 129.355 157.695 129.565 158.515 ;
        RECT 129.795 158.370 129.965 159.170 ;
        RECT 130.250 159.145 130.915 159.315 ;
        RECT 130.250 159.000 130.420 159.145 ;
        RECT 130.135 158.670 130.420 159.000 ;
        RECT 132.100 159.105 132.435 160.075 ;
        RECT 132.605 159.105 132.775 160.245 ;
        RECT 132.945 159.905 134.975 160.075 ;
        RECT 130.250 158.415 130.420 158.670 ;
        RECT 130.655 158.595 130.985 158.965 ;
        RECT 132.100 158.435 132.270 159.105 ;
        RECT 132.945 158.935 133.115 159.905 ;
        RECT 132.440 158.605 132.695 158.935 ;
        RECT 132.920 158.605 133.115 158.935 ;
        RECT 133.285 159.565 134.410 159.735 ;
        RECT 132.525 158.435 132.695 158.605 ;
        RECT 133.285 158.435 133.455 159.565 ;
        RECT 129.795 157.865 130.055 158.370 ;
        RECT 130.250 158.245 130.915 158.415 ;
        RECT 130.235 157.695 130.565 158.075 ;
        RECT 130.745 157.865 130.915 158.245 ;
        RECT 132.100 157.865 132.355 158.435 ;
        RECT 132.525 158.265 133.455 158.435 ;
        RECT 133.625 159.225 134.635 159.395 ;
        RECT 133.625 158.425 133.795 159.225 ;
        RECT 133.280 158.230 133.455 158.265 ;
        RECT 132.525 157.695 132.855 158.095 ;
        RECT 133.280 157.865 133.810 158.230 ;
        RECT 134.000 158.205 134.275 159.025 ;
        RECT 133.995 158.035 134.275 158.205 ;
        RECT 134.000 157.865 134.275 158.035 ;
        RECT 134.445 157.865 134.635 159.225 ;
        RECT 134.805 159.240 134.975 159.905 ;
        RECT 135.145 159.485 135.315 160.245 ;
        RECT 135.550 159.485 136.065 159.895 ;
        RECT 134.805 159.050 135.555 159.240 ;
        RECT 135.725 158.675 136.065 159.485 ;
        RECT 134.835 158.505 136.065 158.675 ;
        RECT 137.160 159.105 137.495 160.075 ;
        RECT 137.665 159.105 137.835 160.245 ;
        RECT 138.005 159.905 140.035 160.075 ;
        RECT 134.815 157.695 135.325 158.230 ;
        RECT 135.545 157.900 135.790 158.505 ;
        RECT 137.160 158.435 137.330 159.105 ;
        RECT 138.005 158.935 138.175 159.905 ;
        RECT 137.500 158.605 137.755 158.935 ;
        RECT 137.980 158.605 138.175 158.935 ;
        RECT 138.345 159.565 139.470 159.735 ;
        RECT 137.585 158.435 137.755 158.605 ;
        RECT 138.345 158.435 138.515 159.565 ;
        RECT 137.160 157.865 137.415 158.435 ;
        RECT 137.585 158.265 138.515 158.435 ;
        RECT 138.685 159.225 139.695 159.395 ;
        RECT 138.685 158.425 138.855 159.225 ;
        RECT 138.340 158.230 138.515 158.265 ;
        RECT 137.585 157.695 137.915 158.095 ;
        RECT 138.340 157.865 138.870 158.230 ;
        RECT 139.060 158.205 139.335 159.025 ;
        RECT 139.055 158.035 139.335 158.205 ;
        RECT 139.060 157.865 139.335 158.035 ;
        RECT 139.505 157.865 139.695 159.225 ;
        RECT 139.865 159.240 140.035 159.905 ;
        RECT 140.205 159.485 140.375 160.245 ;
        RECT 140.610 159.485 141.125 159.895 ;
        RECT 139.865 159.050 140.615 159.240 ;
        RECT 140.785 158.675 141.125 159.485 ;
        RECT 141.295 159.155 143.885 160.245 ;
        RECT 139.895 158.505 141.125 158.675 ;
        RECT 139.875 157.695 140.385 158.230 ;
        RECT 140.605 157.900 140.850 158.505 ;
        RECT 141.295 158.465 142.505 158.985 ;
        RECT 142.675 158.635 143.885 159.155 ;
        RECT 144.515 159.080 144.805 160.245 ;
        RECT 144.975 159.810 150.320 160.245 ;
        RECT 150.495 159.810 155.840 160.245 ;
        RECT 141.295 157.695 143.885 158.465 ;
        RECT 144.515 157.695 144.805 158.420 ;
        RECT 146.560 158.240 146.900 159.070 ;
        RECT 148.380 158.560 148.730 159.810 ;
        RECT 152.080 158.240 152.420 159.070 ;
        RECT 153.900 158.560 154.250 159.810 ;
        RECT 156.935 159.155 158.145 160.245 ;
        RECT 156.935 158.615 157.455 159.155 ;
        RECT 157.625 158.445 158.145 158.985 ;
        RECT 144.975 157.695 150.320 158.240 ;
        RECT 150.495 157.695 155.840 158.240 ;
        RECT 156.935 157.695 158.145 158.445 ;
        RECT 2.750 157.525 158.230 157.695 ;
        RECT 2.835 156.775 4.045 157.525 ;
        RECT 2.835 156.235 3.355 156.775 ;
        RECT 4.215 156.755 5.885 157.525 ;
        RECT 3.525 156.065 4.045 156.605 ;
        RECT 4.215 156.235 4.965 156.755 ;
        RECT 6.790 156.715 7.035 157.320 ;
        RECT 7.255 156.990 7.765 157.525 ;
        RECT 5.135 156.065 5.885 156.585 ;
        RECT 2.835 154.975 4.045 156.065 ;
        RECT 4.215 154.975 5.885 156.065 ;
        RECT 6.515 156.545 7.745 156.715 ;
        RECT 6.515 155.735 6.855 156.545 ;
        RECT 7.025 155.980 7.775 156.170 ;
        RECT 6.515 155.325 7.030 155.735 ;
        RECT 7.265 154.975 7.435 155.735 ;
        RECT 7.605 155.315 7.775 155.980 ;
        RECT 7.945 155.995 8.135 157.355 ;
        RECT 8.305 156.505 8.580 157.355 ;
        RECT 8.770 156.990 9.300 157.355 ;
        RECT 9.725 157.125 10.055 157.525 ;
        RECT 9.125 156.955 9.300 156.990 ;
        RECT 8.305 156.335 8.585 156.505 ;
        RECT 8.305 156.195 8.580 156.335 ;
        RECT 8.785 155.995 8.955 156.795 ;
        RECT 7.945 155.825 8.955 155.995 ;
        RECT 9.125 156.785 10.055 156.955 ;
        RECT 10.225 156.785 10.480 157.355 ;
        RECT 10.660 156.975 10.915 157.265 ;
        RECT 11.085 157.145 11.415 157.525 ;
        RECT 10.660 156.805 11.410 156.975 ;
        RECT 9.125 155.655 9.295 156.785 ;
        RECT 9.885 156.615 10.055 156.785 ;
        RECT 8.170 155.485 9.295 155.655 ;
        RECT 9.465 156.285 9.660 156.615 ;
        RECT 9.885 156.285 10.140 156.615 ;
        RECT 9.465 155.315 9.635 156.285 ;
        RECT 10.310 156.115 10.480 156.785 ;
        RECT 7.605 155.145 9.635 155.315 ;
        RECT 9.805 154.975 9.975 156.115 ;
        RECT 10.145 155.145 10.480 156.115 ;
        RECT 10.660 155.985 11.010 156.635 ;
        RECT 11.180 155.815 11.410 156.805 ;
        RECT 10.660 155.645 11.410 155.815 ;
        RECT 10.660 155.145 10.915 155.645 ;
        RECT 11.085 154.975 11.415 155.475 ;
        RECT 11.585 155.145 11.755 157.265 ;
        RECT 12.115 157.165 12.445 157.525 ;
        RECT 12.615 157.135 13.110 157.305 ;
        RECT 13.315 157.135 14.170 157.305 ;
        RECT 11.985 155.945 12.445 156.995 ;
        RECT 11.925 155.160 12.250 155.945 ;
        RECT 12.615 155.775 12.785 157.135 ;
        RECT 12.955 156.225 13.305 156.845 ;
        RECT 13.475 156.625 13.830 156.845 ;
        RECT 13.475 156.035 13.645 156.625 ;
        RECT 14.000 156.425 14.170 157.135 ;
        RECT 15.045 157.065 15.375 157.525 ;
        RECT 15.585 157.165 15.935 157.335 ;
        RECT 14.375 156.595 15.165 156.845 ;
        RECT 15.585 156.775 15.845 157.165 ;
        RECT 16.155 157.075 17.105 157.355 ;
        RECT 17.275 157.085 17.465 157.525 ;
        RECT 17.635 157.145 18.705 157.315 ;
        RECT 15.335 156.425 15.505 156.605 ;
        RECT 12.615 155.605 13.010 155.775 ;
        RECT 13.180 155.645 13.645 156.035 ;
        RECT 13.815 156.255 15.505 156.425 ;
        RECT 12.840 155.475 13.010 155.605 ;
        RECT 13.815 155.475 13.985 156.255 ;
        RECT 15.675 156.085 15.845 156.775 ;
        RECT 14.345 155.915 15.845 156.085 ;
        RECT 16.035 156.115 16.245 156.905 ;
        RECT 16.415 156.285 16.765 156.905 ;
        RECT 16.935 156.295 17.105 157.075 ;
        RECT 17.635 156.915 17.805 157.145 ;
        RECT 17.275 156.745 17.805 156.915 ;
        RECT 17.275 156.465 17.495 156.745 ;
        RECT 17.975 156.575 18.215 156.975 ;
        RECT 16.935 156.125 17.340 156.295 ;
        RECT 17.675 156.205 18.215 156.575 ;
        RECT 18.385 156.790 18.705 157.145 ;
        RECT 18.950 157.065 19.255 157.525 ;
        RECT 19.425 156.815 19.680 157.345 ;
        RECT 18.385 156.615 18.710 156.790 ;
        RECT 18.385 156.315 19.300 156.615 ;
        RECT 18.560 156.285 19.300 156.315 ;
        RECT 16.035 155.955 16.710 156.115 ;
        RECT 17.170 156.035 17.340 156.125 ;
        RECT 16.035 155.945 17.000 155.955 ;
        RECT 15.675 155.775 15.845 155.915 ;
        RECT 12.420 154.975 12.670 155.435 ;
        RECT 12.840 155.145 13.090 155.475 ;
        RECT 13.305 155.145 13.985 155.475 ;
        RECT 14.155 155.575 15.230 155.745 ;
        RECT 15.675 155.605 16.235 155.775 ;
        RECT 16.540 155.655 17.000 155.945 ;
        RECT 17.170 155.865 18.390 156.035 ;
        RECT 14.155 155.235 14.325 155.575 ;
        RECT 14.560 154.975 14.890 155.405 ;
        RECT 15.060 155.235 15.230 155.575 ;
        RECT 15.525 154.975 15.895 155.435 ;
        RECT 16.065 155.145 16.235 155.605 ;
        RECT 17.170 155.485 17.340 155.865 ;
        RECT 18.560 155.695 18.730 156.285 ;
        RECT 19.470 156.165 19.680 156.815 ;
        RECT 16.470 155.145 17.340 155.485 ;
        RECT 17.930 155.525 18.730 155.695 ;
        RECT 17.510 154.975 17.760 155.435 ;
        RECT 17.930 155.235 18.100 155.525 ;
        RECT 18.280 154.975 18.610 155.355 ;
        RECT 18.950 154.975 19.255 156.115 ;
        RECT 19.425 155.285 19.680 156.165 ;
        RECT 19.855 156.785 20.240 157.355 ;
        RECT 20.410 157.065 20.735 157.525 ;
        RECT 21.255 156.895 21.535 157.355 ;
        RECT 19.855 156.115 20.135 156.785 ;
        RECT 20.410 156.725 21.535 156.895 ;
        RECT 20.410 156.615 20.860 156.725 ;
        RECT 20.305 156.285 20.860 156.615 ;
        RECT 21.725 156.555 22.125 157.355 ;
        RECT 22.525 157.065 22.795 157.525 ;
        RECT 22.965 156.895 23.250 157.355 ;
        RECT 19.855 155.145 20.240 156.115 ;
        RECT 20.410 155.825 20.860 156.285 ;
        RECT 21.030 155.995 22.125 156.555 ;
        RECT 20.410 155.605 21.535 155.825 ;
        RECT 20.410 154.975 20.735 155.435 ;
        RECT 21.255 155.145 21.535 155.605 ;
        RECT 21.725 155.145 22.125 155.995 ;
        RECT 22.295 156.725 23.250 156.895 ;
        RECT 23.535 157.025 23.795 157.355 ;
        RECT 23.965 157.165 24.295 157.525 ;
        RECT 24.550 157.145 25.850 157.355 ;
        RECT 23.535 157.015 23.765 157.025 ;
        RECT 22.295 155.825 22.505 156.725 ;
        RECT 22.675 155.995 23.365 156.555 ;
        RECT 23.535 155.825 23.705 157.015 ;
        RECT 24.550 156.995 24.720 157.145 ;
        RECT 23.965 156.870 24.720 156.995 ;
        RECT 23.875 156.825 24.720 156.870 ;
        RECT 23.875 156.705 24.145 156.825 ;
        RECT 23.875 156.130 24.045 156.705 ;
        RECT 24.275 156.265 24.685 156.570 ;
        RECT 24.975 156.535 25.185 156.935 ;
        RECT 24.855 156.325 25.185 156.535 ;
        RECT 25.430 156.535 25.650 156.935 ;
        RECT 26.125 156.760 26.580 157.525 ;
        RECT 26.755 156.850 27.015 157.355 ;
        RECT 27.195 157.145 27.525 157.525 ;
        RECT 27.705 156.975 27.875 157.355 ;
        RECT 25.430 156.325 25.905 156.535 ;
        RECT 26.095 156.335 26.585 156.535 ;
        RECT 23.875 156.095 24.075 156.130 ;
        RECT 25.405 156.095 26.580 156.155 ;
        RECT 23.875 155.985 26.580 156.095 ;
        RECT 23.935 155.925 25.735 155.985 ;
        RECT 25.405 155.895 25.735 155.925 ;
        RECT 22.295 155.605 23.250 155.825 ;
        RECT 22.525 154.975 22.795 155.435 ;
        RECT 22.965 155.145 23.250 155.605 ;
        RECT 23.535 155.145 23.795 155.825 ;
        RECT 23.965 154.975 24.215 155.755 ;
        RECT 24.465 155.725 25.300 155.735 ;
        RECT 25.890 155.725 26.075 155.815 ;
        RECT 24.465 155.525 26.075 155.725 ;
        RECT 24.465 155.145 24.715 155.525 ;
        RECT 25.845 155.485 26.075 155.525 ;
        RECT 26.325 155.365 26.580 155.985 ;
        RECT 24.885 154.975 25.240 155.355 ;
        RECT 26.245 155.145 26.580 155.365 ;
        RECT 26.755 156.050 26.925 156.850 ;
        RECT 27.210 156.805 27.875 156.975 ;
        RECT 27.210 156.550 27.380 156.805 ;
        RECT 28.595 156.800 28.885 157.525 ;
        RECT 29.060 156.785 29.315 157.355 ;
        RECT 29.485 157.125 29.815 157.525 ;
        RECT 30.240 156.990 30.770 157.355 ;
        RECT 30.240 156.955 30.415 156.990 ;
        RECT 29.485 156.785 30.415 156.955 ;
        RECT 30.960 156.845 31.235 157.355 ;
        RECT 27.095 156.220 27.380 156.550 ;
        RECT 27.615 156.255 27.945 156.625 ;
        RECT 27.210 156.075 27.380 156.220 ;
        RECT 26.755 155.145 27.025 156.050 ;
        RECT 27.210 155.905 27.875 156.075 ;
        RECT 27.195 154.975 27.525 155.735 ;
        RECT 27.705 155.145 27.875 155.905 ;
        RECT 28.595 154.975 28.885 156.140 ;
        RECT 29.060 156.115 29.230 156.785 ;
        RECT 29.485 156.615 29.655 156.785 ;
        RECT 29.400 156.285 29.655 156.615 ;
        RECT 29.880 156.285 30.075 156.615 ;
        RECT 29.060 155.145 29.395 156.115 ;
        RECT 29.565 154.975 29.735 156.115 ;
        RECT 29.905 155.315 30.075 156.285 ;
        RECT 30.245 155.655 30.415 156.785 ;
        RECT 30.585 155.995 30.755 156.795 ;
        RECT 30.955 156.675 31.235 156.845 ;
        RECT 30.960 156.195 31.235 156.675 ;
        RECT 31.405 155.995 31.595 157.355 ;
        RECT 31.775 156.990 32.285 157.525 ;
        RECT 32.505 156.715 32.750 157.320 ;
        RECT 34.205 156.875 34.375 157.355 ;
        RECT 34.545 157.045 34.875 157.525 ;
        RECT 35.100 157.105 36.635 157.355 ;
        RECT 35.100 156.875 35.270 157.105 ;
        RECT 31.795 156.545 33.025 156.715 ;
        RECT 34.205 156.705 35.270 156.875 ;
        RECT 30.585 155.825 31.595 155.995 ;
        RECT 31.765 155.980 32.515 156.170 ;
        RECT 30.245 155.485 31.370 155.655 ;
        RECT 31.765 155.315 31.935 155.980 ;
        RECT 32.685 155.735 33.025 156.545 ;
        RECT 35.450 156.535 35.730 156.935 ;
        RECT 34.120 156.325 34.470 156.535 ;
        RECT 34.640 156.335 35.085 156.535 ;
        RECT 35.255 156.335 35.730 156.535 ;
        RECT 36.000 156.535 36.285 156.935 ;
        RECT 36.465 156.875 36.635 157.105 ;
        RECT 36.805 157.045 37.135 157.525 ;
        RECT 37.350 157.025 37.605 157.355 ;
        RECT 37.420 156.945 37.605 157.025 ;
        RECT 36.465 156.705 37.265 156.875 ;
        RECT 36.000 156.335 36.330 156.535 ;
        RECT 36.500 156.335 36.865 156.535 ;
        RECT 37.095 156.155 37.265 156.705 ;
        RECT 29.905 155.145 31.935 155.315 ;
        RECT 32.105 154.975 32.275 155.735 ;
        RECT 32.510 155.325 33.025 155.735 ;
        RECT 34.205 155.985 37.265 156.155 ;
        RECT 34.205 155.145 34.375 155.985 ;
        RECT 37.435 155.815 37.605 156.945 ;
        RECT 37.795 156.715 38.075 157.525 ;
        RECT 38.245 156.885 38.575 157.355 ;
        RECT 38.745 157.055 38.915 157.525 ;
        RECT 39.085 156.885 39.415 157.355 ;
        RECT 38.245 156.715 39.415 156.885 ;
        RECT 39.585 156.715 39.755 157.525 ;
        RECT 40.105 156.885 40.275 157.165 ;
        RECT 39.925 156.715 40.275 156.885 ;
        RECT 40.485 156.765 40.740 157.525 ;
        RECT 41.475 157.025 41.775 157.355 ;
        RECT 41.945 157.045 42.220 157.525 ;
        RECT 38.775 156.675 38.945 156.715 ;
        RECT 38.190 156.335 38.630 156.545 ;
        RECT 34.545 155.315 34.875 155.815 ;
        RECT 35.045 155.575 36.680 155.815 ;
        RECT 35.045 155.485 35.275 155.575 ;
        RECT 35.385 155.315 35.715 155.355 ;
        RECT 34.545 155.145 35.715 155.315 ;
        RECT 35.905 154.975 36.260 155.395 ;
        RECT 36.430 155.145 36.680 155.575 ;
        RECT 36.850 154.975 37.180 155.735 ;
        RECT 37.350 155.145 37.605 155.815 ;
        RECT 37.795 155.955 38.955 156.165 ;
        RECT 37.795 155.145 38.115 155.955 ;
        RECT 38.285 154.975 38.535 155.785 ;
        RECT 38.705 155.315 38.955 155.955 ;
        RECT 39.125 155.485 39.375 156.715 ;
        RECT 39.925 156.535 40.140 156.715 ;
        RECT 39.585 156.365 40.140 156.535 ;
        RECT 39.970 156.165 40.140 156.365 ;
        RECT 40.310 156.335 40.835 156.545 ;
        RECT 39.545 155.720 39.800 156.165 ;
        RECT 39.970 155.995 40.275 156.165 ;
        RECT 39.545 155.315 39.835 155.720 ;
        RECT 38.705 155.145 39.835 155.315 ;
        RECT 40.105 155.150 40.275 155.995 ;
        RECT 40.620 155.825 40.835 156.335 ;
        RECT 40.615 155.655 40.835 155.825 ;
        RECT 40.620 155.645 40.835 155.655 ;
        RECT 41.475 156.115 41.645 157.025 ;
        RECT 42.400 156.875 42.695 157.265 ;
        RECT 42.865 157.045 43.120 157.525 ;
        RECT 43.295 156.875 43.555 157.265 ;
        RECT 43.725 157.045 44.005 157.525 ;
        RECT 44.235 157.035 44.505 157.525 ;
        RECT 41.815 156.285 42.165 156.855 ;
        RECT 42.400 156.705 44.050 156.875 ;
        RECT 42.335 156.365 43.475 156.535 ;
        RECT 42.335 156.115 42.505 156.365 ;
        RECT 43.645 156.195 44.050 156.705 ;
        RECT 44.295 156.285 44.560 156.865 ;
        RECT 44.730 156.595 45.005 157.305 ;
        RECT 45.205 157.040 45.990 157.305 ;
        RECT 44.730 156.365 45.565 156.595 ;
        RECT 41.475 155.945 42.505 156.115 ;
        RECT 43.295 156.025 44.050 156.195 ;
        RECT 40.485 154.975 40.735 155.465 ;
        RECT 41.475 155.145 41.785 155.945 ;
        RECT 43.295 155.775 43.555 156.025 ;
        RECT 41.955 154.975 42.265 155.775 ;
        RECT 42.435 155.605 43.555 155.775 ;
        RECT 42.435 155.145 42.695 155.605 ;
        RECT 42.865 154.975 43.120 155.435 ;
        RECT 43.295 155.145 43.555 155.605 ;
        RECT 43.725 154.975 44.010 155.845 ;
        RECT 44.235 154.975 44.550 156.035 ;
        RECT 44.730 155.705 45.005 156.365 ;
        RECT 45.735 156.185 45.990 157.040 ;
        RECT 46.160 156.845 46.370 157.305 ;
        RECT 46.560 157.030 46.890 157.525 ;
        RECT 47.065 156.895 47.310 157.355 ;
        RECT 46.160 156.365 46.570 156.845 ;
        RECT 47.140 156.685 47.310 156.895 ;
        RECT 47.480 156.865 47.745 157.525 ;
        RECT 47.915 156.850 48.190 157.195 ;
        RECT 48.380 157.125 48.755 157.525 ;
        RECT 48.925 156.955 49.095 157.305 ;
        RECT 49.265 157.125 49.595 157.525 ;
        RECT 49.765 156.955 50.025 157.355 ;
        RECT 46.740 156.185 46.970 156.615 ;
        RECT 45.200 156.015 46.970 156.185 ;
        RECT 47.140 156.165 47.745 156.685 ;
        RECT 45.200 155.650 45.435 156.015 ;
        RECT 45.605 155.655 45.935 155.845 ;
        RECT 46.160 155.720 46.350 156.015 ;
        RECT 47.140 155.825 47.310 156.165 ;
        RECT 47.915 156.115 48.085 156.850 ;
        RECT 48.360 156.785 50.025 156.955 ;
        RECT 48.360 156.615 48.530 156.785 ;
        RECT 50.205 156.705 50.535 157.125 ;
        RECT 50.705 156.705 50.965 157.525 ;
        RECT 51.135 156.865 51.410 157.525 ;
        RECT 51.580 156.895 51.830 157.355 ;
        RECT 52.005 157.030 52.335 157.525 ;
        RECT 50.205 156.615 50.455 156.705 ;
        RECT 51.580 156.685 51.750 156.895 ;
        RECT 52.515 156.860 52.745 157.305 ;
        RECT 48.255 156.285 48.530 156.615 ;
        RECT 48.700 156.285 49.525 156.615 ;
        RECT 49.740 156.285 50.455 156.615 ;
        RECT 50.625 156.285 50.960 156.535 ;
        RECT 48.360 156.115 48.530 156.285 ;
        RECT 45.605 155.480 45.795 155.655 ;
        RECT 45.180 154.975 45.795 155.480 ;
        RECT 45.965 155.145 46.440 155.485 ;
        RECT 46.610 154.975 46.825 155.820 ;
        RECT 47.055 155.815 47.310 155.825 ;
        RECT 47.025 155.145 47.310 155.815 ;
        RECT 47.480 154.975 47.745 155.985 ;
        RECT 47.915 155.145 48.190 156.115 ;
        RECT 48.360 155.945 49.020 156.115 ;
        RECT 49.280 155.995 49.525 156.285 ;
        RECT 48.850 155.825 49.020 155.945 ;
        RECT 49.695 155.825 50.025 156.115 ;
        RECT 48.400 154.975 48.680 155.775 ;
        RECT 48.850 155.655 50.025 155.825 ;
        RECT 50.285 155.725 50.455 156.285 ;
        RECT 51.135 156.165 51.750 156.685 ;
        RECT 51.920 156.185 52.150 156.615 ;
        RECT 52.335 156.365 52.745 156.860 ;
        RECT 52.915 157.040 53.705 157.305 ;
        RECT 52.915 156.185 53.170 157.040 ;
        RECT 53.340 156.365 53.725 156.845 ;
        RECT 54.355 156.800 54.645 157.525 ;
        RECT 54.815 156.865 55.090 157.525 ;
        RECT 55.260 156.895 55.510 157.355 ;
        RECT 55.685 157.030 56.015 157.525 ;
        RECT 55.260 156.685 55.430 156.895 ;
        RECT 56.195 156.860 56.425 157.305 ;
        RECT 48.850 155.155 50.465 155.485 ;
        RECT 50.705 154.975 50.965 156.115 ;
        RECT 51.135 154.975 51.395 155.985 ;
        RECT 51.565 155.815 51.735 156.165 ;
        RECT 51.920 156.015 53.710 156.185 ;
        RECT 54.815 156.165 55.430 156.685 ;
        RECT 55.600 156.185 55.830 156.615 ;
        RECT 56.015 156.365 56.425 156.860 ;
        RECT 56.595 157.040 57.385 157.305 ;
        RECT 56.595 156.185 56.850 157.040 ;
        RECT 58.035 157.025 58.335 157.355 ;
        RECT 58.505 157.045 58.780 157.525 ;
        RECT 57.020 156.365 57.405 156.845 ;
        RECT 51.565 155.145 51.840 155.815 ;
        RECT 52.040 154.975 52.255 155.820 ;
        RECT 52.480 155.720 52.730 156.015 ;
        RECT 52.955 155.655 53.285 155.845 ;
        RECT 52.440 155.145 52.915 155.485 ;
        RECT 53.095 155.480 53.285 155.655 ;
        RECT 53.455 155.650 53.710 156.015 ;
        RECT 53.095 154.975 53.725 155.480 ;
        RECT 54.355 154.975 54.645 156.140 ;
        RECT 54.815 154.975 55.075 155.985 ;
        RECT 55.245 155.815 55.415 156.165 ;
        RECT 55.600 156.015 57.390 156.185 ;
        RECT 55.245 155.145 55.520 155.815 ;
        RECT 55.720 154.975 55.935 155.820 ;
        RECT 56.160 155.720 56.410 156.015 ;
        RECT 56.635 155.655 56.965 155.845 ;
        RECT 56.120 155.145 56.595 155.485 ;
        RECT 56.775 155.480 56.965 155.655 ;
        RECT 57.135 155.650 57.390 156.015 ;
        RECT 58.035 156.115 58.205 157.025 ;
        RECT 58.960 156.875 59.255 157.265 ;
        RECT 59.425 157.045 59.680 157.525 ;
        RECT 59.855 156.875 60.115 157.265 ;
        RECT 60.285 157.045 60.565 157.525 ;
        RECT 58.375 156.285 58.725 156.855 ;
        RECT 58.960 156.705 60.610 156.875 ;
        RECT 58.895 156.365 60.035 156.535 ;
        RECT 58.895 156.115 59.065 156.365 ;
        RECT 60.205 156.195 60.610 156.705 ;
        RECT 58.035 155.945 59.065 156.115 ;
        RECT 59.855 156.025 60.610 156.195 ;
        RECT 61.720 156.785 61.975 157.355 ;
        RECT 62.145 157.125 62.475 157.525 ;
        RECT 62.900 156.990 63.430 157.355 ;
        RECT 63.620 157.185 63.895 157.355 ;
        RECT 63.615 157.015 63.895 157.185 ;
        RECT 62.900 156.955 63.075 156.990 ;
        RECT 62.145 156.785 63.075 156.955 ;
        RECT 61.720 156.115 61.890 156.785 ;
        RECT 62.145 156.615 62.315 156.785 ;
        RECT 62.060 156.285 62.315 156.615 ;
        RECT 62.540 156.285 62.735 156.615 ;
        RECT 56.775 154.975 57.405 155.480 ;
        RECT 58.035 155.145 58.345 155.945 ;
        RECT 59.855 155.775 60.115 156.025 ;
        RECT 58.515 154.975 58.825 155.775 ;
        RECT 58.995 155.605 60.115 155.775 ;
        RECT 58.995 155.145 59.255 155.605 ;
        RECT 59.425 154.975 59.680 155.435 ;
        RECT 59.855 155.145 60.115 155.605 ;
        RECT 60.285 154.975 60.570 155.845 ;
        RECT 61.720 155.145 62.055 156.115 ;
        RECT 62.225 154.975 62.395 156.115 ;
        RECT 62.565 155.315 62.735 156.285 ;
        RECT 62.905 155.655 63.075 156.785 ;
        RECT 63.245 155.995 63.415 156.795 ;
        RECT 63.620 156.195 63.895 157.015 ;
        RECT 64.065 155.995 64.255 157.355 ;
        RECT 64.435 156.990 64.945 157.525 ;
        RECT 65.165 156.715 65.410 157.320 ;
        RECT 65.860 156.975 66.115 157.265 ;
        RECT 66.285 157.145 66.615 157.525 ;
        RECT 65.860 156.805 66.610 156.975 ;
        RECT 64.455 156.545 65.685 156.715 ;
        RECT 63.245 155.825 64.255 155.995 ;
        RECT 64.425 155.980 65.175 156.170 ;
        RECT 62.905 155.485 64.030 155.655 ;
        RECT 64.425 155.315 64.595 155.980 ;
        RECT 65.345 155.735 65.685 156.545 ;
        RECT 65.860 155.985 66.210 156.635 ;
        RECT 66.380 155.815 66.610 156.805 ;
        RECT 62.565 155.145 64.595 155.315 ;
        RECT 64.765 154.975 64.935 155.735 ;
        RECT 65.170 155.325 65.685 155.735 ;
        RECT 65.860 155.645 66.610 155.815 ;
        RECT 65.860 155.145 66.115 155.645 ;
        RECT 66.285 154.975 66.615 155.475 ;
        RECT 66.785 155.145 66.955 157.265 ;
        RECT 67.315 157.165 67.645 157.525 ;
        RECT 67.815 157.135 68.310 157.305 ;
        RECT 68.515 157.135 69.370 157.305 ;
        RECT 67.185 155.945 67.645 156.995 ;
        RECT 67.125 155.160 67.450 155.945 ;
        RECT 67.815 155.775 67.985 157.135 ;
        RECT 68.155 156.225 68.505 156.845 ;
        RECT 68.675 156.625 69.030 156.845 ;
        RECT 68.675 156.035 68.845 156.625 ;
        RECT 69.200 156.425 69.370 157.135 ;
        RECT 70.245 157.065 70.575 157.525 ;
        RECT 70.785 157.165 71.135 157.335 ;
        RECT 69.575 156.595 70.365 156.845 ;
        RECT 70.785 156.775 71.045 157.165 ;
        RECT 71.355 157.075 72.305 157.355 ;
        RECT 72.475 157.085 72.665 157.525 ;
        RECT 72.835 157.145 73.905 157.315 ;
        RECT 70.535 156.425 70.705 156.605 ;
        RECT 67.815 155.605 68.210 155.775 ;
        RECT 68.380 155.645 68.845 156.035 ;
        RECT 69.015 156.255 70.705 156.425 ;
        RECT 68.040 155.475 68.210 155.605 ;
        RECT 69.015 155.475 69.185 156.255 ;
        RECT 70.875 156.085 71.045 156.775 ;
        RECT 69.545 155.915 71.045 156.085 ;
        RECT 71.235 156.115 71.445 156.905 ;
        RECT 71.615 156.285 71.965 156.905 ;
        RECT 72.135 156.295 72.305 157.075 ;
        RECT 72.835 156.915 73.005 157.145 ;
        RECT 72.475 156.745 73.005 156.915 ;
        RECT 72.475 156.465 72.695 156.745 ;
        RECT 73.175 156.575 73.415 156.975 ;
        RECT 72.135 156.125 72.540 156.295 ;
        RECT 72.875 156.205 73.415 156.575 ;
        RECT 73.585 156.790 73.905 157.145 ;
        RECT 74.150 157.065 74.455 157.525 ;
        RECT 74.625 156.815 74.880 157.345 ;
        RECT 73.585 156.615 73.910 156.790 ;
        RECT 73.585 156.315 74.500 156.615 ;
        RECT 73.760 156.285 74.500 156.315 ;
        RECT 71.235 155.955 71.910 156.115 ;
        RECT 72.370 156.035 72.540 156.125 ;
        RECT 71.235 155.945 72.200 155.955 ;
        RECT 70.875 155.775 71.045 155.915 ;
        RECT 67.620 154.975 67.870 155.435 ;
        RECT 68.040 155.145 68.290 155.475 ;
        RECT 68.505 155.145 69.185 155.475 ;
        RECT 69.355 155.575 70.430 155.745 ;
        RECT 70.875 155.605 71.435 155.775 ;
        RECT 71.740 155.655 72.200 155.945 ;
        RECT 72.370 155.865 73.590 156.035 ;
        RECT 69.355 155.235 69.525 155.575 ;
        RECT 69.760 154.975 70.090 155.405 ;
        RECT 70.260 155.235 70.430 155.575 ;
        RECT 70.725 154.975 71.095 155.435 ;
        RECT 71.265 155.145 71.435 155.605 ;
        RECT 72.370 155.485 72.540 155.865 ;
        RECT 73.760 155.695 73.930 156.285 ;
        RECT 74.670 156.165 74.880 156.815 ;
        RECT 75.980 156.725 76.235 157.525 ;
        RECT 76.405 156.860 76.655 157.355 ;
        RECT 76.825 157.145 77.155 157.525 ;
        RECT 77.325 157.145 78.620 157.315 ;
        RECT 77.325 156.975 77.495 157.145 ;
        RECT 71.670 155.145 72.540 155.485 ;
        RECT 73.130 155.525 73.930 155.695 ;
        RECT 72.710 154.975 72.960 155.435 ;
        RECT 73.130 155.235 73.300 155.525 ;
        RECT 73.480 154.975 73.810 155.355 ;
        RECT 74.150 154.975 74.455 156.115 ;
        RECT 74.625 155.285 74.880 156.165 ;
        RECT 75.980 154.975 76.235 156.115 ;
        RECT 76.405 156.015 76.575 156.860 ;
        RECT 76.885 156.805 77.495 156.975 ;
        RECT 78.790 156.875 78.980 157.190 ;
        RECT 79.240 157.025 79.440 157.525 ;
        RECT 76.885 156.615 77.055 156.805 ;
        RECT 76.745 156.285 77.055 156.615 ;
        RECT 76.405 155.145 76.715 156.015 ;
        RECT 76.885 155.775 77.055 156.285 ;
        RECT 77.225 156.115 77.395 156.615 ;
        RECT 77.705 156.330 78.335 156.845 ;
        RECT 78.515 156.585 78.980 156.875 ;
        RECT 78.165 156.295 78.335 156.330 ;
        RECT 77.225 155.945 77.885 156.115 ;
        RECT 78.165 155.985 78.980 156.295 ;
        RECT 79.250 155.985 79.440 156.855 ;
        RECT 77.715 155.775 77.885 155.945 ;
        RECT 79.610 155.775 79.940 157.355 ;
        RECT 80.115 156.800 80.405 157.525 ;
        RECT 81.125 156.975 81.295 157.355 ;
        RECT 81.510 157.145 81.840 157.525 ;
        RECT 81.125 156.805 81.840 156.975 ;
        RECT 81.035 156.255 81.390 156.625 ;
        RECT 81.670 156.615 81.840 156.805 ;
        RECT 82.010 156.780 82.265 157.355 ;
        RECT 81.670 156.285 81.925 156.615 ;
        RECT 76.885 155.605 77.545 155.775 ;
        RECT 77.715 155.605 79.940 155.775 ;
        RECT 76.915 154.975 77.205 155.435 ;
        RECT 77.375 155.355 77.545 155.605 ;
        RECT 77.375 155.185 78.685 155.355 ;
        RECT 79.215 154.975 79.435 155.435 ;
        RECT 79.605 155.145 79.940 155.605 ;
        RECT 80.115 154.975 80.405 156.140 ;
        RECT 81.670 156.075 81.840 156.285 ;
        RECT 81.125 155.905 81.840 156.075 ;
        RECT 82.095 156.050 82.265 156.780 ;
        RECT 82.440 156.685 82.700 157.525 ;
        RECT 82.880 156.815 83.135 157.345 ;
        RECT 83.305 157.065 83.610 157.525 ;
        RECT 83.855 157.145 84.925 157.315 ;
        RECT 82.880 156.165 83.090 156.815 ;
        RECT 83.855 156.790 84.175 157.145 ;
        RECT 83.850 156.615 84.175 156.790 ;
        RECT 83.260 156.315 84.175 156.615 ;
        RECT 84.345 156.575 84.585 156.975 ;
        RECT 84.755 156.915 84.925 157.145 ;
        RECT 85.095 157.085 85.285 157.525 ;
        RECT 85.455 157.075 86.405 157.355 ;
        RECT 86.625 157.165 86.975 157.335 ;
        RECT 84.755 156.745 85.285 156.915 ;
        RECT 83.260 156.285 84.000 156.315 ;
        RECT 81.125 155.145 81.295 155.905 ;
        RECT 81.510 154.975 81.840 155.735 ;
        RECT 82.010 155.145 82.265 156.050 ;
        RECT 82.440 154.975 82.700 156.125 ;
        RECT 82.880 155.285 83.135 156.165 ;
        RECT 83.305 154.975 83.610 156.115 ;
        RECT 83.830 155.695 84.000 156.285 ;
        RECT 84.345 156.205 84.885 156.575 ;
        RECT 85.065 156.465 85.285 156.745 ;
        RECT 85.455 156.295 85.625 157.075 ;
        RECT 85.220 156.125 85.625 156.295 ;
        RECT 85.795 156.285 86.145 156.905 ;
        RECT 85.220 156.035 85.390 156.125 ;
        RECT 86.315 156.115 86.525 156.905 ;
        RECT 84.170 155.865 85.390 156.035 ;
        RECT 85.850 155.955 86.525 156.115 ;
        RECT 83.830 155.525 84.630 155.695 ;
        RECT 83.950 154.975 84.280 155.355 ;
        RECT 84.460 155.235 84.630 155.525 ;
        RECT 85.220 155.485 85.390 155.865 ;
        RECT 85.560 155.945 86.525 155.955 ;
        RECT 86.715 156.775 86.975 157.165 ;
        RECT 87.185 157.065 87.515 157.525 ;
        RECT 88.390 157.135 89.245 157.305 ;
        RECT 89.450 157.135 89.945 157.305 ;
        RECT 90.115 157.165 90.445 157.525 ;
        RECT 86.715 156.085 86.885 156.775 ;
        RECT 87.055 156.425 87.225 156.605 ;
        RECT 87.395 156.595 88.185 156.845 ;
        RECT 88.390 156.425 88.560 157.135 ;
        RECT 88.730 156.625 89.085 156.845 ;
        RECT 87.055 156.255 88.745 156.425 ;
        RECT 85.560 155.655 86.020 155.945 ;
        RECT 86.715 155.915 88.215 156.085 ;
        RECT 86.715 155.775 86.885 155.915 ;
        RECT 86.325 155.605 86.885 155.775 ;
        RECT 84.800 154.975 85.050 155.435 ;
        RECT 85.220 155.145 86.090 155.485 ;
        RECT 86.325 155.145 86.495 155.605 ;
        RECT 87.330 155.575 88.405 155.745 ;
        RECT 86.665 154.975 87.035 155.435 ;
        RECT 87.330 155.235 87.500 155.575 ;
        RECT 87.670 154.975 88.000 155.405 ;
        RECT 88.235 155.235 88.405 155.575 ;
        RECT 88.575 155.475 88.745 156.255 ;
        RECT 88.915 156.035 89.085 156.625 ;
        RECT 89.255 156.225 89.605 156.845 ;
        RECT 88.915 155.645 89.380 156.035 ;
        RECT 89.775 155.775 89.945 157.135 ;
        RECT 90.115 155.945 90.575 156.995 ;
        RECT 89.550 155.605 89.945 155.775 ;
        RECT 89.550 155.475 89.720 155.605 ;
        RECT 88.575 155.145 89.255 155.475 ;
        RECT 89.470 155.145 89.720 155.475 ;
        RECT 89.890 154.975 90.140 155.435 ;
        RECT 90.310 155.160 90.635 155.945 ;
        RECT 90.805 155.145 90.975 157.265 ;
        RECT 91.145 157.145 91.475 157.525 ;
        RECT 91.645 156.975 91.900 157.265 ;
        RECT 91.150 156.805 91.900 156.975 ;
        RECT 92.075 157.025 92.375 157.355 ;
        RECT 92.545 157.045 92.820 157.525 ;
        RECT 91.150 155.815 91.380 156.805 ;
        RECT 91.550 155.985 91.900 156.635 ;
        RECT 92.075 156.115 92.245 157.025 ;
        RECT 93.000 156.875 93.295 157.265 ;
        RECT 93.465 157.045 93.720 157.525 ;
        RECT 93.895 156.875 94.155 157.265 ;
        RECT 94.325 157.045 94.605 157.525 ;
        RECT 92.415 156.285 92.765 156.855 ;
        RECT 93.000 156.705 94.650 156.875 ;
        RECT 96.030 156.715 96.275 157.320 ;
        RECT 96.495 156.990 97.005 157.525 ;
        RECT 92.935 156.365 94.075 156.535 ;
        RECT 92.935 156.115 93.105 156.365 ;
        RECT 94.245 156.195 94.650 156.705 ;
        RECT 92.075 155.945 93.105 156.115 ;
        RECT 93.895 156.025 94.650 156.195 ;
        RECT 95.755 156.545 96.985 156.715 ;
        RECT 91.150 155.645 91.900 155.815 ;
        RECT 91.145 154.975 91.475 155.475 ;
        RECT 91.645 155.145 91.900 155.645 ;
        RECT 92.075 155.145 92.385 155.945 ;
        RECT 93.895 155.775 94.155 156.025 ;
        RECT 92.555 154.975 92.865 155.775 ;
        RECT 93.035 155.605 94.155 155.775 ;
        RECT 93.035 155.145 93.295 155.605 ;
        RECT 93.465 154.975 93.720 155.435 ;
        RECT 93.895 155.145 94.155 155.605 ;
        RECT 94.325 154.975 94.610 155.845 ;
        RECT 95.755 155.735 96.095 156.545 ;
        RECT 96.265 155.980 97.015 156.170 ;
        RECT 95.755 155.325 96.270 155.735 ;
        RECT 96.505 154.975 96.675 155.735 ;
        RECT 96.845 155.315 97.015 155.980 ;
        RECT 97.185 155.995 97.375 157.355 ;
        RECT 97.545 156.505 97.820 157.355 ;
        RECT 98.010 156.990 98.540 157.355 ;
        RECT 98.965 157.125 99.295 157.525 ;
        RECT 98.365 156.955 98.540 156.990 ;
        RECT 97.545 156.335 97.825 156.505 ;
        RECT 97.545 156.195 97.820 156.335 ;
        RECT 98.025 155.995 98.195 156.795 ;
        RECT 97.185 155.825 98.195 155.995 ;
        RECT 98.365 156.785 99.295 156.955 ;
        RECT 99.465 156.785 99.720 157.355 ;
        RECT 98.365 155.655 98.535 156.785 ;
        RECT 99.125 156.615 99.295 156.785 ;
        RECT 97.410 155.485 98.535 155.655 ;
        RECT 98.705 156.285 98.900 156.615 ;
        RECT 99.125 156.285 99.380 156.615 ;
        RECT 98.705 155.315 98.875 156.285 ;
        RECT 99.550 156.115 99.720 156.785 ;
        RECT 96.845 155.145 98.875 155.315 ;
        RECT 99.045 154.975 99.215 156.115 ;
        RECT 99.385 155.145 99.720 156.115 ;
        RECT 99.895 156.850 100.155 157.355 ;
        RECT 100.335 157.145 100.665 157.525 ;
        RECT 100.845 156.975 101.015 157.355 ;
        RECT 99.895 156.050 100.065 156.850 ;
        RECT 100.350 156.805 101.015 156.975 ;
        RECT 101.825 156.975 101.995 157.355 ;
        RECT 102.175 157.145 102.505 157.525 ;
        RECT 101.825 156.805 102.490 156.975 ;
        RECT 102.685 156.850 102.945 157.355 ;
        RECT 103.175 157.045 103.455 157.525 ;
        RECT 103.625 156.875 103.885 157.265 ;
        RECT 104.060 157.045 104.315 157.525 ;
        RECT 104.485 156.875 104.780 157.265 ;
        RECT 104.960 157.045 105.235 157.525 ;
        RECT 105.405 157.025 105.705 157.355 ;
        RECT 100.350 156.550 100.520 156.805 ;
        RECT 100.235 156.220 100.520 156.550 ;
        RECT 100.755 156.255 101.085 156.625 ;
        RECT 101.755 156.255 102.085 156.625 ;
        RECT 102.320 156.550 102.490 156.805 ;
        RECT 100.350 156.075 100.520 156.220 ;
        RECT 102.320 156.220 102.605 156.550 ;
        RECT 102.320 156.075 102.490 156.220 ;
        RECT 99.895 155.145 100.165 156.050 ;
        RECT 100.350 155.905 101.015 156.075 ;
        RECT 100.335 154.975 100.665 155.735 ;
        RECT 100.845 155.145 101.015 155.905 ;
        RECT 101.825 155.905 102.490 156.075 ;
        RECT 102.775 156.050 102.945 156.850 ;
        RECT 101.825 155.145 101.995 155.905 ;
        RECT 102.175 154.975 102.505 155.735 ;
        RECT 102.675 155.145 102.945 156.050 ;
        RECT 103.130 156.705 104.780 156.875 ;
        RECT 103.130 156.195 103.535 156.705 ;
        RECT 103.705 156.365 104.845 156.535 ;
        RECT 103.130 156.025 103.885 156.195 ;
        RECT 103.170 154.975 103.455 155.845 ;
        RECT 103.625 155.775 103.885 156.025 ;
        RECT 104.675 156.115 104.845 156.365 ;
        RECT 105.015 156.285 105.365 156.855 ;
        RECT 105.535 156.115 105.705 157.025 ;
        RECT 105.875 156.800 106.165 157.525 ;
        RECT 106.340 156.785 106.595 157.355 ;
        RECT 106.765 157.125 107.095 157.525 ;
        RECT 107.520 156.990 108.050 157.355 ;
        RECT 108.240 157.185 108.515 157.355 ;
        RECT 108.235 157.015 108.515 157.185 ;
        RECT 107.520 156.955 107.695 156.990 ;
        RECT 106.765 156.785 107.695 156.955 ;
        RECT 104.675 155.945 105.705 156.115 ;
        RECT 103.625 155.605 104.745 155.775 ;
        RECT 103.625 155.145 103.885 155.605 ;
        RECT 104.060 154.975 104.315 155.435 ;
        RECT 104.485 155.145 104.745 155.605 ;
        RECT 104.915 154.975 105.225 155.775 ;
        RECT 105.395 155.145 105.705 155.945 ;
        RECT 105.875 154.975 106.165 156.140 ;
        RECT 106.340 156.115 106.510 156.785 ;
        RECT 106.765 156.615 106.935 156.785 ;
        RECT 106.680 156.285 106.935 156.615 ;
        RECT 107.160 156.285 107.355 156.615 ;
        RECT 106.340 155.145 106.675 156.115 ;
        RECT 106.845 154.975 107.015 156.115 ;
        RECT 107.185 155.315 107.355 156.285 ;
        RECT 107.525 155.655 107.695 156.785 ;
        RECT 107.865 155.995 108.035 156.795 ;
        RECT 108.240 156.195 108.515 157.015 ;
        RECT 108.685 155.995 108.875 157.355 ;
        RECT 109.055 156.990 109.565 157.525 ;
        RECT 109.785 156.715 110.030 157.320 ;
        RECT 110.935 156.715 111.215 157.525 ;
        RECT 111.385 156.885 111.715 157.355 ;
        RECT 111.885 157.055 112.055 157.525 ;
        RECT 112.225 156.885 112.555 157.355 ;
        RECT 111.385 156.715 112.555 156.885 ;
        RECT 112.725 156.715 112.895 157.525 ;
        RECT 113.245 156.885 113.415 157.165 ;
        RECT 113.065 156.715 113.415 156.885 ;
        RECT 113.625 156.765 113.880 157.525 ;
        RECT 114.160 156.975 114.415 157.265 ;
        RECT 114.585 157.145 114.915 157.525 ;
        RECT 114.160 156.805 114.910 156.975 ;
        RECT 109.075 156.545 110.305 156.715 ;
        RECT 107.865 155.825 108.875 155.995 ;
        RECT 109.045 155.980 109.795 156.170 ;
        RECT 107.525 155.485 108.650 155.655 ;
        RECT 109.045 155.315 109.215 155.980 ;
        RECT 109.965 155.735 110.305 156.545 ;
        RECT 111.330 156.335 111.770 156.545 ;
        RECT 112.265 156.505 112.515 156.715 ;
        RECT 113.065 156.535 113.280 156.715 ;
        RECT 112.265 156.335 112.545 156.505 ;
        RECT 112.725 156.365 113.280 156.535 ;
        RECT 107.185 155.145 109.215 155.315 ;
        RECT 109.385 154.975 109.555 155.735 ;
        RECT 109.790 155.325 110.305 155.735 ;
        RECT 110.935 155.955 112.095 156.165 ;
        RECT 110.935 155.145 111.255 155.955 ;
        RECT 111.425 154.975 111.675 155.785 ;
        RECT 111.845 155.315 112.095 155.955 ;
        RECT 112.265 155.485 112.515 156.335 ;
        RECT 113.110 156.165 113.280 156.365 ;
        RECT 113.450 156.335 113.975 156.545 ;
        RECT 112.685 155.720 112.940 156.165 ;
        RECT 113.110 155.995 113.415 156.165 ;
        RECT 112.685 155.315 112.975 155.720 ;
        RECT 111.845 155.145 112.975 155.315 ;
        RECT 113.245 155.150 113.415 155.995 ;
        RECT 113.760 155.825 113.975 156.335 ;
        RECT 114.160 155.985 114.510 156.635 ;
        RECT 113.755 155.655 113.975 155.825 ;
        RECT 114.680 155.815 114.910 156.805 ;
        RECT 113.760 155.645 113.975 155.655 ;
        RECT 114.160 155.645 114.910 155.815 ;
        RECT 113.625 154.975 113.875 155.465 ;
        RECT 114.160 155.145 114.415 155.645 ;
        RECT 114.585 154.975 114.915 155.475 ;
        RECT 115.085 155.145 115.255 157.265 ;
        RECT 115.615 157.165 115.945 157.525 ;
        RECT 116.115 157.135 116.610 157.305 ;
        RECT 116.815 157.135 117.670 157.305 ;
        RECT 115.485 155.945 115.945 156.995 ;
        RECT 115.425 155.160 115.750 155.945 ;
        RECT 116.115 155.775 116.285 157.135 ;
        RECT 116.455 156.225 116.805 156.845 ;
        RECT 116.975 156.625 117.330 156.845 ;
        RECT 116.975 156.035 117.145 156.625 ;
        RECT 117.500 156.425 117.670 157.135 ;
        RECT 118.545 157.065 118.875 157.525 ;
        RECT 119.085 157.165 119.435 157.335 ;
        RECT 117.875 156.595 118.665 156.845 ;
        RECT 119.085 156.775 119.345 157.165 ;
        RECT 119.655 157.075 120.605 157.355 ;
        RECT 120.775 157.085 120.965 157.525 ;
        RECT 121.135 157.145 122.205 157.315 ;
        RECT 118.835 156.425 119.005 156.605 ;
        RECT 116.115 155.605 116.510 155.775 ;
        RECT 116.680 155.645 117.145 156.035 ;
        RECT 117.315 156.255 119.005 156.425 ;
        RECT 116.340 155.475 116.510 155.605 ;
        RECT 117.315 155.475 117.485 156.255 ;
        RECT 119.175 156.085 119.345 156.775 ;
        RECT 117.845 155.915 119.345 156.085 ;
        RECT 119.535 156.115 119.745 156.905 ;
        RECT 119.915 156.285 120.265 156.905 ;
        RECT 120.435 156.295 120.605 157.075 ;
        RECT 121.135 156.915 121.305 157.145 ;
        RECT 120.775 156.745 121.305 156.915 ;
        RECT 120.775 156.465 120.995 156.745 ;
        RECT 121.475 156.575 121.715 156.975 ;
        RECT 120.435 156.125 120.840 156.295 ;
        RECT 121.175 156.205 121.715 156.575 ;
        RECT 121.885 156.790 122.205 157.145 ;
        RECT 122.450 157.065 122.755 157.525 ;
        RECT 122.925 156.815 123.175 157.345 ;
        RECT 121.885 156.615 122.210 156.790 ;
        RECT 121.885 156.315 122.800 156.615 ;
        RECT 122.060 156.285 122.800 156.315 ;
        RECT 119.535 155.955 120.210 156.115 ;
        RECT 120.670 156.035 120.840 156.125 ;
        RECT 119.535 155.945 120.500 155.955 ;
        RECT 119.175 155.775 119.345 155.915 ;
        RECT 115.920 154.975 116.170 155.435 ;
        RECT 116.340 155.145 116.590 155.475 ;
        RECT 116.805 155.145 117.485 155.475 ;
        RECT 117.655 155.575 118.730 155.745 ;
        RECT 119.175 155.605 119.735 155.775 ;
        RECT 120.040 155.655 120.500 155.945 ;
        RECT 120.670 155.865 121.890 156.035 ;
        RECT 117.655 155.235 117.825 155.575 ;
        RECT 118.060 154.975 118.390 155.405 ;
        RECT 118.560 155.235 118.730 155.575 ;
        RECT 119.025 154.975 119.395 155.435 ;
        RECT 119.565 155.145 119.735 155.605 ;
        RECT 120.670 155.485 120.840 155.865 ;
        RECT 122.060 155.695 122.230 156.285 ;
        RECT 122.970 156.165 123.175 156.815 ;
        RECT 123.345 156.770 123.595 157.525 ;
        RECT 124.275 156.850 124.535 157.355 ;
        RECT 124.715 157.145 125.045 157.525 ;
        RECT 125.225 156.975 125.395 157.355 ;
        RECT 119.970 155.145 120.840 155.485 ;
        RECT 121.430 155.525 122.230 155.695 ;
        RECT 121.010 154.975 121.260 155.435 ;
        RECT 121.430 155.235 121.600 155.525 ;
        RECT 121.780 154.975 122.110 155.355 ;
        RECT 122.450 154.975 122.755 156.115 ;
        RECT 122.925 155.285 123.175 156.165 ;
        RECT 123.345 154.975 123.595 156.115 ;
        RECT 124.275 156.050 124.445 156.850 ;
        RECT 124.730 156.805 125.395 156.975 ;
        RECT 124.730 156.550 124.900 156.805 ;
        RECT 125.660 156.785 125.915 157.355 ;
        RECT 126.085 157.125 126.415 157.525 ;
        RECT 126.840 156.990 127.370 157.355 ;
        RECT 126.840 156.955 127.015 156.990 ;
        RECT 126.085 156.785 127.015 156.955 ;
        RECT 127.560 156.845 127.835 157.355 ;
        RECT 124.615 156.220 124.900 156.550 ;
        RECT 125.135 156.255 125.465 156.625 ;
        RECT 124.730 156.075 124.900 156.220 ;
        RECT 125.660 156.115 125.830 156.785 ;
        RECT 126.085 156.615 126.255 156.785 ;
        RECT 126.000 156.285 126.255 156.615 ;
        RECT 126.480 156.285 126.675 156.615 ;
        RECT 124.275 155.145 124.545 156.050 ;
        RECT 124.730 155.905 125.395 156.075 ;
        RECT 124.715 154.975 125.045 155.735 ;
        RECT 125.225 155.145 125.395 155.905 ;
        RECT 125.660 155.145 125.995 156.115 ;
        RECT 126.165 154.975 126.335 156.115 ;
        RECT 126.505 155.315 126.675 156.285 ;
        RECT 126.845 155.655 127.015 156.785 ;
        RECT 127.185 155.995 127.355 156.795 ;
        RECT 127.555 156.675 127.835 156.845 ;
        RECT 127.560 156.195 127.835 156.675 ;
        RECT 128.005 155.995 128.195 157.355 ;
        RECT 128.375 156.990 128.885 157.525 ;
        RECT 129.105 156.715 129.350 157.320 ;
        RECT 130.345 156.975 130.515 157.355 ;
        RECT 130.695 157.145 131.025 157.525 ;
        RECT 130.345 156.805 131.010 156.975 ;
        RECT 131.205 156.850 131.465 157.355 ;
        RECT 128.395 156.545 129.625 156.715 ;
        RECT 127.185 155.825 128.195 155.995 ;
        RECT 128.365 155.980 129.115 156.170 ;
        RECT 126.845 155.485 127.970 155.655 ;
        RECT 128.365 155.315 128.535 155.980 ;
        RECT 129.285 155.735 129.625 156.545 ;
        RECT 130.275 156.255 130.605 156.625 ;
        RECT 130.840 156.550 131.010 156.805 ;
        RECT 130.840 156.220 131.125 156.550 ;
        RECT 130.840 156.075 131.010 156.220 ;
        RECT 126.505 155.145 128.535 155.315 ;
        RECT 128.705 154.975 128.875 155.735 ;
        RECT 129.110 155.325 129.625 155.735 ;
        RECT 130.345 155.905 131.010 156.075 ;
        RECT 131.295 156.050 131.465 156.850 ;
        RECT 131.635 156.800 131.925 157.525 ;
        RECT 132.145 156.770 132.395 157.525 ;
        RECT 132.565 156.815 132.815 157.345 ;
        RECT 132.985 157.065 133.290 157.525 ;
        RECT 133.535 157.145 134.605 157.315 ;
        RECT 132.565 156.165 132.770 156.815 ;
        RECT 133.535 156.790 133.855 157.145 ;
        RECT 133.530 156.615 133.855 156.790 ;
        RECT 132.940 156.315 133.855 156.615 ;
        RECT 134.025 156.575 134.265 156.975 ;
        RECT 134.435 156.915 134.605 157.145 ;
        RECT 134.775 157.085 134.965 157.525 ;
        RECT 135.135 157.075 136.085 157.355 ;
        RECT 136.305 157.165 136.655 157.335 ;
        RECT 134.435 156.745 134.965 156.915 ;
        RECT 132.940 156.285 133.680 156.315 ;
        RECT 130.345 155.145 130.515 155.905 ;
        RECT 130.695 154.975 131.025 155.735 ;
        RECT 131.195 155.145 131.465 156.050 ;
        RECT 131.635 154.975 131.925 156.140 ;
        RECT 132.145 154.975 132.395 156.115 ;
        RECT 132.565 155.285 132.815 156.165 ;
        RECT 132.985 154.975 133.290 156.115 ;
        RECT 133.510 155.695 133.680 156.285 ;
        RECT 134.025 156.205 134.565 156.575 ;
        RECT 134.745 156.465 134.965 156.745 ;
        RECT 135.135 156.295 135.305 157.075 ;
        RECT 134.900 156.125 135.305 156.295 ;
        RECT 135.475 156.285 135.825 156.905 ;
        RECT 134.900 156.035 135.070 156.125 ;
        RECT 135.995 156.115 136.205 156.905 ;
        RECT 133.850 155.865 135.070 156.035 ;
        RECT 135.530 155.955 136.205 156.115 ;
        RECT 133.510 155.525 134.310 155.695 ;
        RECT 133.630 154.975 133.960 155.355 ;
        RECT 134.140 155.235 134.310 155.525 ;
        RECT 134.900 155.485 135.070 155.865 ;
        RECT 135.240 155.945 136.205 155.955 ;
        RECT 136.395 156.775 136.655 157.165 ;
        RECT 136.865 157.065 137.195 157.525 ;
        RECT 138.070 157.135 138.925 157.305 ;
        RECT 139.130 157.135 139.625 157.305 ;
        RECT 139.795 157.165 140.125 157.525 ;
        RECT 136.395 156.085 136.565 156.775 ;
        RECT 136.735 156.425 136.905 156.605 ;
        RECT 137.075 156.595 137.865 156.845 ;
        RECT 138.070 156.425 138.240 157.135 ;
        RECT 138.410 156.625 138.765 156.845 ;
        RECT 136.735 156.255 138.425 156.425 ;
        RECT 135.240 155.655 135.700 155.945 ;
        RECT 136.395 155.915 137.895 156.085 ;
        RECT 136.395 155.775 136.565 155.915 ;
        RECT 136.005 155.605 136.565 155.775 ;
        RECT 134.480 154.975 134.730 155.435 ;
        RECT 134.900 155.145 135.770 155.485 ;
        RECT 136.005 155.145 136.175 155.605 ;
        RECT 137.010 155.575 138.085 155.745 ;
        RECT 136.345 154.975 136.715 155.435 ;
        RECT 137.010 155.235 137.180 155.575 ;
        RECT 137.350 154.975 137.680 155.405 ;
        RECT 137.915 155.235 138.085 155.575 ;
        RECT 138.255 155.475 138.425 156.255 ;
        RECT 138.595 156.035 138.765 156.625 ;
        RECT 138.935 156.225 139.285 156.845 ;
        RECT 138.595 155.645 139.060 156.035 ;
        RECT 139.455 155.775 139.625 157.135 ;
        RECT 139.795 155.945 140.255 156.995 ;
        RECT 139.230 155.605 139.625 155.775 ;
        RECT 139.230 155.475 139.400 155.605 ;
        RECT 138.255 155.145 138.935 155.475 ;
        RECT 139.150 155.145 139.400 155.475 ;
        RECT 139.570 154.975 139.820 155.435 ;
        RECT 139.990 155.160 140.315 155.945 ;
        RECT 140.485 155.145 140.655 157.265 ;
        RECT 140.825 157.145 141.155 157.525 ;
        RECT 141.325 156.975 141.580 157.265 ;
        RECT 140.830 156.805 141.580 156.975 ;
        RECT 141.760 156.975 142.015 157.265 ;
        RECT 142.185 157.145 142.515 157.525 ;
        RECT 141.760 156.805 142.510 156.975 ;
        RECT 140.830 155.815 141.060 156.805 ;
        RECT 141.230 155.985 141.580 156.635 ;
        RECT 141.760 155.985 142.110 156.635 ;
        RECT 142.280 155.815 142.510 156.805 ;
        RECT 140.830 155.645 141.580 155.815 ;
        RECT 140.825 154.975 141.155 155.475 ;
        RECT 141.325 155.145 141.580 155.645 ;
        RECT 141.760 155.645 142.510 155.815 ;
        RECT 141.760 155.145 142.015 155.645 ;
        RECT 142.185 154.975 142.515 155.475 ;
        RECT 142.685 155.145 142.855 157.265 ;
        RECT 143.215 157.165 143.545 157.525 ;
        RECT 143.715 157.135 144.210 157.305 ;
        RECT 144.415 157.135 145.270 157.305 ;
        RECT 143.085 155.945 143.545 156.995 ;
        RECT 143.025 155.160 143.350 155.945 ;
        RECT 143.715 155.775 143.885 157.135 ;
        RECT 144.055 156.225 144.405 156.845 ;
        RECT 144.575 156.625 144.930 156.845 ;
        RECT 144.575 156.035 144.745 156.625 ;
        RECT 145.100 156.425 145.270 157.135 ;
        RECT 146.145 157.065 146.475 157.525 ;
        RECT 146.685 157.165 147.035 157.335 ;
        RECT 145.475 156.595 146.265 156.845 ;
        RECT 146.685 156.775 146.945 157.165 ;
        RECT 147.255 157.075 148.205 157.355 ;
        RECT 148.375 157.085 148.565 157.525 ;
        RECT 148.735 157.145 149.805 157.315 ;
        RECT 146.435 156.425 146.605 156.605 ;
        RECT 143.715 155.605 144.110 155.775 ;
        RECT 144.280 155.645 144.745 156.035 ;
        RECT 144.915 156.255 146.605 156.425 ;
        RECT 143.940 155.475 144.110 155.605 ;
        RECT 144.915 155.475 145.085 156.255 ;
        RECT 146.775 156.085 146.945 156.775 ;
        RECT 145.445 155.915 146.945 156.085 ;
        RECT 147.135 156.115 147.345 156.905 ;
        RECT 147.515 156.285 147.865 156.905 ;
        RECT 148.035 156.295 148.205 157.075 ;
        RECT 148.735 156.915 148.905 157.145 ;
        RECT 148.375 156.745 148.905 156.915 ;
        RECT 148.375 156.465 148.595 156.745 ;
        RECT 149.075 156.575 149.315 156.975 ;
        RECT 148.035 156.125 148.440 156.295 ;
        RECT 148.775 156.205 149.315 156.575 ;
        RECT 149.485 156.790 149.805 157.145 ;
        RECT 150.050 157.065 150.355 157.525 ;
        RECT 150.525 156.815 150.775 157.345 ;
        RECT 149.485 156.615 149.810 156.790 ;
        RECT 149.485 156.315 150.400 156.615 ;
        RECT 149.660 156.285 150.400 156.315 ;
        RECT 147.135 155.955 147.810 156.115 ;
        RECT 148.270 156.035 148.440 156.125 ;
        RECT 147.135 155.945 148.100 155.955 ;
        RECT 146.775 155.775 146.945 155.915 ;
        RECT 143.520 154.975 143.770 155.435 ;
        RECT 143.940 155.145 144.190 155.475 ;
        RECT 144.405 155.145 145.085 155.475 ;
        RECT 145.255 155.575 146.330 155.745 ;
        RECT 146.775 155.605 147.335 155.775 ;
        RECT 147.640 155.655 148.100 155.945 ;
        RECT 148.270 155.865 149.490 156.035 ;
        RECT 145.255 155.235 145.425 155.575 ;
        RECT 145.660 154.975 145.990 155.405 ;
        RECT 146.160 155.235 146.330 155.575 ;
        RECT 146.625 154.975 146.995 155.435 ;
        RECT 147.165 155.145 147.335 155.605 ;
        RECT 148.270 155.485 148.440 155.865 ;
        RECT 149.660 155.695 149.830 156.285 ;
        RECT 150.570 156.165 150.775 156.815 ;
        RECT 150.945 156.770 151.195 157.525 ;
        RECT 151.415 156.980 156.760 157.525 ;
        RECT 147.570 155.145 148.440 155.485 ;
        RECT 149.030 155.525 149.830 155.695 ;
        RECT 148.610 154.975 148.860 155.435 ;
        RECT 149.030 155.235 149.200 155.525 ;
        RECT 149.380 154.975 149.710 155.355 ;
        RECT 150.050 154.975 150.355 156.115 ;
        RECT 150.525 155.285 150.775 156.165 ;
        RECT 153.000 156.150 153.340 156.980 ;
        RECT 156.935 156.775 158.145 157.525 ;
        RECT 150.945 154.975 151.195 156.115 ;
        RECT 154.820 155.410 155.170 156.660 ;
        RECT 156.935 156.065 157.455 156.605 ;
        RECT 157.625 156.235 158.145 156.775 ;
        RECT 151.415 154.975 156.760 155.410 ;
        RECT 156.935 154.975 158.145 156.065 ;
        RECT 2.750 154.805 158.230 154.975 ;
        RECT 2.835 153.715 4.045 154.805 ;
        RECT 4.220 154.135 4.475 154.635 ;
        RECT 4.645 154.305 4.975 154.805 ;
        RECT 4.220 153.965 4.970 154.135 ;
        RECT 2.835 153.005 3.355 153.545 ;
        RECT 3.525 153.175 4.045 153.715 ;
        RECT 4.220 153.145 4.570 153.795 ;
        RECT 2.835 152.255 4.045 153.005 ;
        RECT 4.740 152.975 4.970 153.965 ;
        RECT 4.220 152.805 4.970 152.975 ;
        RECT 4.220 152.515 4.475 152.805 ;
        RECT 4.645 152.255 4.975 152.635 ;
        RECT 5.145 152.515 5.315 154.635 ;
        RECT 5.485 153.835 5.810 154.620 ;
        RECT 5.980 154.345 6.230 154.805 ;
        RECT 6.400 154.305 6.650 154.635 ;
        RECT 6.865 154.305 7.545 154.635 ;
        RECT 6.400 154.175 6.570 154.305 ;
        RECT 6.175 154.005 6.570 154.175 ;
        RECT 5.545 152.785 6.005 153.835 ;
        RECT 6.175 152.645 6.345 154.005 ;
        RECT 6.740 153.745 7.205 154.135 ;
        RECT 6.515 152.935 6.865 153.555 ;
        RECT 7.035 153.155 7.205 153.745 ;
        RECT 7.375 153.525 7.545 154.305 ;
        RECT 7.715 154.205 7.885 154.545 ;
        RECT 8.120 154.375 8.450 154.805 ;
        RECT 8.620 154.205 8.790 154.545 ;
        RECT 9.085 154.345 9.455 154.805 ;
        RECT 7.715 154.035 8.790 154.205 ;
        RECT 9.625 154.175 9.795 154.635 ;
        RECT 10.030 154.295 10.900 154.635 ;
        RECT 11.070 154.345 11.320 154.805 ;
        RECT 9.235 154.005 9.795 154.175 ;
        RECT 9.235 153.865 9.405 154.005 ;
        RECT 7.905 153.695 9.405 153.865 ;
        RECT 10.100 153.835 10.560 154.125 ;
        RECT 7.375 153.355 9.065 153.525 ;
        RECT 7.035 152.935 7.390 153.155 ;
        RECT 7.560 152.645 7.730 153.355 ;
        RECT 7.935 152.935 8.725 153.185 ;
        RECT 8.895 153.175 9.065 153.355 ;
        RECT 9.235 153.005 9.405 153.695 ;
        RECT 5.675 152.255 6.005 152.615 ;
        RECT 6.175 152.475 6.670 152.645 ;
        RECT 6.875 152.475 7.730 152.645 ;
        RECT 8.605 152.255 8.935 152.715 ;
        RECT 9.145 152.615 9.405 153.005 ;
        RECT 9.595 153.825 10.560 153.835 ;
        RECT 10.730 153.915 10.900 154.295 ;
        RECT 11.490 154.255 11.660 154.545 ;
        RECT 11.840 154.425 12.170 154.805 ;
        RECT 11.490 154.085 12.290 154.255 ;
        RECT 9.595 153.665 10.270 153.825 ;
        RECT 10.730 153.745 11.950 153.915 ;
        RECT 9.595 152.875 9.805 153.665 ;
        RECT 10.730 153.655 10.900 153.745 ;
        RECT 9.975 152.875 10.325 153.495 ;
        RECT 10.495 153.485 10.900 153.655 ;
        RECT 10.495 152.705 10.665 153.485 ;
        RECT 10.835 153.035 11.055 153.315 ;
        RECT 11.235 153.205 11.775 153.575 ;
        RECT 12.120 153.495 12.290 154.085 ;
        RECT 12.510 153.665 12.815 154.805 ;
        RECT 12.985 153.615 13.240 154.495 ;
        RECT 12.120 153.465 12.860 153.495 ;
        RECT 10.835 152.865 11.365 153.035 ;
        RECT 9.145 152.445 9.495 152.615 ;
        RECT 9.715 152.425 10.665 152.705 ;
        RECT 10.835 152.255 11.025 152.695 ;
        RECT 11.195 152.635 11.365 152.865 ;
        RECT 11.535 152.805 11.775 153.205 ;
        RECT 11.945 153.165 12.860 153.465 ;
        RECT 11.945 152.990 12.270 153.165 ;
        RECT 11.945 152.635 12.265 152.990 ;
        RECT 13.030 152.965 13.240 153.615 ;
        RECT 11.195 152.465 12.265 152.635 ;
        RECT 12.510 152.255 12.815 152.715 ;
        RECT 12.985 152.435 13.240 152.965 ;
        RECT 13.415 153.730 13.685 154.635 ;
        RECT 13.855 154.045 14.185 154.805 ;
        RECT 14.365 153.875 14.535 154.635 ;
        RECT 13.415 152.930 13.585 153.730 ;
        RECT 13.870 153.705 14.535 153.875 ;
        RECT 13.870 153.560 14.040 153.705 ;
        RECT 15.715 153.640 16.005 154.805 ;
        RECT 16.180 153.665 16.515 154.635 ;
        RECT 16.685 153.665 16.855 154.805 ;
        RECT 17.025 154.465 19.055 154.635 ;
        RECT 13.755 153.230 14.040 153.560 ;
        RECT 13.870 152.975 14.040 153.230 ;
        RECT 14.275 153.155 14.605 153.525 ;
        RECT 16.180 152.995 16.350 153.665 ;
        RECT 17.025 153.495 17.195 154.465 ;
        RECT 16.520 153.165 16.775 153.495 ;
        RECT 17.000 153.165 17.195 153.495 ;
        RECT 17.365 154.125 18.490 154.295 ;
        RECT 16.605 152.995 16.775 153.165 ;
        RECT 17.365 152.995 17.535 154.125 ;
        RECT 13.415 152.425 13.675 152.930 ;
        RECT 13.870 152.805 14.535 152.975 ;
        RECT 13.855 152.255 14.185 152.635 ;
        RECT 14.365 152.425 14.535 152.805 ;
        RECT 15.715 152.255 16.005 152.980 ;
        RECT 16.180 152.425 16.435 152.995 ;
        RECT 16.605 152.825 17.535 152.995 ;
        RECT 17.705 153.785 18.715 153.955 ;
        RECT 17.705 152.985 17.875 153.785 ;
        RECT 18.080 153.445 18.355 153.585 ;
        RECT 18.075 153.275 18.355 153.445 ;
        RECT 17.360 152.790 17.535 152.825 ;
        RECT 16.605 152.255 16.935 152.655 ;
        RECT 17.360 152.425 17.890 152.790 ;
        RECT 18.080 152.425 18.355 153.275 ;
        RECT 18.525 152.425 18.715 153.785 ;
        RECT 18.885 153.800 19.055 154.465 ;
        RECT 19.225 154.045 19.395 154.805 ;
        RECT 19.630 154.045 20.145 154.455 ;
        RECT 18.885 153.610 19.635 153.800 ;
        RECT 19.805 153.235 20.145 154.045 ;
        RECT 20.320 154.415 20.655 154.635 ;
        RECT 21.660 154.425 22.015 154.805 ;
        RECT 20.320 153.795 20.575 154.415 ;
        RECT 20.825 154.255 21.055 154.295 ;
        RECT 22.185 154.255 22.435 154.635 ;
        RECT 20.825 154.055 22.435 154.255 ;
        RECT 20.825 153.965 21.010 154.055 ;
        RECT 21.600 154.045 22.435 154.055 ;
        RECT 22.685 154.025 22.935 154.805 ;
        RECT 23.105 153.955 23.365 154.635 ;
        RECT 24.000 154.135 24.255 154.635 ;
        RECT 24.425 154.305 24.755 154.805 ;
        RECT 24.000 153.965 24.750 154.135 ;
        RECT 21.165 153.855 21.495 153.885 ;
        RECT 21.165 153.795 22.965 153.855 ;
        RECT 20.320 153.685 23.025 153.795 ;
        RECT 20.320 153.625 21.495 153.685 ;
        RECT 22.825 153.650 23.025 153.685 ;
        RECT 20.315 153.245 20.805 153.445 ;
        RECT 20.995 153.245 21.470 153.455 ;
        RECT 18.915 153.065 20.145 153.235 ;
        RECT 18.895 152.255 19.405 152.790 ;
        RECT 19.625 152.460 19.870 153.065 ;
        RECT 20.320 152.255 20.775 153.020 ;
        RECT 21.250 152.845 21.470 153.245 ;
        RECT 21.715 153.245 22.045 153.455 ;
        RECT 21.715 152.845 21.925 153.245 ;
        RECT 22.215 153.210 22.625 153.515 ;
        RECT 22.855 153.075 23.025 153.650 ;
        RECT 22.755 152.955 23.025 153.075 ;
        RECT 22.180 152.910 23.025 152.955 ;
        RECT 22.180 152.785 22.935 152.910 ;
        RECT 22.180 152.635 22.350 152.785 ;
        RECT 23.195 152.765 23.365 153.955 ;
        RECT 24.000 153.145 24.350 153.795 ;
        RECT 24.520 152.975 24.750 153.965 ;
        RECT 23.135 152.755 23.365 152.765 ;
        RECT 21.050 152.425 22.350 152.635 ;
        RECT 22.605 152.255 22.935 152.615 ;
        RECT 23.105 152.425 23.365 152.755 ;
        RECT 24.000 152.805 24.750 152.975 ;
        RECT 24.000 152.515 24.255 152.805 ;
        RECT 24.425 152.255 24.755 152.635 ;
        RECT 24.925 152.515 25.095 154.635 ;
        RECT 25.265 153.835 25.590 154.620 ;
        RECT 25.760 154.345 26.010 154.805 ;
        RECT 26.180 154.305 26.430 154.635 ;
        RECT 26.645 154.305 27.325 154.635 ;
        RECT 26.180 154.175 26.350 154.305 ;
        RECT 25.955 154.005 26.350 154.175 ;
        RECT 25.325 152.785 25.785 153.835 ;
        RECT 25.955 152.645 26.125 154.005 ;
        RECT 26.520 153.745 26.985 154.135 ;
        RECT 26.295 152.935 26.645 153.555 ;
        RECT 26.815 153.155 26.985 153.745 ;
        RECT 27.155 153.525 27.325 154.305 ;
        RECT 27.495 154.205 27.665 154.545 ;
        RECT 27.900 154.375 28.230 154.805 ;
        RECT 28.400 154.205 28.570 154.545 ;
        RECT 28.865 154.345 29.235 154.805 ;
        RECT 27.495 154.035 28.570 154.205 ;
        RECT 29.405 154.175 29.575 154.635 ;
        RECT 29.810 154.295 30.680 154.635 ;
        RECT 30.850 154.345 31.100 154.805 ;
        RECT 29.015 154.005 29.575 154.175 ;
        RECT 29.015 153.865 29.185 154.005 ;
        RECT 27.685 153.695 29.185 153.865 ;
        RECT 29.880 153.835 30.340 154.125 ;
        RECT 27.155 153.355 28.845 153.525 ;
        RECT 26.815 152.935 27.170 153.155 ;
        RECT 27.340 152.645 27.510 153.355 ;
        RECT 27.715 152.935 28.505 153.185 ;
        RECT 28.675 153.175 28.845 153.355 ;
        RECT 29.015 153.005 29.185 153.695 ;
        RECT 25.455 152.255 25.785 152.615 ;
        RECT 25.955 152.475 26.450 152.645 ;
        RECT 26.655 152.475 27.510 152.645 ;
        RECT 28.385 152.255 28.715 152.715 ;
        RECT 28.925 152.615 29.185 153.005 ;
        RECT 29.375 153.825 30.340 153.835 ;
        RECT 30.510 153.915 30.680 154.295 ;
        RECT 31.270 154.255 31.440 154.545 ;
        RECT 31.620 154.425 31.950 154.805 ;
        RECT 31.270 154.085 32.070 154.255 ;
        RECT 29.375 153.665 30.050 153.825 ;
        RECT 30.510 153.745 31.730 153.915 ;
        RECT 29.375 152.875 29.585 153.665 ;
        RECT 30.510 153.655 30.680 153.745 ;
        RECT 29.755 152.875 30.105 153.495 ;
        RECT 30.275 153.485 30.680 153.655 ;
        RECT 30.275 152.705 30.445 153.485 ;
        RECT 30.615 153.035 30.835 153.315 ;
        RECT 31.015 153.205 31.555 153.575 ;
        RECT 31.900 153.495 32.070 154.085 ;
        RECT 32.290 153.665 32.595 154.805 ;
        RECT 32.765 153.615 33.020 154.495 ;
        RECT 31.900 153.465 32.640 153.495 ;
        RECT 30.615 152.865 31.145 153.035 ;
        RECT 28.925 152.445 29.275 152.615 ;
        RECT 29.495 152.425 30.445 152.705 ;
        RECT 30.615 152.255 30.805 152.695 ;
        RECT 30.975 152.635 31.145 152.865 ;
        RECT 31.315 152.805 31.555 153.205 ;
        RECT 31.725 153.165 32.640 153.465 ;
        RECT 31.725 152.990 32.050 153.165 ;
        RECT 31.725 152.635 32.045 152.990 ;
        RECT 32.810 152.965 33.020 153.615 ;
        RECT 30.975 152.465 32.045 152.635 ;
        RECT 32.290 152.255 32.595 152.715 ;
        RECT 32.765 152.435 33.020 152.965 ;
        RECT 33.195 153.665 33.580 154.635 ;
        RECT 33.750 154.345 34.075 154.805 ;
        RECT 34.595 154.175 34.875 154.635 ;
        RECT 33.750 153.955 34.875 154.175 ;
        RECT 33.195 152.995 33.475 153.665 ;
        RECT 33.750 153.495 34.200 153.955 ;
        RECT 35.065 153.785 35.465 154.635 ;
        RECT 35.865 154.345 36.135 154.805 ;
        RECT 36.305 154.175 36.590 154.635 ;
        RECT 33.645 153.165 34.200 153.495 ;
        RECT 34.370 153.225 35.465 153.785 ;
        RECT 33.750 153.055 34.200 153.165 ;
        RECT 33.195 152.425 33.580 152.995 ;
        RECT 33.750 152.885 34.875 153.055 ;
        RECT 33.750 152.255 34.075 152.715 ;
        RECT 34.595 152.425 34.875 152.885 ;
        RECT 35.065 152.425 35.465 153.225 ;
        RECT 35.635 153.955 36.590 154.175 ;
        RECT 35.635 153.055 35.845 153.955 ;
        RECT 36.015 153.225 36.705 153.785 ;
        RECT 36.875 153.745 37.190 154.805 ;
        RECT 37.820 154.300 38.435 154.805 ;
        RECT 35.635 152.885 36.590 153.055 ;
        RECT 36.935 152.915 37.200 153.495 ;
        RECT 37.370 153.415 37.645 154.075 ;
        RECT 37.840 153.765 38.075 154.130 ;
        RECT 38.245 154.125 38.435 154.300 ;
        RECT 38.605 154.295 39.080 154.635 ;
        RECT 38.245 153.935 38.575 154.125 ;
        RECT 38.800 153.765 38.990 154.060 ;
        RECT 39.250 153.960 39.465 154.805 ;
        RECT 39.665 153.965 39.950 154.635 ;
        RECT 37.840 153.595 39.610 153.765 ;
        RECT 37.370 153.185 38.205 153.415 ;
        RECT 35.865 152.255 36.135 152.715 ;
        RECT 36.305 152.425 36.590 152.885 ;
        RECT 36.875 152.255 37.145 152.745 ;
        RECT 37.370 152.475 37.645 153.185 ;
        RECT 38.375 152.740 38.630 153.595 ;
        RECT 37.845 152.475 38.630 152.740 ;
        RECT 38.800 152.935 39.210 153.415 ;
        RECT 39.380 153.165 39.610 153.595 ;
        RECT 39.780 153.615 39.950 153.965 ;
        RECT 40.120 153.795 40.385 154.805 ;
        RECT 41.475 153.640 41.765 154.805 ;
        RECT 41.935 153.795 42.200 154.805 ;
        RECT 42.370 153.965 42.655 154.635 ;
        RECT 42.370 153.955 42.625 153.965 ;
        RECT 42.855 153.960 43.070 154.805 ;
        RECT 43.240 154.295 43.715 154.635 ;
        RECT 43.885 154.300 44.500 154.805 ;
        RECT 43.885 154.125 44.075 154.300 ;
        RECT 42.370 153.615 42.540 153.955 ;
        RECT 43.330 153.765 43.520 154.060 ;
        RECT 43.745 153.935 44.075 154.125 ;
        RECT 44.245 153.765 44.480 154.130 ;
        RECT 39.780 153.095 40.385 153.615 ;
        RECT 41.935 153.095 42.540 153.615 ;
        RECT 42.710 153.595 44.480 153.765 ;
        RECT 42.710 153.165 42.940 153.595 ;
        RECT 38.800 152.475 39.010 152.935 ;
        RECT 39.780 152.885 39.950 153.095 ;
        RECT 39.200 152.255 39.530 152.750 ;
        RECT 39.705 152.425 39.950 152.885 ;
        RECT 40.120 152.255 40.385 152.915 ;
        RECT 41.475 152.255 41.765 152.980 ;
        RECT 41.935 152.255 42.200 152.915 ;
        RECT 42.370 152.885 42.540 153.095 ;
        RECT 43.110 152.935 43.520 153.415 ;
        RECT 42.370 152.425 42.615 152.885 ;
        RECT 42.790 152.255 43.120 152.750 ;
        RECT 43.310 152.475 43.520 152.935 ;
        RECT 43.690 152.740 43.945 153.595 ;
        RECT 44.675 153.415 44.950 154.075 ;
        RECT 45.130 153.745 45.445 154.805 ;
        RECT 45.705 153.875 45.875 154.635 ;
        RECT 46.055 154.045 46.385 154.805 ;
        RECT 45.705 153.705 46.370 153.875 ;
        RECT 46.555 153.730 46.825 154.635 ;
        RECT 46.200 153.560 46.370 153.705 ;
        RECT 44.115 153.185 44.950 153.415 ;
        RECT 43.690 152.475 44.475 152.740 ;
        RECT 44.675 152.475 44.950 153.185 ;
        RECT 45.120 152.915 45.385 153.495 ;
        RECT 45.635 153.155 45.965 153.525 ;
        RECT 46.200 153.230 46.485 153.560 ;
        RECT 46.200 152.975 46.370 153.230 ;
        RECT 45.705 152.805 46.370 152.975 ;
        RECT 46.655 152.930 46.825 153.730 ;
        RECT 45.175 152.255 45.445 152.745 ;
        RECT 45.705 152.425 45.875 152.805 ;
        RECT 46.055 152.255 46.385 152.635 ;
        RECT 46.565 152.425 46.825 152.930 ;
        RECT 46.995 153.665 47.270 154.635 ;
        RECT 47.480 154.005 47.760 154.805 ;
        RECT 47.930 154.295 49.545 154.625 ;
        RECT 47.930 153.955 49.105 154.125 ;
        RECT 47.930 153.835 48.100 153.955 ;
        RECT 47.440 153.665 48.100 153.835 ;
        RECT 46.995 152.930 47.165 153.665 ;
        RECT 47.440 153.495 47.610 153.665 ;
        RECT 48.360 153.495 48.605 153.785 ;
        RECT 48.775 153.665 49.105 153.955 ;
        RECT 49.365 153.495 49.535 154.055 ;
        RECT 49.785 153.665 50.045 154.805 ;
        RECT 51.335 153.965 51.585 154.805 ;
        RECT 51.755 153.795 52.005 154.635 ;
        RECT 52.175 153.965 52.425 154.805 ;
        RECT 52.595 153.795 52.845 154.635 ;
        RECT 53.055 154.005 53.755 154.805 ;
        RECT 53.925 154.465 55.105 154.635 ;
        RECT 53.925 153.835 54.190 154.465 ;
        RECT 51.135 153.625 52.845 153.795 ;
        RECT 53.100 153.665 54.190 153.835 ;
        RECT 47.335 153.165 47.610 153.495 ;
        RECT 47.780 153.165 48.605 153.495 ;
        RECT 48.820 153.165 49.535 153.495 ;
        RECT 49.705 153.245 50.040 153.495 ;
        RECT 47.440 152.995 47.610 153.165 ;
        RECT 49.285 153.075 49.535 153.165 ;
        RECT 51.135 153.075 51.425 153.625 ;
        RECT 53.100 153.415 53.320 153.665 ;
        RECT 54.360 153.495 54.595 154.220 ;
        RECT 54.765 153.665 55.105 154.465 ;
        RECT 55.280 154.135 55.535 154.635 ;
        RECT 55.705 154.305 56.035 154.805 ;
        RECT 55.280 153.965 56.030 154.135 ;
        RECT 51.595 153.245 53.320 153.415 ;
        RECT 53.490 153.245 53.965 153.495 ;
        RECT 54.135 153.245 54.595 153.495 ;
        RECT 54.765 153.245 55.105 153.495 ;
        RECT 53.100 153.075 53.320 153.245 ;
        RECT 55.280 153.145 55.630 153.795 ;
        RECT 46.995 152.585 47.270 152.930 ;
        RECT 47.440 152.825 49.105 152.995 ;
        RECT 47.460 152.255 47.835 152.655 ;
        RECT 48.005 152.475 48.175 152.825 ;
        RECT 48.345 152.255 48.675 152.655 ;
        RECT 48.845 152.425 49.105 152.825 ;
        RECT 49.285 152.655 49.615 153.075 ;
        RECT 49.785 152.255 50.045 153.075 ;
        RECT 51.135 152.905 52.885 153.075 ;
        RECT 51.375 152.255 51.545 152.725 ;
        RECT 51.715 152.435 52.045 152.905 ;
        RECT 52.215 152.255 52.385 152.725 ;
        RECT 52.555 152.435 52.885 152.905 ;
        RECT 53.100 152.895 55.105 153.075 ;
        RECT 55.800 152.975 56.030 153.965 ;
        RECT 53.055 152.255 53.755 152.725 ;
        RECT 53.925 152.425 54.255 152.895 ;
        RECT 54.425 152.255 54.595 152.725 ;
        RECT 54.765 152.425 55.105 152.895 ;
        RECT 55.280 152.805 56.030 152.975 ;
        RECT 55.280 152.515 55.535 152.805 ;
        RECT 55.705 152.255 56.035 152.635 ;
        RECT 56.205 152.515 56.375 154.635 ;
        RECT 56.545 153.835 56.870 154.620 ;
        RECT 57.040 154.345 57.290 154.805 ;
        RECT 57.460 154.305 57.710 154.635 ;
        RECT 57.925 154.305 58.605 154.635 ;
        RECT 57.460 154.175 57.630 154.305 ;
        RECT 57.235 154.005 57.630 154.175 ;
        RECT 56.605 152.785 57.065 153.835 ;
        RECT 57.235 152.645 57.405 154.005 ;
        RECT 57.800 153.745 58.265 154.135 ;
        RECT 57.575 152.935 57.925 153.555 ;
        RECT 58.095 153.155 58.265 153.745 ;
        RECT 58.435 153.525 58.605 154.305 ;
        RECT 58.775 154.205 58.945 154.545 ;
        RECT 59.180 154.375 59.510 154.805 ;
        RECT 59.680 154.205 59.850 154.545 ;
        RECT 60.145 154.345 60.515 154.805 ;
        RECT 58.775 154.035 59.850 154.205 ;
        RECT 60.685 154.175 60.855 154.635 ;
        RECT 61.090 154.295 61.960 154.635 ;
        RECT 62.130 154.345 62.380 154.805 ;
        RECT 60.295 154.005 60.855 154.175 ;
        RECT 60.295 153.865 60.465 154.005 ;
        RECT 58.965 153.695 60.465 153.865 ;
        RECT 61.160 153.835 61.620 154.125 ;
        RECT 58.435 153.355 60.125 153.525 ;
        RECT 58.095 152.935 58.450 153.155 ;
        RECT 58.620 152.645 58.790 153.355 ;
        RECT 58.995 152.935 59.785 153.185 ;
        RECT 59.955 153.175 60.125 153.355 ;
        RECT 60.295 153.005 60.465 153.695 ;
        RECT 56.735 152.255 57.065 152.615 ;
        RECT 57.235 152.475 57.730 152.645 ;
        RECT 57.935 152.475 58.790 152.645 ;
        RECT 59.665 152.255 59.995 152.715 ;
        RECT 60.205 152.615 60.465 153.005 ;
        RECT 60.655 153.825 61.620 153.835 ;
        RECT 61.790 153.915 61.960 154.295 ;
        RECT 62.550 154.255 62.720 154.545 ;
        RECT 62.900 154.425 63.230 154.805 ;
        RECT 62.550 154.085 63.350 154.255 ;
        RECT 60.655 153.665 61.330 153.825 ;
        RECT 61.790 153.745 63.010 153.915 ;
        RECT 60.655 152.875 60.865 153.665 ;
        RECT 61.790 153.655 61.960 153.745 ;
        RECT 61.035 152.875 61.385 153.495 ;
        RECT 61.555 153.485 61.960 153.655 ;
        RECT 61.555 152.705 61.725 153.485 ;
        RECT 61.895 153.035 62.115 153.315 ;
        RECT 62.295 153.205 62.835 153.575 ;
        RECT 63.180 153.495 63.350 154.085 ;
        RECT 63.570 153.665 63.875 154.805 ;
        RECT 64.045 153.615 64.300 154.495 ;
        RECT 64.480 154.295 66.135 154.585 ;
        RECT 64.480 153.955 66.070 154.125 ;
        RECT 66.305 154.005 66.585 154.805 ;
        RECT 64.480 153.665 64.800 153.955 ;
        RECT 65.900 153.835 66.070 153.955 ;
        RECT 64.995 153.615 65.710 153.785 ;
        RECT 65.900 153.665 66.625 153.835 ;
        RECT 66.795 153.665 67.065 154.635 ;
        RECT 63.180 153.465 63.920 153.495 ;
        RECT 61.895 152.865 62.425 153.035 ;
        RECT 60.205 152.445 60.555 152.615 ;
        RECT 60.775 152.425 61.725 152.705 ;
        RECT 61.895 152.255 62.085 152.695 ;
        RECT 62.255 152.635 62.425 152.865 ;
        RECT 62.595 152.805 62.835 153.205 ;
        RECT 63.005 153.165 63.920 153.465 ;
        RECT 63.005 152.990 63.330 153.165 ;
        RECT 63.005 152.635 63.325 152.990 ;
        RECT 64.090 152.965 64.300 153.615 ;
        RECT 62.255 152.465 63.325 152.635 ;
        RECT 63.570 152.255 63.875 152.715 ;
        RECT 64.045 152.435 64.300 152.965 ;
        RECT 64.480 152.925 64.830 153.495 ;
        RECT 65.000 153.165 65.710 153.615 ;
        RECT 66.455 153.495 66.625 153.665 ;
        RECT 65.880 153.165 66.285 153.495 ;
        RECT 66.455 153.165 66.725 153.495 ;
        RECT 66.455 152.995 66.625 153.165 ;
        RECT 65.015 152.825 66.625 152.995 ;
        RECT 66.895 152.930 67.065 153.665 ;
        RECT 67.235 153.640 67.525 154.805 ;
        RECT 67.700 153.665 68.035 154.635 ;
        RECT 68.205 153.665 68.375 154.805 ;
        RECT 68.545 154.465 70.575 154.635 ;
        RECT 67.700 152.995 67.870 153.665 ;
        RECT 68.545 153.495 68.715 154.465 ;
        RECT 68.040 153.165 68.295 153.495 ;
        RECT 68.520 153.165 68.715 153.495 ;
        RECT 68.885 154.125 70.010 154.295 ;
        RECT 68.125 152.995 68.295 153.165 ;
        RECT 68.885 152.995 69.055 154.125 ;
        RECT 64.485 152.255 64.815 152.755 ;
        RECT 65.015 152.475 65.185 152.825 ;
        RECT 65.385 152.255 65.715 152.655 ;
        RECT 65.885 152.475 66.055 152.825 ;
        RECT 66.225 152.255 66.605 152.655 ;
        RECT 66.795 152.585 67.065 152.930 ;
        RECT 67.235 152.255 67.525 152.980 ;
        RECT 67.700 152.425 67.955 152.995 ;
        RECT 68.125 152.825 69.055 152.995 ;
        RECT 69.225 153.785 70.235 153.955 ;
        RECT 69.225 152.985 69.395 153.785 ;
        RECT 68.880 152.790 69.055 152.825 ;
        RECT 68.125 152.255 68.455 152.655 ;
        RECT 68.880 152.425 69.410 152.790 ;
        RECT 69.600 152.765 69.875 153.585 ;
        RECT 69.595 152.595 69.875 152.765 ;
        RECT 69.600 152.425 69.875 152.595 ;
        RECT 70.045 152.425 70.235 153.785 ;
        RECT 70.405 153.800 70.575 154.465 ;
        RECT 70.745 154.045 70.915 154.805 ;
        RECT 71.150 154.045 71.665 154.455 ;
        RECT 70.405 153.610 71.155 153.800 ;
        RECT 71.325 153.235 71.665 154.045 ;
        RECT 70.435 153.065 71.665 153.235 ;
        RECT 71.835 153.665 72.220 154.635 ;
        RECT 72.390 154.345 72.715 154.805 ;
        RECT 73.235 154.175 73.515 154.635 ;
        RECT 72.390 153.955 73.515 154.175 ;
        RECT 70.415 152.255 70.925 152.790 ;
        RECT 71.145 152.460 71.390 153.065 ;
        RECT 71.835 152.995 72.115 153.665 ;
        RECT 72.390 153.495 72.840 153.955 ;
        RECT 73.705 153.785 74.105 154.635 ;
        RECT 74.505 154.345 74.775 154.805 ;
        RECT 74.945 154.175 75.230 154.635 ;
        RECT 72.285 153.165 72.840 153.495 ;
        RECT 73.010 153.225 74.105 153.785 ;
        RECT 72.390 153.055 72.840 153.165 ;
        RECT 71.835 152.425 72.220 152.995 ;
        RECT 72.390 152.885 73.515 153.055 ;
        RECT 72.390 152.255 72.715 152.715 ;
        RECT 73.235 152.425 73.515 152.885 ;
        RECT 73.705 152.425 74.105 153.225 ;
        RECT 74.275 153.955 75.230 154.175 ;
        RECT 74.275 153.055 74.485 153.955 ;
        RECT 75.570 153.935 75.855 154.805 ;
        RECT 76.025 154.175 76.285 154.635 ;
        RECT 76.460 154.345 76.715 154.805 ;
        RECT 76.885 154.175 77.145 154.635 ;
        RECT 76.025 154.005 77.145 154.175 ;
        RECT 77.315 154.005 77.625 154.805 ;
        RECT 74.655 153.225 75.345 153.785 ;
        RECT 76.025 153.755 76.285 154.005 ;
        RECT 77.795 153.835 78.105 154.635 ;
        RECT 78.275 154.295 79.465 154.585 ;
        RECT 75.530 153.585 76.285 153.755 ;
        RECT 77.075 153.665 78.105 153.835 ;
        RECT 78.295 153.955 79.465 154.125 ;
        RECT 79.635 154.005 79.915 154.805 ;
        RECT 78.295 153.665 78.620 153.955 ;
        RECT 79.295 153.835 79.465 153.955 ;
        RECT 75.530 153.075 75.935 153.585 ;
        RECT 77.075 153.415 77.245 153.665 ;
        RECT 76.105 153.245 77.245 153.415 ;
        RECT 74.275 152.885 75.230 153.055 ;
        RECT 75.530 152.905 77.180 153.075 ;
        RECT 77.415 152.925 77.765 153.495 ;
        RECT 74.505 152.255 74.775 152.715 ;
        RECT 74.945 152.425 75.230 152.885 ;
        RECT 75.575 152.255 75.855 152.735 ;
        RECT 76.025 152.515 76.285 152.905 ;
        RECT 76.460 152.255 76.715 152.735 ;
        RECT 76.885 152.515 77.180 152.905 ;
        RECT 77.935 152.755 78.105 153.665 ;
        RECT 78.790 153.495 78.985 153.785 ;
        RECT 79.295 153.665 79.955 153.835 ;
        RECT 80.125 153.665 80.400 154.635 ;
        RECT 79.785 153.495 79.955 153.665 ;
        RECT 78.275 153.165 78.620 153.495 ;
        RECT 78.790 153.165 79.615 153.495 ;
        RECT 79.785 153.165 80.060 153.495 ;
        RECT 79.785 152.995 79.955 153.165 ;
        RECT 77.360 152.255 77.635 152.735 ;
        RECT 77.805 152.425 78.105 152.755 ;
        RECT 78.290 152.825 79.955 152.995 ;
        RECT 80.230 152.930 80.400 153.665 ;
        RECT 78.290 152.475 78.545 152.825 ;
        RECT 78.715 152.255 79.045 152.655 ;
        RECT 79.215 152.475 79.385 152.825 ;
        RECT 79.555 152.255 79.935 152.655 ;
        RECT 80.125 152.585 80.400 152.930 ;
        RECT 80.580 153.665 80.855 154.635 ;
        RECT 81.065 154.005 81.345 154.805 ;
        RECT 81.515 154.295 82.705 154.585 ;
        RECT 81.515 153.955 82.685 154.125 ;
        RECT 81.515 153.835 81.685 153.955 ;
        RECT 81.025 153.665 81.685 153.835 ;
        RECT 80.580 152.930 80.750 153.665 ;
        RECT 81.025 153.495 81.195 153.665 ;
        RECT 81.995 153.495 82.190 153.785 ;
        RECT 82.360 153.665 82.685 153.955 ;
        RECT 83.335 154.045 83.850 154.455 ;
        RECT 84.085 154.045 84.255 154.805 ;
        RECT 84.425 154.465 86.455 154.635 ;
        RECT 80.920 153.165 81.195 153.495 ;
        RECT 81.365 153.165 82.190 153.495 ;
        RECT 82.360 153.165 82.705 153.495 ;
        RECT 83.335 153.235 83.675 154.045 ;
        RECT 84.425 153.800 84.595 154.465 ;
        RECT 84.990 154.125 86.115 154.295 ;
        RECT 83.845 153.610 84.595 153.800 ;
        RECT 84.765 153.785 85.775 153.955 ;
        RECT 81.025 152.995 81.195 153.165 ;
        RECT 83.335 153.065 84.565 153.235 ;
        RECT 80.580 152.585 80.855 152.930 ;
        RECT 81.025 152.825 82.690 152.995 ;
        RECT 81.045 152.255 81.425 152.655 ;
        RECT 81.595 152.475 81.765 152.825 ;
        RECT 81.935 152.255 82.265 152.655 ;
        RECT 82.435 152.475 82.690 152.825 ;
        RECT 83.610 152.460 83.855 153.065 ;
        RECT 84.075 152.255 84.585 152.790 ;
        RECT 84.765 152.425 84.955 153.785 ;
        RECT 85.125 153.445 85.400 153.585 ;
        RECT 85.125 153.275 85.405 153.445 ;
        RECT 85.125 152.425 85.400 153.275 ;
        RECT 85.605 152.985 85.775 153.785 ;
        RECT 85.945 152.995 86.115 154.125 ;
        RECT 86.285 153.495 86.455 154.465 ;
        RECT 86.625 153.665 86.795 154.805 ;
        RECT 86.965 153.665 87.300 154.635 ;
        RECT 87.475 153.715 88.685 154.805 ;
        RECT 86.285 153.165 86.480 153.495 ;
        RECT 86.705 153.165 86.960 153.495 ;
        RECT 86.705 152.995 86.875 153.165 ;
        RECT 87.130 152.995 87.300 153.665 ;
        RECT 85.945 152.825 86.875 152.995 ;
        RECT 85.945 152.790 86.120 152.825 ;
        RECT 85.590 152.425 86.120 152.790 ;
        RECT 86.545 152.255 86.875 152.655 ;
        RECT 87.045 152.425 87.300 152.995 ;
        RECT 87.475 153.005 87.995 153.545 ;
        RECT 88.165 153.175 88.685 153.715 ;
        RECT 88.860 153.665 89.195 154.635 ;
        RECT 89.365 153.665 89.535 154.805 ;
        RECT 89.705 154.465 91.735 154.635 ;
        RECT 87.475 152.255 88.685 153.005 ;
        RECT 88.860 152.995 89.030 153.665 ;
        RECT 89.705 153.495 89.875 154.465 ;
        RECT 89.200 153.165 89.455 153.495 ;
        RECT 89.680 153.165 89.875 153.495 ;
        RECT 90.045 154.125 91.170 154.295 ;
        RECT 89.285 152.995 89.455 153.165 ;
        RECT 90.045 152.995 90.215 154.125 ;
        RECT 88.860 152.425 89.115 152.995 ;
        RECT 89.285 152.825 90.215 152.995 ;
        RECT 90.385 153.785 91.395 153.955 ;
        RECT 90.385 152.985 90.555 153.785 ;
        RECT 90.760 153.105 91.035 153.585 ;
        RECT 90.755 152.935 91.035 153.105 ;
        RECT 90.040 152.790 90.215 152.825 ;
        RECT 89.285 152.255 89.615 152.655 ;
        RECT 90.040 152.425 90.570 152.790 ;
        RECT 90.760 152.425 91.035 152.935 ;
        RECT 91.205 152.425 91.395 153.785 ;
        RECT 91.565 153.800 91.735 154.465 ;
        RECT 91.905 154.045 92.075 154.805 ;
        RECT 92.310 154.045 92.825 154.455 ;
        RECT 91.565 153.610 92.315 153.800 ;
        RECT 92.485 153.235 92.825 154.045 ;
        RECT 92.995 153.640 93.285 154.805 ;
        RECT 93.455 153.730 93.725 154.635 ;
        RECT 93.895 154.045 94.225 154.805 ;
        RECT 94.405 153.875 94.575 154.635 ;
        RECT 91.595 153.065 92.825 153.235 ;
        RECT 91.575 152.255 92.085 152.790 ;
        RECT 92.305 152.460 92.550 153.065 ;
        RECT 92.995 152.255 93.285 152.980 ;
        RECT 93.455 152.930 93.625 153.730 ;
        RECT 93.910 153.705 94.575 153.875 ;
        RECT 93.910 153.560 94.080 153.705 ;
        RECT 93.795 153.230 94.080 153.560 ;
        RECT 93.910 152.975 94.080 153.230 ;
        RECT 94.315 153.155 94.645 153.525 ;
        RECT 93.455 152.425 93.715 152.930 ;
        RECT 93.910 152.805 94.575 152.975 ;
        RECT 93.895 152.255 94.225 152.635 ;
        RECT 94.405 152.425 94.575 152.805 ;
        RECT 95.755 152.425 96.505 154.635 ;
        RECT 97.595 154.045 98.110 154.455 ;
        RECT 98.345 154.045 98.515 154.805 ;
        RECT 98.685 154.465 100.715 154.635 ;
        RECT 97.595 153.235 97.935 154.045 ;
        RECT 98.685 153.800 98.855 154.465 ;
        RECT 99.250 154.125 100.375 154.295 ;
        RECT 98.105 153.610 98.855 153.800 ;
        RECT 99.025 153.785 100.035 153.955 ;
        RECT 97.595 153.065 98.825 153.235 ;
        RECT 97.870 152.460 98.115 153.065 ;
        RECT 98.335 152.255 98.845 152.790 ;
        RECT 99.025 152.425 99.215 153.785 ;
        RECT 99.385 153.105 99.660 153.585 ;
        RECT 99.385 152.935 99.665 153.105 ;
        RECT 99.865 152.985 100.035 153.785 ;
        RECT 100.205 152.995 100.375 154.125 ;
        RECT 100.545 153.495 100.715 154.465 ;
        RECT 100.885 153.665 101.055 154.805 ;
        RECT 101.225 153.665 101.560 154.635 ;
        RECT 101.735 153.715 103.405 154.805 ;
        RECT 103.580 154.135 103.835 154.635 ;
        RECT 104.005 154.305 104.335 154.805 ;
        RECT 103.580 153.965 104.330 154.135 ;
        RECT 100.545 153.165 100.740 153.495 ;
        RECT 100.965 153.165 101.220 153.495 ;
        RECT 100.965 152.995 101.135 153.165 ;
        RECT 101.390 152.995 101.560 153.665 ;
        RECT 99.385 152.425 99.660 152.935 ;
        RECT 100.205 152.825 101.135 152.995 ;
        RECT 100.205 152.790 100.380 152.825 ;
        RECT 99.850 152.425 100.380 152.790 ;
        RECT 100.805 152.255 101.135 152.655 ;
        RECT 101.305 152.425 101.560 152.995 ;
        RECT 101.735 153.025 102.485 153.545 ;
        RECT 102.655 153.195 103.405 153.715 ;
        RECT 103.580 153.145 103.930 153.795 ;
        RECT 101.735 152.255 103.405 153.025 ;
        RECT 104.100 152.975 104.330 153.965 ;
        RECT 103.580 152.805 104.330 152.975 ;
        RECT 103.580 152.515 103.835 152.805 ;
        RECT 104.005 152.255 104.335 152.635 ;
        RECT 104.505 152.515 104.675 154.635 ;
        RECT 104.845 153.835 105.170 154.620 ;
        RECT 105.340 154.345 105.590 154.805 ;
        RECT 105.760 154.305 106.010 154.635 ;
        RECT 106.225 154.305 106.905 154.635 ;
        RECT 105.760 154.175 105.930 154.305 ;
        RECT 105.535 154.005 105.930 154.175 ;
        RECT 104.905 152.785 105.365 153.835 ;
        RECT 105.535 152.645 105.705 154.005 ;
        RECT 106.100 153.745 106.565 154.135 ;
        RECT 105.875 152.935 106.225 153.555 ;
        RECT 106.395 153.155 106.565 153.745 ;
        RECT 106.735 153.525 106.905 154.305 ;
        RECT 107.075 154.205 107.245 154.545 ;
        RECT 107.480 154.375 107.810 154.805 ;
        RECT 107.980 154.205 108.150 154.545 ;
        RECT 108.445 154.345 108.815 154.805 ;
        RECT 107.075 154.035 108.150 154.205 ;
        RECT 108.985 154.175 109.155 154.635 ;
        RECT 109.390 154.295 110.260 154.635 ;
        RECT 110.430 154.345 110.680 154.805 ;
        RECT 108.595 154.005 109.155 154.175 ;
        RECT 108.595 153.865 108.765 154.005 ;
        RECT 107.265 153.695 108.765 153.865 ;
        RECT 109.460 153.835 109.920 154.125 ;
        RECT 106.735 153.355 108.425 153.525 ;
        RECT 106.395 152.935 106.750 153.155 ;
        RECT 106.920 152.645 107.090 153.355 ;
        RECT 107.295 152.935 108.085 153.185 ;
        RECT 108.255 153.175 108.425 153.355 ;
        RECT 108.595 153.005 108.765 153.695 ;
        RECT 105.035 152.255 105.365 152.615 ;
        RECT 105.535 152.475 106.030 152.645 ;
        RECT 106.235 152.475 107.090 152.645 ;
        RECT 107.965 152.255 108.295 152.715 ;
        RECT 108.505 152.615 108.765 153.005 ;
        RECT 108.955 153.825 109.920 153.835 ;
        RECT 110.090 153.915 110.260 154.295 ;
        RECT 110.850 154.255 111.020 154.545 ;
        RECT 111.200 154.425 111.530 154.805 ;
        RECT 110.850 154.085 111.650 154.255 ;
        RECT 108.955 153.665 109.630 153.825 ;
        RECT 110.090 153.745 111.310 153.915 ;
        RECT 108.955 152.875 109.165 153.665 ;
        RECT 110.090 153.655 110.260 153.745 ;
        RECT 109.335 152.875 109.685 153.495 ;
        RECT 109.855 153.485 110.260 153.655 ;
        RECT 109.855 152.705 110.025 153.485 ;
        RECT 110.195 153.035 110.415 153.315 ;
        RECT 110.595 153.205 111.135 153.575 ;
        RECT 111.480 153.495 111.650 154.085 ;
        RECT 111.870 153.665 112.175 154.805 ;
        RECT 112.345 153.615 112.595 154.495 ;
        RECT 112.765 153.665 113.015 154.805 ;
        RECT 113.325 153.875 113.495 154.635 ;
        RECT 113.675 154.045 114.005 154.805 ;
        RECT 113.325 153.705 113.990 153.875 ;
        RECT 114.175 153.730 114.445 154.635 ;
        RECT 111.480 153.465 112.220 153.495 ;
        RECT 110.195 152.865 110.725 153.035 ;
        RECT 108.505 152.445 108.855 152.615 ;
        RECT 109.075 152.425 110.025 152.705 ;
        RECT 110.195 152.255 110.385 152.695 ;
        RECT 110.555 152.635 110.725 152.865 ;
        RECT 110.895 152.805 111.135 153.205 ;
        RECT 111.305 153.165 112.220 153.465 ;
        RECT 111.305 152.990 111.630 153.165 ;
        RECT 111.305 152.635 111.625 152.990 ;
        RECT 112.390 152.965 112.595 153.615 ;
        RECT 113.820 153.560 113.990 153.705 ;
        RECT 113.255 153.155 113.585 153.525 ;
        RECT 113.820 153.230 114.105 153.560 ;
        RECT 110.555 152.465 111.625 152.635 ;
        RECT 111.870 152.255 112.175 152.715 ;
        RECT 112.345 152.435 112.595 152.965 ;
        RECT 112.765 152.255 113.015 153.010 ;
        RECT 113.820 152.975 113.990 153.230 ;
        RECT 113.325 152.805 113.990 152.975 ;
        RECT 114.275 152.930 114.445 153.730 ;
        RECT 114.615 154.045 115.130 154.455 ;
        RECT 115.365 154.045 115.535 154.805 ;
        RECT 115.705 154.465 117.735 154.635 ;
        RECT 114.615 153.235 114.955 154.045 ;
        RECT 115.705 153.800 115.875 154.465 ;
        RECT 116.270 154.125 117.395 154.295 ;
        RECT 115.125 153.610 115.875 153.800 ;
        RECT 116.045 153.785 117.055 153.955 ;
        RECT 114.615 153.065 115.845 153.235 ;
        RECT 113.325 152.425 113.495 152.805 ;
        RECT 113.675 152.255 114.005 152.635 ;
        RECT 114.185 152.425 114.445 152.930 ;
        RECT 114.890 152.460 115.135 153.065 ;
        RECT 115.355 152.255 115.865 152.790 ;
        RECT 116.045 152.425 116.235 153.785 ;
        RECT 116.405 152.765 116.680 153.585 ;
        RECT 116.885 152.985 117.055 153.785 ;
        RECT 117.225 152.995 117.395 154.125 ;
        RECT 117.565 153.495 117.735 154.465 ;
        RECT 117.905 153.665 118.075 154.805 ;
        RECT 118.245 153.665 118.580 154.635 ;
        RECT 117.565 153.165 117.760 153.495 ;
        RECT 117.985 153.165 118.240 153.495 ;
        RECT 117.985 152.995 118.155 153.165 ;
        RECT 118.410 152.995 118.580 153.665 ;
        RECT 118.755 153.640 119.045 154.805 ;
        RECT 119.220 153.665 119.475 154.805 ;
        RECT 119.670 154.255 120.865 154.585 ;
        RECT 119.725 153.495 119.895 154.055 ;
        RECT 120.120 153.835 120.540 154.085 ;
        RECT 121.045 154.005 121.325 154.805 ;
        RECT 120.120 153.665 121.365 153.835 ;
        RECT 121.535 153.665 121.805 154.635 ;
        RECT 121.980 154.135 122.235 154.635 ;
        RECT 122.405 154.305 122.735 154.805 ;
        RECT 121.980 153.965 122.730 154.135 ;
        RECT 121.195 153.495 121.365 153.665 ;
        RECT 119.220 153.245 119.555 153.495 ;
        RECT 119.725 153.165 120.465 153.495 ;
        RECT 121.195 153.165 121.425 153.495 ;
        RECT 119.725 153.075 119.975 153.165 ;
        RECT 117.225 152.825 118.155 152.995 ;
        RECT 117.225 152.790 117.400 152.825 ;
        RECT 116.405 152.595 116.685 152.765 ;
        RECT 116.405 152.425 116.680 152.595 ;
        RECT 116.870 152.425 117.400 152.790 ;
        RECT 117.825 152.255 118.155 152.655 ;
        RECT 118.325 152.425 118.580 152.995 ;
        RECT 118.755 152.255 119.045 152.980 ;
        RECT 119.240 152.905 119.975 153.075 ;
        RECT 121.195 152.995 121.365 153.165 ;
        RECT 119.240 152.435 119.550 152.905 ;
        RECT 120.625 152.825 121.365 152.995 ;
        RECT 121.635 152.930 121.805 153.665 ;
        RECT 121.980 153.145 122.330 153.795 ;
        RECT 122.500 152.975 122.730 153.965 ;
        RECT 119.720 152.255 120.455 152.735 ;
        RECT 120.625 152.475 120.795 152.825 ;
        RECT 120.965 152.255 121.345 152.655 ;
        RECT 121.535 152.585 121.805 152.930 ;
        RECT 121.980 152.805 122.730 152.975 ;
        RECT 121.980 152.515 122.235 152.805 ;
        RECT 122.405 152.255 122.735 152.635 ;
        RECT 122.905 152.515 123.075 154.635 ;
        RECT 123.245 153.835 123.570 154.620 ;
        RECT 123.740 154.345 123.990 154.805 ;
        RECT 124.160 154.305 124.410 154.635 ;
        RECT 124.625 154.305 125.305 154.635 ;
        RECT 124.160 154.175 124.330 154.305 ;
        RECT 123.935 154.005 124.330 154.175 ;
        RECT 123.305 152.785 123.765 153.835 ;
        RECT 123.935 152.645 124.105 154.005 ;
        RECT 124.500 153.745 124.965 154.135 ;
        RECT 124.275 152.935 124.625 153.555 ;
        RECT 124.795 153.155 124.965 153.745 ;
        RECT 125.135 153.525 125.305 154.305 ;
        RECT 125.475 154.205 125.645 154.545 ;
        RECT 125.880 154.375 126.210 154.805 ;
        RECT 126.380 154.205 126.550 154.545 ;
        RECT 126.845 154.345 127.215 154.805 ;
        RECT 125.475 154.035 126.550 154.205 ;
        RECT 127.385 154.175 127.555 154.635 ;
        RECT 127.790 154.295 128.660 154.635 ;
        RECT 128.830 154.345 129.080 154.805 ;
        RECT 126.995 154.005 127.555 154.175 ;
        RECT 126.995 153.865 127.165 154.005 ;
        RECT 125.665 153.695 127.165 153.865 ;
        RECT 127.860 153.835 128.320 154.125 ;
        RECT 125.135 153.355 126.825 153.525 ;
        RECT 124.795 152.935 125.150 153.155 ;
        RECT 125.320 152.645 125.490 153.355 ;
        RECT 125.695 152.935 126.485 153.185 ;
        RECT 126.655 153.175 126.825 153.355 ;
        RECT 126.995 153.005 127.165 153.695 ;
        RECT 123.435 152.255 123.765 152.615 ;
        RECT 123.935 152.475 124.430 152.645 ;
        RECT 124.635 152.475 125.490 152.645 ;
        RECT 126.365 152.255 126.695 152.715 ;
        RECT 126.905 152.615 127.165 153.005 ;
        RECT 127.355 153.825 128.320 153.835 ;
        RECT 128.490 153.915 128.660 154.295 ;
        RECT 129.250 154.255 129.420 154.545 ;
        RECT 129.600 154.425 129.930 154.805 ;
        RECT 129.250 154.085 130.050 154.255 ;
        RECT 127.355 153.665 128.030 153.825 ;
        RECT 128.490 153.745 129.710 153.915 ;
        RECT 127.355 152.875 127.565 153.665 ;
        RECT 128.490 153.655 128.660 153.745 ;
        RECT 127.735 152.875 128.085 153.495 ;
        RECT 128.255 153.485 128.660 153.655 ;
        RECT 128.255 152.705 128.425 153.485 ;
        RECT 128.595 153.035 128.815 153.315 ;
        RECT 128.995 153.205 129.535 153.575 ;
        RECT 129.880 153.495 130.050 154.085 ;
        RECT 130.270 153.665 130.575 154.805 ;
        RECT 130.745 153.615 131.000 154.495 ;
        RECT 129.880 153.465 130.620 153.495 ;
        RECT 128.595 152.865 129.125 153.035 ;
        RECT 126.905 152.445 127.255 152.615 ;
        RECT 127.475 152.425 128.425 152.705 ;
        RECT 128.595 152.255 128.785 152.695 ;
        RECT 128.955 152.635 129.125 152.865 ;
        RECT 129.295 152.805 129.535 153.205 ;
        RECT 129.705 153.165 130.620 153.465 ;
        RECT 129.705 152.990 130.030 153.165 ;
        RECT 129.705 152.635 130.025 152.990 ;
        RECT 130.790 152.965 131.000 153.615 ;
        RECT 128.955 152.465 130.025 152.635 ;
        RECT 130.270 152.255 130.575 152.715 ;
        RECT 130.745 152.435 131.000 152.965 ;
        RECT 132.095 152.425 132.845 154.635 ;
        RECT 133.940 154.175 134.275 154.635 ;
        RECT 134.445 154.345 134.665 154.805 ;
        RECT 135.195 154.425 136.505 154.595 ;
        RECT 136.335 154.175 136.505 154.425 ;
        RECT 136.675 154.345 136.965 154.805 ;
        RECT 133.940 154.005 136.165 154.175 ;
        RECT 136.335 154.005 136.995 154.175 ;
        RECT 133.940 152.425 134.270 154.005 ;
        RECT 135.995 153.835 136.165 154.005 ;
        RECT 134.440 152.925 134.630 153.795 ;
        RECT 134.900 153.485 135.715 153.795 ;
        RECT 135.995 153.665 136.655 153.835 ;
        RECT 135.545 153.450 135.715 153.485 ;
        RECT 134.900 152.905 135.365 153.195 ;
        RECT 135.545 152.935 136.175 153.450 ;
        RECT 136.485 153.165 136.655 153.665 ;
        RECT 136.825 153.495 136.995 154.005 ;
        RECT 137.165 153.765 137.475 154.635 ;
        RECT 136.825 153.165 137.135 153.495 ;
        RECT 136.825 152.975 136.995 153.165 ;
        RECT 134.440 152.255 134.640 152.755 ;
        RECT 134.900 152.590 135.090 152.905 ;
        RECT 136.385 152.805 136.995 152.975 ;
        RECT 137.305 152.920 137.475 153.765 ;
        RECT 137.645 153.665 137.900 154.805 ;
        RECT 138.165 153.875 138.335 154.635 ;
        RECT 138.515 154.045 138.845 154.805 ;
        RECT 138.165 153.705 138.830 153.875 ;
        RECT 139.015 153.730 139.285 154.635 ;
        RECT 138.660 153.560 138.830 153.705 ;
        RECT 138.095 153.155 138.425 153.525 ;
        RECT 138.660 153.230 138.945 153.560 ;
        RECT 136.385 152.635 136.555 152.805 ;
        RECT 135.260 152.465 136.555 152.635 ;
        RECT 136.725 152.255 137.055 152.635 ;
        RECT 137.225 152.425 137.475 152.920 ;
        RECT 137.645 152.255 137.900 153.055 ;
        RECT 138.660 152.975 138.830 153.230 ;
        RECT 138.165 152.805 138.830 152.975 ;
        RECT 139.115 152.930 139.285 153.730 ;
        RECT 138.165 152.425 138.335 152.805 ;
        RECT 138.515 152.255 138.845 152.635 ;
        RECT 139.025 152.425 139.285 152.930 ;
        RECT 139.455 153.730 139.725 154.635 ;
        RECT 139.895 154.045 140.225 154.805 ;
        RECT 140.405 153.875 140.575 154.635 ;
        RECT 139.455 152.930 139.625 153.730 ;
        RECT 139.910 153.705 140.575 153.875 ;
        RECT 140.835 153.715 144.345 154.805 ;
        RECT 139.910 153.560 140.080 153.705 ;
        RECT 139.795 153.230 140.080 153.560 ;
        RECT 139.910 152.975 140.080 153.230 ;
        RECT 140.315 153.155 140.645 153.525 ;
        RECT 140.835 153.025 142.485 153.545 ;
        RECT 142.655 153.195 144.345 153.715 ;
        RECT 144.515 153.640 144.805 154.805 ;
        RECT 144.975 154.370 150.320 154.805 ;
        RECT 150.495 154.370 155.840 154.805 ;
        RECT 139.455 152.425 139.715 152.930 ;
        RECT 139.910 152.805 140.575 152.975 ;
        RECT 139.895 152.255 140.225 152.635 ;
        RECT 140.405 152.425 140.575 152.805 ;
        RECT 140.835 152.255 144.345 153.025 ;
        RECT 144.515 152.255 144.805 152.980 ;
        RECT 146.560 152.800 146.900 153.630 ;
        RECT 148.380 153.120 148.730 154.370 ;
        RECT 152.080 152.800 152.420 153.630 ;
        RECT 153.900 153.120 154.250 154.370 ;
        RECT 156.935 153.715 158.145 154.805 ;
        RECT 156.935 153.175 157.455 153.715 ;
        RECT 157.625 153.005 158.145 153.545 ;
        RECT 144.975 152.255 150.320 152.800 ;
        RECT 150.495 152.255 155.840 152.800 ;
        RECT 156.935 152.255 158.145 153.005 ;
        RECT 2.750 152.085 158.230 152.255 ;
        RECT 2.835 151.335 4.045 152.085 ;
        RECT 5.225 151.535 5.395 151.915 ;
        RECT 5.575 151.705 5.905 152.085 ;
        RECT 5.225 151.365 5.890 151.535 ;
        RECT 6.085 151.410 6.345 151.915 ;
        RECT 2.835 150.795 3.355 151.335 ;
        RECT 3.525 150.625 4.045 151.165 ;
        RECT 5.155 150.815 5.485 151.185 ;
        RECT 5.720 151.110 5.890 151.365 ;
        RECT 5.720 150.780 6.005 151.110 ;
        RECT 5.720 150.635 5.890 150.780 ;
        RECT 2.835 149.535 4.045 150.625 ;
        RECT 5.225 150.465 5.890 150.635 ;
        RECT 6.175 150.610 6.345 151.410 ;
        RECT 6.565 151.545 6.790 151.905 ;
        RECT 6.970 151.715 7.300 152.085 ;
        RECT 7.480 151.545 7.735 151.905 ;
        RECT 8.300 151.715 9.045 152.085 ;
        RECT 6.565 151.355 9.050 151.545 ;
        RECT 6.525 150.845 6.795 151.175 ;
        RECT 6.975 150.845 7.410 151.175 ;
        RECT 7.590 150.845 8.165 151.175 ;
        RECT 8.345 150.845 8.625 151.175 ;
        RECT 8.825 150.665 9.050 151.355 ;
        RECT 5.225 149.705 5.395 150.465 ;
        RECT 5.575 149.535 5.905 150.295 ;
        RECT 6.075 149.705 6.345 150.610 ;
        RECT 6.555 150.485 9.050 150.665 ;
        RECT 9.225 150.485 9.560 151.905 ;
        RECT 9.740 151.535 9.995 151.825 ;
        RECT 10.165 151.705 10.495 152.085 ;
        RECT 9.740 151.365 10.490 151.535 ;
        RECT 9.740 150.545 10.090 151.195 ;
        RECT 6.555 149.715 6.845 150.485 ;
        RECT 7.415 150.075 8.605 150.305 ;
        RECT 7.415 149.715 7.675 150.075 ;
        RECT 7.845 149.535 8.175 149.905 ;
        RECT 8.345 149.715 8.605 150.075 ;
        RECT 8.795 149.535 9.125 150.255 ;
        RECT 9.295 149.715 9.560 150.485 ;
        RECT 10.260 150.375 10.490 151.365 ;
        RECT 9.740 150.205 10.490 150.375 ;
        RECT 9.740 149.705 9.995 150.205 ;
        RECT 10.165 149.535 10.495 150.035 ;
        RECT 10.665 149.705 10.835 151.825 ;
        RECT 11.195 151.725 11.525 152.085 ;
        RECT 11.695 151.695 12.190 151.865 ;
        RECT 12.395 151.695 13.250 151.865 ;
        RECT 11.065 150.505 11.525 151.555 ;
        RECT 11.005 149.720 11.330 150.505 ;
        RECT 11.695 150.335 11.865 151.695 ;
        RECT 12.035 150.785 12.385 151.405 ;
        RECT 12.555 151.185 12.910 151.405 ;
        RECT 12.555 150.595 12.725 151.185 ;
        RECT 13.080 150.985 13.250 151.695 ;
        RECT 14.125 151.625 14.455 152.085 ;
        RECT 14.665 151.725 15.015 151.895 ;
        RECT 13.455 151.155 14.245 151.405 ;
        RECT 14.665 151.335 14.925 151.725 ;
        RECT 15.235 151.635 16.185 151.915 ;
        RECT 16.355 151.645 16.545 152.085 ;
        RECT 16.715 151.705 17.785 151.875 ;
        RECT 14.415 150.985 14.585 151.165 ;
        RECT 11.695 150.165 12.090 150.335 ;
        RECT 12.260 150.205 12.725 150.595 ;
        RECT 12.895 150.815 14.585 150.985 ;
        RECT 11.920 150.035 12.090 150.165 ;
        RECT 12.895 150.035 13.065 150.815 ;
        RECT 14.755 150.645 14.925 151.335 ;
        RECT 13.425 150.475 14.925 150.645 ;
        RECT 15.115 150.675 15.325 151.465 ;
        RECT 15.495 150.845 15.845 151.465 ;
        RECT 16.015 150.855 16.185 151.635 ;
        RECT 16.715 151.475 16.885 151.705 ;
        RECT 16.355 151.305 16.885 151.475 ;
        RECT 16.355 151.025 16.575 151.305 ;
        RECT 17.055 151.135 17.295 151.535 ;
        RECT 16.015 150.685 16.420 150.855 ;
        RECT 16.755 150.765 17.295 151.135 ;
        RECT 17.465 151.350 17.785 151.705 ;
        RECT 18.030 151.625 18.335 152.085 ;
        RECT 18.505 151.375 18.760 151.905 ;
        RECT 17.465 151.175 17.790 151.350 ;
        RECT 17.465 150.875 18.380 151.175 ;
        RECT 17.640 150.845 18.380 150.875 ;
        RECT 15.115 150.515 15.790 150.675 ;
        RECT 16.250 150.595 16.420 150.685 ;
        RECT 15.115 150.505 16.080 150.515 ;
        RECT 14.755 150.335 14.925 150.475 ;
        RECT 11.500 149.535 11.750 149.995 ;
        RECT 11.920 149.705 12.170 150.035 ;
        RECT 12.385 149.705 13.065 150.035 ;
        RECT 13.235 150.135 14.310 150.305 ;
        RECT 14.755 150.165 15.315 150.335 ;
        RECT 15.620 150.215 16.080 150.505 ;
        RECT 16.250 150.425 17.470 150.595 ;
        RECT 13.235 149.795 13.405 150.135 ;
        RECT 13.640 149.535 13.970 149.965 ;
        RECT 14.140 149.795 14.310 150.135 ;
        RECT 14.605 149.535 14.975 149.995 ;
        RECT 15.145 149.705 15.315 150.165 ;
        RECT 16.250 150.045 16.420 150.425 ;
        RECT 17.640 150.255 17.810 150.845 ;
        RECT 18.550 150.725 18.760 151.375 ;
        RECT 15.550 149.705 16.420 150.045 ;
        RECT 17.010 150.085 17.810 150.255 ;
        RECT 16.590 149.535 16.840 149.995 ;
        RECT 17.010 149.795 17.180 150.085 ;
        RECT 17.360 149.535 17.690 149.915 ;
        RECT 18.030 149.535 18.335 150.675 ;
        RECT 18.505 149.845 18.760 150.725 ;
        RECT 18.935 151.345 19.320 151.915 ;
        RECT 19.490 151.625 19.815 152.085 ;
        RECT 20.335 151.455 20.615 151.915 ;
        RECT 18.935 150.675 19.215 151.345 ;
        RECT 19.490 151.285 20.615 151.455 ;
        RECT 19.490 151.175 19.940 151.285 ;
        RECT 19.385 150.845 19.940 151.175 ;
        RECT 20.805 151.115 21.205 151.915 ;
        RECT 21.605 151.625 21.875 152.085 ;
        RECT 22.045 151.455 22.330 151.915 ;
        RECT 18.935 149.705 19.320 150.675 ;
        RECT 19.490 150.385 19.940 150.845 ;
        RECT 20.110 150.555 21.205 151.115 ;
        RECT 19.490 150.165 20.615 150.385 ;
        RECT 19.490 149.535 19.815 149.995 ;
        RECT 20.335 149.705 20.615 150.165 ;
        RECT 20.805 149.705 21.205 150.555 ;
        RECT 21.375 151.285 22.330 151.455 ;
        RECT 21.375 150.385 21.585 151.285 ;
        RECT 23.595 151.265 23.805 152.085 ;
        RECT 23.975 151.285 24.305 151.915 ;
        RECT 21.755 150.555 22.445 151.115 ;
        RECT 23.975 150.685 24.225 151.285 ;
        RECT 24.475 151.265 24.705 152.085 ;
        RECT 25.015 151.285 25.185 152.085 ;
        RECT 24.395 150.845 24.725 151.095 ;
        RECT 21.375 150.165 22.330 150.385 ;
        RECT 21.605 149.535 21.875 149.995 ;
        RECT 22.045 149.705 22.330 150.165 ;
        RECT 23.595 149.535 23.805 150.675 ;
        RECT 23.975 149.705 24.305 150.685 ;
        RECT 24.475 149.535 24.705 150.675 ;
        RECT 24.945 149.535 25.195 150.725 ;
        RECT 25.420 149.705 25.635 151.805 ;
        RECT 25.855 151.625 26.035 152.085 ;
        RECT 26.295 151.695 27.560 151.875 ;
        RECT 26.680 151.455 27.045 151.525 ;
        RECT 25.805 151.275 27.045 151.455 ;
        RECT 27.220 151.475 27.560 151.695 ;
        RECT 27.745 151.645 27.915 152.085 ;
        RECT 28.085 151.475 28.420 151.890 ;
        RECT 27.220 151.345 28.420 151.475 ;
        RECT 28.595 151.360 28.885 152.085 ;
        RECT 27.390 151.305 28.420 151.345 ;
        RECT 29.155 151.285 29.325 152.085 ;
        RECT 25.805 150.675 26.085 151.275 ;
        RECT 26.265 150.845 26.620 151.095 ;
        RECT 26.790 150.845 27.255 151.095 ;
        RECT 27.425 150.845 27.755 151.095 ;
        RECT 27.925 150.895 28.420 151.095 ;
        RECT 27.575 150.725 27.755 150.845 ;
        RECT 25.805 150.465 27.405 150.675 ;
        RECT 27.575 150.555 27.930 150.725 ;
        RECT 28.100 150.555 28.420 150.895 ;
        RECT 25.825 149.535 26.625 150.295 ;
        RECT 27.020 149.705 27.405 150.465 ;
        RECT 27.730 149.765 27.930 150.555 ;
        RECT 28.100 149.535 28.420 150.375 ;
        RECT 28.595 149.535 28.885 150.700 ;
        RECT 29.085 149.535 29.335 150.725 ;
        RECT 29.560 149.705 29.775 151.805 ;
        RECT 29.995 151.625 30.175 152.085 ;
        RECT 30.435 151.695 31.700 151.875 ;
        RECT 30.820 151.455 31.185 151.525 ;
        RECT 29.945 151.275 31.185 151.455 ;
        RECT 31.360 151.475 31.700 151.695 ;
        RECT 31.885 151.645 32.055 152.085 ;
        RECT 32.225 151.475 32.560 151.890 ;
        RECT 31.360 151.345 32.560 151.475 ;
        RECT 31.530 151.305 32.560 151.345 ;
        RECT 29.945 150.675 30.225 151.275 ;
        RECT 30.405 150.845 30.760 151.095 ;
        RECT 30.930 150.845 31.395 151.095 ;
        RECT 31.565 150.845 31.895 151.095 ;
        RECT 32.065 150.895 32.560 151.095 ;
        RECT 31.715 150.725 31.895 150.845 ;
        RECT 29.945 150.465 31.545 150.675 ;
        RECT 31.715 150.555 32.070 150.725 ;
        RECT 32.240 150.555 32.560 150.895 ;
        RECT 29.965 149.535 30.765 150.295 ;
        RECT 31.160 149.705 31.545 150.465 ;
        RECT 31.870 149.765 32.070 150.555 ;
        RECT 32.740 150.485 33.075 151.905 ;
        RECT 33.255 151.715 34.000 152.085 ;
        RECT 34.565 151.545 34.820 151.905 ;
        RECT 35.000 151.715 35.330 152.085 ;
        RECT 35.510 151.545 35.735 151.905 ;
        RECT 33.250 151.355 35.735 151.545 ;
        RECT 33.250 150.665 33.475 151.355 ;
        RECT 36.875 151.345 37.260 151.915 ;
        RECT 37.430 151.625 37.755 152.085 ;
        RECT 38.275 151.455 38.555 151.915 ;
        RECT 33.675 150.845 33.955 151.175 ;
        RECT 34.135 150.845 34.710 151.175 ;
        RECT 34.890 150.845 35.325 151.175 ;
        RECT 35.505 150.845 35.775 151.175 ;
        RECT 36.875 150.675 37.155 151.345 ;
        RECT 37.430 151.285 38.555 151.455 ;
        RECT 37.430 151.175 37.880 151.285 ;
        RECT 37.325 150.845 37.880 151.175 ;
        RECT 38.745 151.115 39.145 151.915 ;
        RECT 39.545 151.625 39.815 152.085 ;
        RECT 39.985 151.455 40.270 151.915 ;
        RECT 33.250 150.485 35.745 150.665 ;
        RECT 32.240 149.535 32.560 150.375 ;
        RECT 32.740 149.715 33.005 150.485 ;
        RECT 33.175 149.535 33.505 150.255 ;
        RECT 33.695 150.075 34.885 150.305 ;
        RECT 33.695 149.715 33.955 150.075 ;
        RECT 34.125 149.535 34.455 149.905 ;
        RECT 34.625 149.715 34.885 150.075 ;
        RECT 35.455 149.715 35.745 150.485 ;
        RECT 36.875 149.705 37.260 150.675 ;
        RECT 37.430 150.385 37.880 150.845 ;
        RECT 38.050 150.555 39.145 151.115 ;
        RECT 37.430 150.165 38.555 150.385 ;
        RECT 37.430 149.535 37.755 149.995 ;
        RECT 38.275 149.705 38.555 150.165 ;
        RECT 38.745 149.705 39.145 150.555 ;
        RECT 39.315 151.285 40.270 151.455 ;
        RECT 41.015 151.585 41.275 151.915 ;
        RECT 41.445 151.725 41.775 152.085 ;
        RECT 42.030 151.705 43.330 151.915 ;
        RECT 39.315 150.385 39.525 151.285 ;
        RECT 39.695 150.555 40.385 151.115 ;
        RECT 41.015 150.385 41.185 151.585 ;
        RECT 42.030 151.555 42.200 151.705 ;
        RECT 41.445 151.430 42.200 151.555 ;
        RECT 41.355 151.385 42.200 151.430 ;
        RECT 41.355 151.265 41.625 151.385 ;
        RECT 41.355 150.690 41.525 151.265 ;
        RECT 41.755 150.825 42.165 151.130 ;
        RECT 42.455 151.095 42.665 151.495 ;
        RECT 42.335 150.885 42.665 151.095 ;
        RECT 42.910 151.095 43.130 151.495 ;
        RECT 43.605 151.320 44.060 152.085 ;
        RECT 44.335 151.285 44.505 152.085 ;
        RECT 42.910 150.885 43.385 151.095 ;
        RECT 43.575 150.895 44.065 151.095 ;
        RECT 41.355 150.655 41.555 150.690 ;
        RECT 42.885 150.655 44.060 150.715 ;
        RECT 41.355 150.545 44.060 150.655 ;
        RECT 41.415 150.485 43.215 150.545 ;
        RECT 42.885 150.455 43.215 150.485 ;
        RECT 39.315 150.165 40.270 150.385 ;
        RECT 39.545 149.535 39.815 149.995 ;
        RECT 39.985 149.705 40.270 150.165 ;
        RECT 41.015 149.705 41.275 150.385 ;
        RECT 41.445 149.535 41.695 150.315 ;
        RECT 41.945 150.285 42.780 150.295 ;
        RECT 43.370 150.285 43.555 150.375 ;
        RECT 41.945 150.085 43.555 150.285 ;
        RECT 41.945 149.705 42.195 150.085 ;
        RECT 43.325 150.045 43.555 150.085 ;
        RECT 43.805 149.925 44.060 150.545 ;
        RECT 42.365 149.535 42.720 149.915 ;
        RECT 43.725 149.705 44.060 149.925 ;
        RECT 44.265 149.535 44.515 150.725 ;
        RECT 44.740 149.705 44.955 151.805 ;
        RECT 45.175 151.625 45.355 152.085 ;
        RECT 45.615 151.695 46.880 151.875 ;
        RECT 46.000 151.455 46.365 151.525 ;
        RECT 45.125 151.275 46.365 151.455 ;
        RECT 46.540 151.475 46.880 151.695 ;
        RECT 47.065 151.645 47.235 152.085 ;
        RECT 47.405 151.475 47.740 151.890 ;
        RECT 46.540 151.345 47.740 151.475 ;
        RECT 46.710 151.305 47.740 151.345 ;
        RECT 48.380 151.320 48.835 152.085 ;
        RECT 49.110 151.705 50.410 151.915 ;
        RECT 50.665 151.725 50.995 152.085 ;
        RECT 50.240 151.555 50.410 151.705 ;
        RECT 51.165 151.585 51.425 151.915 ;
        RECT 45.125 150.675 45.405 151.275 ;
        RECT 49.310 151.095 49.530 151.495 ;
        RECT 45.585 150.845 45.940 151.095 ;
        RECT 46.110 150.845 46.575 151.095 ;
        RECT 46.745 150.845 47.075 151.095 ;
        RECT 47.245 150.895 47.740 151.095 ;
        RECT 48.375 150.895 48.865 151.095 ;
        RECT 46.895 150.725 47.075 150.845 ;
        RECT 45.125 150.465 46.725 150.675 ;
        RECT 46.895 150.555 47.250 150.725 ;
        RECT 47.420 150.555 47.740 150.895 ;
        RECT 49.055 150.885 49.530 151.095 ;
        RECT 49.775 151.095 49.985 151.495 ;
        RECT 50.240 151.430 50.995 151.555 ;
        RECT 50.240 151.385 51.085 151.430 ;
        RECT 50.815 151.265 51.085 151.385 ;
        RECT 49.775 150.885 50.105 151.095 ;
        RECT 50.275 150.825 50.685 151.130 ;
        RECT 48.380 150.655 49.555 150.715 ;
        RECT 50.915 150.690 51.085 151.265 ;
        RECT 50.885 150.655 51.085 150.690 ;
        RECT 45.145 149.535 45.945 150.295 ;
        RECT 46.340 149.705 46.725 150.465 ;
        RECT 47.050 149.765 47.250 150.555 ;
        RECT 48.380 150.545 51.085 150.655 ;
        RECT 47.420 149.535 47.740 150.375 ;
        RECT 48.380 149.925 48.635 150.545 ;
        RECT 49.225 150.485 51.025 150.545 ;
        RECT 49.225 150.455 49.555 150.485 ;
        RECT 51.255 150.385 51.425 151.585 ;
        RECT 48.885 150.285 49.070 150.375 ;
        RECT 49.660 150.285 50.495 150.295 ;
        RECT 48.885 150.085 50.495 150.285 ;
        RECT 48.885 150.045 49.115 150.085 ;
        RECT 48.380 149.705 48.715 149.925 ;
        RECT 49.720 149.535 50.075 149.915 ;
        RECT 50.245 149.705 50.495 150.085 ;
        RECT 50.745 149.535 50.995 150.315 ;
        RECT 51.165 149.705 51.425 150.385 ;
        RECT 51.605 149.715 51.865 151.905 ;
        RECT 52.125 151.715 52.795 152.085 ;
        RECT 52.975 151.535 53.285 151.905 ;
        RECT 52.055 151.335 53.285 151.535 ;
        RECT 52.055 150.665 52.345 151.335 ;
        RECT 53.465 151.155 53.695 151.795 ;
        RECT 53.875 151.355 54.165 152.085 ;
        RECT 54.355 151.360 54.645 152.085 ;
        RECT 54.905 151.535 55.075 151.915 ;
        RECT 55.255 151.705 55.585 152.085 ;
        RECT 54.905 151.365 55.570 151.535 ;
        RECT 55.765 151.410 56.025 151.915 ;
        RECT 52.525 150.845 52.990 151.155 ;
        RECT 53.170 150.845 53.695 151.155 ;
        RECT 53.875 150.845 54.175 151.175 ;
        RECT 54.835 150.815 55.165 151.185 ;
        RECT 55.400 151.110 55.570 151.365 ;
        RECT 55.400 150.780 55.685 151.110 ;
        RECT 52.055 150.445 52.825 150.665 ;
        RECT 52.035 149.535 52.375 150.265 ;
        RECT 52.555 149.715 52.825 150.445 ;
        RECT 53.005 150.425 54.165 150.665 ;
        RECT 53.005 149.715 53.235 150.425 ;
        RECT 53.405 149.535 53.735 150.245 ;
        RECT 53.905 149.715 54.165 150.425 ;
        RECT 54.355 149.535 54.645 150.700 ;
        RECT 55.400 150.635 55.570 150.780 ;
        RECT 54.905 150.465 55.570 150.635 ;
        RECT 55.855 150.610 56.025 151.410 ;
        RECT 54.905 149.705 55.075 150.465 ;
        RECT 55.255 149.535 55.585 150.295 ;
        RECT 55.755 149.705 56.025 150.610 ;
        RECT 56.200 151.345 56.455 151.915 ;
        RECT 56.625 151.685 56.955 152.085 ;
        RECT 57.380 151.550 57.910 151.915 ;
        RECT 57.380 151.515 57.555 151.550 ;
        RECT 56.625 151.345 57.555 151.515 ;
        RECT 56.200 150.675 56.370 151.345 ;
        RECT 56.625 151.175 56.795 151.345 ;
        RECT 56.540 150.845 56.795 151.175 ;
        RECT 57.020 150.845 57.215 151.175 ;
        RECT 56.200 149.705 56.535 150.675 ;
        RECT 56.705 149.535 56.875 150.675 ;
        RECT 57.045 149.875 57.215 150.845 ;
        RECT 57.385 150.215 57.555 151.345 ;
        RECT 57.725 150.555 57.895 151.355 ;
        RECT 58.100 151.065 58.375 151.915 ;
        RECT 58.095 150.895 58.375 151.065 ;
        RECT 58.100 150.755 58.375 150.895 ;
        RECT 58.545 150.555 58.735 151.915 ;
        RECT 58.915 151.550 59.425 152.085 ;
        RECT 59.645 151.275 59.890 151.880 ;
        RECT 60.340 151.345 60.595 151.915 ;
        RECT 60.765 151.685 61.095 152.085 ;
        RECT 61.520 151.550 62.050 151.915 ;
        RECT 62.240 151.745 62.515 151.915 ;
        RECT 62.235 151.575 62.515 151.745 ;
        RECT 61.520 151.515 61.695 151.550 ;
        RECT 60.765 151.345 61.695 151.515 ;
        RECT 58.935 151.105 60.165 151.275 ;
        RECT 57.725 150.385 58.735 150.555 ;
        RECT 58.905 150.540 59.655 150.730 ;
        RECT 57.385 150.045 58.510 150.215 ;
        RECT 58.905 149.875 59.075 150.540 ;
        RECT 59.825 150.295 60.165 151.105 ;
        RECT 57.045 149.705 59.075 149.875 ;
        RECT 59.245 149.535 59.415 150.295 ;
        RECT 59.650 149.885 60.165 150.295 ;
        RECT 60.340 150.675 60.510 151.345 ;
        RECT 60.765 151.175 60.935 151.345 ;
        RECT 60.680 150.845 60.935 151.175 ;
        RECT 61.160 150.845 61.355 151.175 ;
        RECT 60.340 149.705 60.675 150.675 ;
        RECT 60.845 149.535 61.015 150.675 ;
        RECT 61.185 149.875 61.355 150.845 ;
        RECT 61.525 150.215 61.695 151.345 ;
        RECT 61.865 150.555 62.035 151.355 ;
        RECT 62.240 150.755 62.515 151.575 ;
        RECT 62.685 150.555 62.875 151.915 ;
        RECT 63.055 151.550 63.565 152.085 ;
        RECT 63.785 151.275 64.030 151.880 ;
        RECT 64.475 151.345 64.860 151.915 ;
        RECT 65.030 151.625 65.355 152.085 ;
        RECT 65.875 151.455 66.155 151.915 ;
        RECT 63.075 151.105 64.305 151.275 ;
        RECT 61.865 150.385 62.875 150.555 ;
        RECT 63.045 150.540 63.795 150.730 ;
        RECT 61.525 150.045 62.650 150.215 ;
        RECT 63.045 149.875 63.215 150.540 ;
        RECT 63.965 150.295 64.305 151.105 ;
        RECT 61.185 149.705 63.215 149.875 ;
        RECT 63.385 149.535 63.555 150.295 ;
        RECT 63.790 149.885 64.305 150.295 ;
        RECT 64.475 150.675 64.755 151.345 ;
        RECT 65.030 151.285 66.155 151.455 ;
        RECT 65.030 151.175 65.480 151.285 ;
        RECT 64.925 150.845 65.480 151.175 ;
        RECT 66.345 151.115 66.745 151.915 ;
        RECT 67.145 151.625 67.415 152.085 ;
        RECT 67.585 151.455 67.870 151.915 ;
        RECT 64.475 149.705 64.860 150.675 ;
        RECT 65.030 150.385 65.480 150.845 ;
        RECT 65.650 150.555 66.745 151.115 ;
        RECT 65.030 150.165 66.155 150.385 ;
        RECT 65.030 149.535 65.355 149.995 ;
        RECT 65.875 149.705 66.155 150.165 ;
        RECT 66.345 149.705 66.745 150.555 ;
        RECT 66.915 151.285 67.870 151.455 ;
        RECT 68.155 151.285 68.465 152.085 ;
        RECT 68.670 151.285 69.365 151.915 ;
        RECT 69.625 151.605 69.925 152.085 ;
        RECT 70.095 151.435 70.355 151.890 ;
        RECT 70.525 151.605 70.785 152.085 ;
        RECT 70.965 151.435 71.225 151.890 ;
        RECT 71.395 151.605 71.645 152.085 ;
        RECT 71.825 151.435 72.085 151.890 ;
        RECT 72.255 151.605 72.505 152.085 ;
        RECT 72.685 151.435 72.945 151.890 ;
        RECT 73.115 151.605 73.360 152.085 ;
        RECT 73.530 151.435 73.805 151.890 ;
        RECT 73.975 151.605 74.220 152.085 ;
        RECT 74.390 151.435 74.650 151.890 ;
        RECT 74.820 151.605 75.080 152.085 ;
        RECT 75.250 151.435 75.510 151.890 ;
        RECT 75.680 151.605 75.940 152.085 ;
        RECT 76.110 151.435 76.370 151.890 ;
        RECT 76.540 151.525 76.800 152.085 ;
        RECT 66.915 150.385 67.125 151.285 ;
        RECT 67.295 150.555 67.985 151.115 ;
        RECT 68.165 150.845 68.500 151.115 ;
        RECT 68.670 150.685 68.840 151.285 ;
        RECT 69.625 151.265 76.370 151.435 ;
        RECT 69.010 150.845 69.345 151.095 ;
        RECT 66.915 150.165 67.870 150.385 ;
        RECT 67.145 149.535 67.415 149.995 ;
        RECT 67.585 149.705 67.870 150.165 ;
        RECT 68.155 149.535 68.435 150.675 ;
        RECT 68.605 149.705 68.935 150.685 ;
        RECT 69.625 150.675 70.790 151.265 ;
        RECT 76.970 151.095 77.220 151.905 ;
        RECT 77.400 151.560 77.660 152.085 ;
        RECT 77.830 151.095 78.080 151.905 ;
        RECT 78.260 151.575 78.565 152.085 ;
        RECT 70.960 150.845 78.080 151.095 ;
        RECT 78.250 150.845 78.565 151.405 ;
        RECT 78.735 151.335 79.945 152.085 ;
        RECT 80.115 151.360 80.405 152.085 ;
        RECT 80.580 151.535 80.835 151.825 ;
        RECT 81.005 151.705 81.335 152.085 ;
        RECT 80.580 151.365 81.330 151.535 ;
        RECT 69.105 149.535 69.365 150.675 ;
        RECT 69.625 150.450 76.370 150.675 ;
        RECT 69.625 149.535 69.895 150.280 ;
        RECT 70.065 149.710 70.355 150.450 ;
        RECT 70.965 150.435 76.370 150.450 ;
        RECT 70.525 149.540 70.780 150.265 ;
        RECT 70.965 149.710 71.225 150.435 ;
        RECT 71.395 149.540 71.640 150.265 ;
        RECT 71.825 149.710 72.085 150.435 ;
        RECT 72.255 149.540 72.500 150.265 ;
        RECT 72.685 149.710 72.945 150.435 ;
        RECT 73.115 149.540 73.360 150.265 ;
        RECT 73.530 149.710 73.790 150.435 ;
        RECT 73.960 149.540 74.220 150.265 ;
        RECT 74.390 149.710 74.650 150.435 ;
        RECT 74.820 149.540 75.080 150.265 ;
        RECT 75.250 149.710 75.510 150.435 ;
        RECT 75.680 149.540 75.940 150.265 ;
        RECT 76.110 149.710 76.370 150.435 ;
        RECT 76.540 149.540 76.800 150.335 ;
        RECT 76.970 149.710 77.220 150.845 ;
        RECT 70.525 149.535 76.800 149.540 ;
        RECT 77.400 149.535 77.660 150.345 ;
        RECT 77.835 149.705 78.080 150.845 ;
        RECT 78.735 150.795 79.255 151.335 ;
        RECT 79.425 150.625 79.945 151.165 ;
        RECT 78.260 149.535 78.555 150.345 ;
        RECT 78.735 149.535 79.945 150.625 ;
        RECT 80.115 149.535 80.405 150.700 ;
        RECT 80.580 150.545 80.930 151.195 ;
        RECT 81.100 150.375 81.330 151.365 ;
        RECT 80.580 150.205 81.330 150.375 ;
        RECT 80.580 149.705 80.835 150.205 ;
        RECT 81.005 149.535 81.335 150.035 ;
        RECT 81.505 149.705 81.675 151.825 ;
        RECT 82.035 151.725 82.365 152.085 ;
        RECT 82.535 151.695 83.030 151.865 ;
        RECT 83.235 151.695 84.090 151.865 ;
        RECT 81.905 150.505 82.365 151.555 ;
        RECT 81.845 149.720 82.170 150.505 ;
        RECT 82.535 150.335 82.705 151.695 ;
        RECT 82.875 150.785 83.225 151.405 ;
        RECT 83.395 151.185 83.750 151.405 ;
        RECT 83.395 150.595 83.565 151.185 ;
        RECT 83.920 150.985 84.090 151.695 ;
        RECT 84.965 151.625 85.295 152.085 ;
        RECT 85.505 151.725 85.855 151.895 ;
        RECT 84.295 151.155 85.085 151.405 ;
        RECT 85.505 151.335 85.765 151.725 ;
        RECT 86.075 151.635 87.025 151.915 ;
        RECT 87.195 151.645 87.385 152.085 ;
        RECT 87.555 151.705 88.625 151.875 ;
        RECT 85.255 150.985 85.425 151.165 ;
        RECT 82.535 150.165 82.930 150.335 ;
        RECT 83.100 150.205 83.565 150.595 ;
        RECT 83.735 150.815 85.425 150.985 ;
        RECT 82.760 150.035 82.930 150.165 ;
        RECT 83.735 150.035 83.905 150.815 ;
        RECT 85.595 150.645 85.765 151.335 ;
        RECT 84.265 150.475 85.765 150.645 ;
        RECT 85.955 150.675 86.165 151.465 ;
        RECT 86.335 150.845 86.685 151.465 ;
        RECT 86.855 150.855 87.025 151.635 ;
        RECT 87.555 151.475 87.725 151.705 ;
        RECT 87.195 151.305 87.725 151.475 ;
        RECT 87.195 151.025 87.415 151.305 ;
        RECT 87.895 151.135 88.135 151.535 ;
        RECT 86.855 150.685 87.260 150.855 ;
        RECT 87.595 150.765 88.135 151.135 ;
        RECT 88.305 151.350 88.625 151.705 ;
        RECT 88.870 151.625 89.175 152.085 ;
        RECT 89.345 151.375 89.600 151.905 ;
        RECT 88.305 151.175 88.630 151.350 ;
        RECT 88.305 150.875 89.220 151.175 ;
        RECT 88.480 150.845 89.220 150.875 ;
        RECT 85.955 150.515 86.630 150.675 ;
        RECT 87.090 150.595 87.260 150.685 ;
        RECT 85.955 150.505 86.920 150.515 ;
        RECT 85.595 150.335 85.765 150.475 ;
        RECT 82.340 149.535 82.590 149.995 ;
        RECT 82.760 149.705 83.010 150.035 ;
        RECT 83.225 149.705 83.905 150.035 ;
        RECT 84.075 150.135 85.150 150.305 ;
        RECT 85.595 150.165 86.155 150.335 ;
        RECT 86.460 150.215 86.920 150.505 ;
        RECT 87.090 150.425 88.310 150.595 ;
        RECT 84.075 149.795 84.245 150.135 ;
        RECT 84.480 149.535 84.810 149.965 ;
        RECT 84.980 149.795 85.150 150.135 ;
        RECT 85.445 149.535 85.815 149.995 ;
        RECT 85.985 149.705 86.155 150.165 ;
        RECT 87.090 150.045 87.260 150.425 ;
        RECT 88.480 150.255 88.650 150.845 ;
        RECT 89.390 150.725 89.600 151.375 ;
        RECT 86.390 149.705 87.260 150.045 ;
        RECT 87.850 150.085 88.650 150.255 ;
        RECT 87.430 149.535 87.680 149.995 ;
        RECT 87.850 149.795 88.020 150.085 ;
        RECT 88.200 149.535 88.530 149.915 ;
        RECT 88.870 149.535 89.175 150.675 ;
        RECT 89.345 149.845 89.600 150.725 ;
        RECT 89.780 151.545 90.035 151.875 ;
        RECT 90.205 151.705 90.535 152.085 ;
        RECT 91.665 151.705 92.920 151.875 ;
        RECT 93.105 151.705 93.435 152.085 ;
        RECT 89.780 150.675 89.950 151.545 ;
        RECT 90.260 151.365 92.540 151.535 ;
        RECT 90.260 151.175 90.430 151.365 ;
        RECT 92.370 151.175 92.540 151.365 ;
        RECT 92.750 151.515 92.920 151.705 ;
        RECT 93.605 151.535 93.775 151.915 ;
        RECT 93.945 151.705 94.275 152.085 ;
        RECT 94.445 151.535 94.615 151.915 ;
        RECT 94.785 151.705 95.115 152.085 ;
        RECT 92.750 151.345 93.425 151.515 ;
        RECT 93.605 151.365 95.120 151.535 ;
        RECT 90.120 150.845 90.430 151.175 ;
        RECT 90.600 150.675 90.770 151.175 ;
        RECT 89.780 150.505 90.770 150.675 ;
        RECT 91.170 150.555 91.440 151.175 ;
        RECT 91.655 150.845 92.125 151.175 ;
        RECT 92.370 150.845 93.085 151.175 ;
        RECT 93.255 151.095 93.425 151.345 ;
        RECT 93.255 150.925 94.720 151.095 ;
        RECT 93.255 150.575 93.425 150.925 ;
        RECT 94.890 150.595 95.120 151.365 ;
        RECT 89.780 149.705 90.035 150.505 ;
        RECT 91.670 150.405 93.425 150.575 ;
        RECT 93.255 150.385 93.425 150.405 ;
        RECT 93.605 150.425 95.120 150.595 ;
        RECT 90.205 149.535 90.510 150.335 ;
        RECT 90.680 149.895 91.030 150.235 ;
        RECT 91.220 150.065 92.935 150.235 ;
        RECT 90.680 149.725 92.460 149.895 ;
        RECT 92.765 149.705 92.935 150.065 ;
        RECT 93.105 149.535 93.435 149.915 ;
        RECT 93.605 149.705 93.775 150.425 ;
        RECT 93.945 149.535 94.275 150.255 ;
        RECT 94.445 149.705 94.615 150.425 ;
        RECT 94.785 149.535 95.115 150.255 ;
        RECT 96.215 149.705 96.965 151.915 ;
        RECT 98.060 151.285 98.315 152.085 ;
        RECT 98.485 151.420 98.735 151.915 ;
        RECT 98.905 151.705 99.235 152.085 ;
        RECT 99.405 151.705 100.700 151.875 ;
        RECT 99.405 151.535 99.575 151.705 ;
        RECT 98.060 149.535 98.315 150.675 ;
        RECT 98.485 150.575 98.655 151.420 ;
        RECT 98.965 151.365 99.575 151.535 ;
        RECT 100.870 151.435 101.060 151.750 ;
        RECT 101.320 151.585 101.520 152.085 ;
        RECT 98.965 151.175 99.135 151.365 ;
        RECT 98.825 150.845 99.135 151.175 ;
        RECT 98.485 149.705 98.795 150.575 ;
        RECT 98.965 150.335 99.135 150.845 ;
        RECT 99.305 150.675 99.475 151.175 ;
        RECT 99.785 150.890 100.415 151.405 ;
        RECT 100.595 151.145 101.060 151.435 ;
        RECT 100.245 150.855 100.415 150.890 ;
        RECT 99.305 150.505 99.965 150.675 ;
        RECT 100.245 150.545 101.060 150.855 ;
        RECT 101.330 150.545 101.520 151.415 ;
        RECT 99.795 150.335 99.965 150.505 ;
        RECT 101.690 150.335 102.020 151.915 ;
        RECT 102.360 151.575 102.600 152.085 ;
        RECT 102.780 151.575 103.060 151.905 ;
        RECT 103.290 151.575 103.505 152.085 ;
        RECT 102.255 150.845 102.610 151.405 ;
        RECT 102.780 150.675 102.950 151.575 ;
        RECT 103.120 150.845 103.385 151.405 ;
        RECT 103.675 151.345 104.290 151.915 ;
        RECT 103.635 150.675 103.805 151.175 ;
        RECT 98.965 150.165 99.625 150.335 ;
        RECT 99.795 150.165 102.020 150.335 ;
        RECT 102.380 150.505 103.805 150.675 ;
        RECT 102.380 150.330 102.770 150.505 ;
        RECT 98.995 149.535 99.285 149.995 ;
        RECT 99.455 149.915 99.625 150.165 ;
        RECT 99.455 149.745 100.765 149.915 ;
        RECT 101.295 149.535 101.515 149.995 ;
        RECT 101.685 149.705 102.020 150.165 ;
        RECT 103.255 149.535 103.585 150.335 ;
        RECT 103.975 150.325 104.290 151.345 ;
        RECT 104.495 151.335 105.705 152.085 ;
        RECT 105.875 151.360 106.165 152.085 ;
        RECT 104.495 150.795 105.015 151.335 ;
        RECT 105.185 150.625 105.705 151.165 ;
        RECT 103.755 149.705 104.290 150.325 ;
        RECT 104.495 149.535 105.705 150.625 ;
        RECT 105.875 149.535 106.165 150.700 ;
        RECT 107.255 149.705 108.005 151.915 ;
        RECT 108.420 151.725 110.440 151.915 ;
        RECT 110.610 151.725 110.940 152.085 ;
        RECT 111.470 151.725 111.800 152.085 ;
        RECT 112.330 151.725 112.660 152.085 ;
        RECT 113.190 151.725 113.520 152.085 ;
        RECT 110.210 151.555 110.440 151.725 ;
        RECT 114.320 151.575 114.560 152.085 ;
        RECT 114.740 151.575 115.020 151.905 ;
        RECT 115.250 151.575 115.465 152.085 ;
        RECT 108.235 151.325 110.040 151.555 ;
        RECT 110.210 151.350 113.950 151.555 ;
        RECT 108.235 150.725 108.645 151.325 ;
        RECT 108.815 150.895 110.165 151.155 ;
        RECT 108.235 150.470 110.135 150.725 ;
        RECT 110.375 150.655 110.625 151.180 ;
        RECT 110.795 150.825 112.085 151.100 ;
        RECT 112.595 150.850 113.945 151.155 ;
        RECT 112.595 150.655 113.495 150.850 ;
        RECT 114.215 150.845 114.570 151.405 ;
        RECT 114.740 150.675 114.910 151.575 ;
        RECT 115.080 150.845 115.345 151.405 ;
        RECT 115.635 151.345 116.250 151.915 ;
        RECT 115.595 150.675 115.765 151.175 ;
        RECT 110.375 150.485 113.495 150.655 ;
        RECT 114.340 150.505 115.765 150.675 ;
        RECT 108.920 150.315 110.135 150.470 ;
        RECT 108.420 149.535 108.750 150.290 ;
        RECT 108.920 150.145 112.230 150.315 ;
        RECT 108.920 150.085 109.990 150.145 ;
        RECT 108.920 149.705 109.110 150.085 ;
        RECT 109.280 149.535 109.610 149.915 ;
        RECT 109.780 149.705 109.990 150.085 ;
        RECT 112.400 150.085 113.495 150.255 ;
        RECT 110.160 149.535 110.440 149.975 ;
        RECT 112.400 149.895 112.590 150.085 ;
        RECT 110.610 149.705 112.590 149.895 ;
        RECT 112.760 149.535 113.090 149.915 ;
        RECT 113.260 149.705 113.495 150.085 ;
        RECT 113.665 149.535 113.950 150.350 ;
        RECT 114.340 150.330 114.730 150.505 ;
        RECT 115.215 149.535 115.545 150.335 ;
        RECT 115.935 150.325 116.250 151.345 ;
        RECT 116.505 151.330 116.755 152.085 ;
        RECT 116.925 151.375 117.175 151.905 ;
        RECT 117.345 151.625 117.650 152.085 ;
        RECT 117.895 151.705 118.965 151.875 ;
        RECT 116.925 150.725 117.130 151.375 ;
        RECT 117.895 151.350 118.215 151.705 ;
        RECT 117.890 151.175 118.215 151.350 ;
        RECT 117.300 150.875 118.215 151.175 ;
        RECT 118.385 151.135 118.625 151.535 ;
        RECT 118.795 151.475 118.965 151.705 ;
        RECT 119.135 151.645 119.325 152.085 ;
        RECT 119.495 151.635 120.445 151.915 ;
        RECT 120.665 151.725 121.015 151.895 ;
        RECT 118.795 151.305 119.325 151.475 ;
        RECT 117.300 150.845 118.040 150.875 ;
        RECT 115.715 149.705 116.250 150.325 ;
        RECT 116.505 149.535 116.755 150.675 ;
        RECT 116.925 149.845 117.175 150.725 ;
        RECT 117.345 149.535 117.650 150.675 ;
        RECT 117.870 150.255 118.040 150.845 ;
        RECT 118.385 150.765 118.925 151.135 ;
        RECT 119.105 151.025 119.325 151.305 ;
        RECT 119.495 150.855 119.665 151.635 ;
        RECT 119.260 150.685 119.665 150.855 ;
        RECT 119.835 150.845 120.185 151.465 ;
        RECT 119.260 150.595 119.430 150.685 ;
        RECT 120.355 150.675 120.565 151.465 ;
        RECT 118.210 150.425 119.430 150.595 ;
        RECT 119.890 150.515 120.565 150.675 ;
        RECT 117.870 150.085 118.670 150.255 ;
        RECT 117.990 149.535 118.320 149.915 ;
        RECT 118.500 149.795 118.670 150.085 ;
        RECT 119.260 150.045 119.430 150.425 ;
        RECT 119.600 150.505 120.565 150.515 ;
        RECT 120.755 151.335 121.015 151.725 ;
        RECT 121.225 151.625 121.555 152.085 ;
        RECT 122.430 151.695 123.285 151.865 ;
        RECT 123.490 151.695 123.985 151.865 ;
        RECT 124.155 151.725 124.485 152.085 ;
        RECT 120.755 150.645 120.925 151.335 ;
        RECT 121.095 150.985 121.265 151.165 ;
        RECT 121.435 151.155 122.225 151.405 ;
        RECT 122.430 150.985 122.600 151.695 ;
        RECT 122.770 151.185 123.125 151.405 ;
        RECT 121.095 150.815 122.785 150.985 ;
        RECT 119.600 150.215 120.060 150.505 ;
        RECT 120.755 150.475 122.255 150.645 ;
        RECT 120.755 150.335 120.925 150.475 ;
        RECT 120.365 150.165 120.925 150.335 ;
        RECT 118.840 149.535 119.090 149.995 ;
        RECT 119.260 149.705 120.130 150.045 ;
        RECT 120.365 149.705 120.535 150.165 ;
        RECT 121.370 150.135 122.445 150.305 ;
        RECT 120.705 149.535 121.075 149.995 ;
        RECT 121.370 149.795 121.540 150.135 ;
        RECT 121.710 149.535 122.040 149.965 ;
        RECT 122.275 149.795 122.445 150.135 ;
        RECT 122.615 150.035 122.785 150.815 ;
        RECT 122.955 150.595 123.125 151.185 ;
        RECT 123.295 150.785 123.645 151.405 ;
        RECT 122.955 150.205 123.420 150.595 ;
        RECT 123.815 150.335 123.985 151.695 ;
        RECT 124.155 150.505 124.615 151.555 ;
        RECT 123.590 150.165 123.985 150.335 ;
        RECT 123.590 150.035 123.760 150.165 ;
        RECT 122.615 149.705 123.295 150.035 ;
        RECT 123.510 149.705 123.760 150.035 ;
        RECT 123.930 149.535 124.180 149.995 ;
        RECT 124.350 149.720 124.675 150.505 ;
        RECT 124.845 149.705 125.015 151.825 ;
        RECT 125.185 151.705 125.515 152.085 ;
        RECT 125.685 151.535 125.940 151.825 ;
        RECT 125.190 151.365 125.940 151.535 ;
        RECT 125.190 150.375 125.420 151.365 ;
        RECT 126.115 151.285 126.425 152.085 ;
        RECT 126.630 151.285 127.325 151.915 ;
        RECT 125.590 150.545 125.940 151.195 ;
        RECT 126.125 150.845 126.460 151.115 ;
        RECT 126.630 150.685 126.800 151.285 ;
        RECT 127.770 151.275 128.015 151.880 ;
        RECT 128.235 151.550 128.745 152.085 ;
        RECT 127.495 151.105 128.725 151.275 ;
        RECT 126.970 150.845 127.305 151.095 ;
        RECT 125.190 150.205 125.940 150.375 ;
        RECT 125.185 149.535 125.515 150.035 ;
        RECT 125.685 149.705 125.940 150.205 ;
        RECT 126.115 149.535 126.395 150.675 ;
        RECT 126.565 149.705 126.895 150.685 ;
        RECT 127.065 149.535 127.325 150.675 ;
        RECT 127.495 150.295 127.835 151.105 ;
        RECT 128.005 150.540 128.755 150.730 ;
        RECT 127.495 149.885 128.010 150.295 ;
        RECT 128.245 149.535 128.415 150.295 ;
        RECT 128.585 149.875 128.755 150.540 ;
        RECT 128.925 150.555 129.115 151.915 ;
        RECT 129.285 151.065 129.560 151.915 ;
        RECT 129.750 151.550 130.280 151.915 ;
        RECT 130.705 151.685 131.035 152.085 ;
        RECT 130.105 151.515 130.280 151.550 ;
        RECT 129.285 150.895 129.565 151.065 ;
        RECT 129.285 150.755 129.560 150.895 ;
        RECT 129.765 150.555 129.935 151.355 ;
        RECT 128.925 150.385 129.935 150.555 ;
        RECT 130.105 151.345 131.035 151.515 ;
        RECT 131.205 151.345 131.460 151.915 ;
        RECT 131.635 151.360 131.925 152.085 ;
        RECT 132.560 151.535 132.815 151.825 ;
        RECT 132.985 151.705 133.315 152.085 ;
        RECT 132.560 151.365 133.310 151.535 ;
        RECT 130.105 150.215 130.275 151.345 ;
        RECT 130.865 151.175 131.035 151.345 ;
        RECT 129.150 150.045 130.275 150.215 ;
        RECT 130.445 150.845 130.640 151.175 ;
        RECT 130.865 150.845 131.120 151.175 ;
        RECT 130.445 149.875 130.615 150.845 ;
        RECT 131.290 150.675 131.460 151.345 ;
        RECT 128.585 149.705 130.615 149.875 ;
        RECT 130.785 149.535 130.955 150.675 ;
        RECT 131.125 149.705 131.460 150.675 ;
        RECT 131.635 149.535 131.925 150.700 ;
        RECT 132.560 150.545 132.910 151.195 ;
        RECT 133.080 150.375 133.310 151.365 ;
        RECT 132.560 150.205 133.310 150.375 ;
        RECT 132.560 149.705 132.815 150.205 ;
        RECT 132.985 149.535 133.315 150.035 ;
        RECT 133.485 149.705 133.655 151.825 ;
        RECT 134.015 151.725 134.345 152.085 ;
        RECT 134.515 151.695 135.010 151.865 ;
        RECT 135.215 151.695 136.070 151.865 ;
        RECT 133.885 150.505 134.345 151.555 ;
        RECT 133.825 149.720 134.150 150.505 ;
        RECT 134.515 150.335 134.685 151.695 ;
        RECT 134.855 150.785 135.205 151.405 ;
        RECT 135.375 151.185 135.730 151.405 ;
        RECT 135.375 150.595 135.545 151.185 ;
        RECT 135.900 150.985 136.070 151.695 ;
        RECT 136.945 151.625 137.275 152.085 ;
        RECT 137.485 151.725 137.835 151.895 ;
        RECT 136.275 151.155 137.065 151.405 ;
        RECT 137.485 151.335 137.745 151.725 ;
        RECT 138.055 151.635 139.005 151.915 ;
        RECT 139.175 151.645 139.365 152.085 ;
        RECT 139.535 151.705 140.605 151.875 ;
        RECT 137.235 150.985 137.405 151.165 ;
        RECT 134.515 150.165 134.910 150.335 ;
        RECT 135.080 150.205 135.545 150.595 ;
        RECT 135.715 150.815 137.405 150.985 ;
        RECT 134.740 150.035 134.910 150.165 ;
        RECT 135.715 150.035 135.885 150.815 ;
        RECT 137.575 150.645 137.745 151.335 ;
        RECT 136.245 150.475 137.745 150.645 ;
        RECT 137.935 150.675 138.145 151.465 ;
        RECT 138.315 150.845 138.665 151.465 ;
        RECT 138.835 150.855 139.005 151.635 ;
        RECT 139.535 151.475 139.705 151.705 ;
        RECT 139.175 151.305 139.705 151.475 ;
        RECT 139.175 151.025 139.395 151.305 ;
        RECT 139.875 151.135 140.115 151.535 ;
        RECT 138.835 150.685 139.240 150.855 ;
        RECT 139.575 150.765 140.115 151.135 ;
        RECT 140.285 151.350 140.605 151.705 ;
        RECT 140.850 151.625 141.155 152.085 ;
        RECT 141.325 151.375 141.580 151.905 ;
        RECT 141.815 151.605 142.095 152.085 ;
        RECT 142.265 151.435 142.525 151.825 ;
        RECT 142.700 151.605 142.955 152.085 ;
        RECT 143.125 151.435 143.420 151.825 ;
        RECT 143.600 151.605 143.875 152.085 ;
        RECT 144.045 151.585 144.345 151.915 ;
        RECT 140.285 151.175 140.610 151.350 ;
        RECT 140.285 150.875 141.200 151.175 ;
        RECT 140.460 150.845 141.200 150.875 ;
        RECT 137.935 150.515 138.610 150.675 ;
        RECT 139.070 150.595 139.240 150.685 ;
        RECT 137.935 150.505 138.900 150.515 ;
        RECT 137.575 150.335 137.745 150.475 ;
        RECT 134.320 149.535 134.570 149.995 ;
        RECT 134.740 149.705 134.990 150.035 ;
        RECT 135.205 149.705 135.885 150.035 ;
        RECT 136.055 150.135 137.130 150.305 ;
        RECT 137.575 150.165 138.135 150.335 ;
        RECT 138.440 150.215 138.900 150.505 ;
        RECT 139.070 150.425 140.290 150.595 ;
        RECT 136.055 149.795 136.225 150.135 ;
        RECT 136.460 149.535 136.790 149.965 ;
        RECT 136.960 149.795 137.130 150.135 ;
        RECT 137.425 149.535 137.795 149.995 ;
        RECT 137.965 149.705 138.135 150.165 ;
        RECT 139.070 150.045 139.240 150.425 ;
        RECT 140.460 150.255 140.630 150.845 ;
        RECT 141.370 150.725 141.580 151.375 ;
        RECT 138.370 149.705 139.240 150.045 ;
        RECT 139.830 150.085 140.630 150.255 ;
        RECT 139.410 149.535 139.660 149.995 ;
        RECT 139.830 149.795 140.000 150.085 ;
        RECT 140.180 149.535 140.510 149.915 ;
        RECT 140.850 149.535 141.155 150.675 ;
        RECT 141.325 149.845 141.580 150.725 ;
        RECT 141.770 151.265 143.420 151.435 ;
        RECT 141.770 150.755 142.175 151.265 ;
        RECT 142.345 150.925 143.485 151.095 ;
        RECT 141.770 150.585 142.525 150.755 ;
        RECT 141.810 149.535 142.095 150.405 ;
        RECT 142.265 150.335 142.525 150.585 ;
        RECT 143.315 150.675 143.485 150.925 ;
        RECT 143.655 150.845 144.005 151.415 ;
        RECT 144.175 150.675 144.345 151.585 ;
        RECT 144.515 151.540 149.860 152.085 ;
        RECT 150.035 151.540 155.380 152.085 ;
        RECT 146.100 150.710 146.440 151.540 ;
        RECT 143.315 150.505 144.345 150.675 ;
        RECT 142.265 150.165 143.385 150.335 ;
        RECT 142.265 149.705 142.525 150.165 ;
        RECT 142.700 149.535 142.955 149.995 ;
        RECT 143.125 149.705 143.385 150.165 ;
        RECT 143.555 149.535 143.865 150.335 ;
        RECT 144.035 149.705 144.345 150.505 ;
        RECT 147.920 149.970 148.270 151.220 ;
        RECT 151.620 150.710 151.960 151.540 ;
        RECT 155.555 151.335 156.765 152.085 ;
        RECT 156.935 151.335 158.145 152.085 ;
        RECT 153.440 149.970 153.790 151.220 ;
        RECT 155.555 150.795 156.075 151.335 ;
        RECT 156.245 150.625 156.765 151.165 ;
        RECT 144.515 149.535 149.860 149.970 ;
        RECT 150.035 149.535 155.380 149.970 ;
        RECT 155.555 149.535 156.765 150.625 ;
        RECT 156.935 150.625 157.455 151.165 ;
        RECT 157.625 150.795 158.145 151.335 ;
        RECT 156.935 149.535 158.145 150.625 ;
        RECT 2.750 149.365 158.230 149.535 ;
        RECT 2.835 148.275 4.045 149.365 ;
        RECT 4.220 148.695 4.475 149.195 ;
        RECT 4.645 148.865 4.975 149.365 ;
        RECT 4.220 148.525 4.970 148.695 ;
        RECT 2.835 147.565 3.355 148.105 ;
        RECT 3.525 147.735 4.045 148.275 ;
        RECT 4.220 147.705 4.570 148.355 ;
        RECT 2.835 146.815 4.045 147.565 ;
        RECT 4.740 147.535 4.970 148.525 ;
        RECT 4.220 147.365 4.970 147.535 ;
        RECT 4.220 147.075 4.475 147.365 ;
        RECT 4.645 146.815 4.975 147.195 ;
        RECT 5.145 147.075 5.315 149.195 ;
        RECT 5.485 148.395 5.810 149.180 ;
        RECT 5.980 148.905 6.230 149.365 ;
        RECT 6.400 148.865 6.650 149.195 ;
        RECT 6.865 148.865 7.545 149.195 ;
        RECT 6.400 148.735 6.570 148.865 ;
        RECT 6.175 148.565 6.570 148.735 ;
        RECT 5.545 147.345 6.005 148.395 ;
        RECT 6.175 147.205 6.345 148.565 ;
        RECT 6.740 148.305 7.205 148.695 ;
        RECT 6.515 147.495 6.865 148.115 ;
        RECT 7.035 147.715 7.205 148.305 ;
        RECT 7.375 148.085 7.545 148.865 ;
        RECT 7.715 148.765 7.885 149.105 ;
        RECT 8.120 148.935 8.450 149.365 ;
        RECT 8.620 148.765 8.790 149.105 ;
        RECT 9.085 148.905 9.455 149.365 ;
        RECT 7.715 148.595 8.790 148.765 ;
        RECT 9.625 148.735 9.795 149.195 ;
        RECT 10.030 148.855 10.900 149.195 ;
        RECT 11.070 148.905 11.320 149.365 ;
        RECT 9.235 148.565 9.795 148.735 ;
        RECT 9.235 148.425 9.405 148.565 ;
        RECT 7.905 148.255 9.405 148.425 ;
        RECT 10.100 148.395 10.560 148.685 ;
        RECT 7.375 147.915 9.065 148.085 ;
        RECT 7.035 147.495 7.390 147.715 ;
        RECT 7.560 147.205 7.730 147.915 ;
        RECT 7.935 147.495 8.725 147.745 ;
        RECT 8.895 147.735 9.065 147.915 ;
        RECT 9.235 147.565 9.405 148.255 ;
        RECT 5.675 146.815 6.005 147.175 ;
        RECT 6.175 147.035 6.670 147.205 ;
        RECT 6.875 147.035 7.730 147.205 ;
        RECT 8.605 146.815 8.935 147.275 ;
        RECT 9.145 147.175 9.405 147.565 ;
        RECT 9.595 148.385 10.560 148.395 ;
        RECT 10.730 148.475 10.900 148.855 ;
        RECT 11.490 148.815 11.660 149.105 ;
        RECT 11.840 148.985 12.170 149.365 ;
        RECT 11.490 148.645 12.290 148.815 ;
        RECT 9.595 148.225 10.270 148.385 ;
        RECT 10.730 148.305 11.950 148.475 ;
        RECT 9.595 147.435 9.805 148.225 ;
        RECT 10.730 148.215 10.900 148.305 ;
        RECT 9.975 147.435 10.325 148.055 ;
        RECT 10.495 148.045 10.900 148.215 ;
        RECT 10.495 147.265 10.665 148.045 ;
        RECT 10.835 147.595 11.055 147.875 ;
        RECT 11.235 147.765 11.775 148.135 ;
        RECT 12.120 148.055 12.290 148.645 ;
        RECT 12.510 148.225 12.815 149.365 ;
        RECT 12.985 148.175 13.240 149.055 ;
        RECT 12.120 148.025 12.860 148.055 ;
        RECT 10.835 147.425 11.365 147.595 ;
        RECT 9.145 147.005 9.495 147.175 ;
        RECT 9.715 146.985 10.665 147.265 ;
        RECT 10.835 146.815 11.025 147.255 ;
        RECT 11.195 147.195 11.365 147.425 ;
        RECT 11.535 147.365 11.775 147.765 ;
        RECT 11.945 147.725 12.860 148.025 ;
        RECT 11.945 147.550 12.270 147.725 ;
        RECT 11.945 147.195 12.265 147.550 ;
        RECT 13.030 147.525 13.240 148.175 ;
        RECT 11.195 147.025 12.265 147.195 ;
        RECT 12.510 146.815 12.815 147.275 ;
        RECT 12.985 146.995 13.240 147.525 ;
        RECT 13.415 148.290 13.685 149.195 ;
        RECT 13.855 148.605 14.185 149.365 ;
        RECT 14.365 148.435 14.535 149.195 ;
        RECT 13.415 147.490 13.585 148.290 ;
        RECT 13.870 148.265 14.535 148.435 ;
        RECT 13.870 148.120 14.040 148.265 ;
        RECT 15.715 148.200 16.005 149.365 ;
        RECT 16.180 148.225 16.515 149.195 ;
        RECT 16.685 148.225 16.855 149.365 ;
        RECT 17.025 149.025 19.055 149.195 ;
        RECT 13.755 147.790 14.040 148.120 ;
        RECT 13.870 147.535 14.040 147.790 ;
        RECT 14.275 147.715 14.605 148.085 ;
        RECT 16.180 147.555 16.350 148.225 ;
        RECT 17.025 148.055 17.195 149.025 ;
        RECT 16.520 147.725 16.775 148.055 ;
        RECT 17.000 147.725 17.195 148.055 ;
        RECT 17.365 148.685 18.490 148.855 ;
        RECT 16.605 147.555 16.775 147.725 ;
        RECT 17.365 147.555 17.535 148.685 ;
        RECT 13.415 146.985 13.675 147.490 ;
        RECT 13.870 147.365 14.535 147.535 ;
        RECT 13.855 146.815 14.185 147.195 ;
        RECT 14.365 146.985 14.535 147.365 ;
        RECT 15.715 146.815 16.005 147.540 ;
        RECT 16.180 146.985 16.435 147.555 ;
        RECT 16.605 147.385 17.535 147.555 ;
        RECT 17.705 148.345 18.715 148.515 ;
        RECT 17.705 147.545 17.875 148.345 ;
        RECT 17.360 147.350 17.535 147.385 ;
        RECT 16.605 146.815 16.935 147.215 ;
        RECT 17.360 146.985 17.890 147.350 ;
        RECT 18.080 147.325 18.355 148.145 ;
        RECT 18.075 147.155 18.355 147.325 ;
        RECT 18.080 146.985 18.355 147.155 ;
        RECT 18.525 146.985 18.715 148.345 ;
        RECT 18.885 148.360 19.055 149.025 ;
        RECT 19.225 148.605 19.395 149.365 ;
        RECT 19.630 148.605 20.145 149.015 ;
        RECT 18.885 148.170 19.635 148.360 ;
        RECT 19.805 147.795 20.145 148.605 ;
        RECT 18.915 147.625 20.145 147.795 ;
        RECT 20.315 148.225 20.700 149.195 ;
        RECT 20.870 148.905 21.195 149.365 ;
        RECT 21.715 148.735 21.995 149.195 ;
        RECT 20.870 148.515 21.995 148.735 ;
        RECT 18.895 146.815 19.405 147.350 ;
        RECT 19.625 147.020 19.870 147.625 ;
        RECT 20.315 147.555 20.595 148.225 ;
        RECT 20.870 148.055 21.320 148.515 ;
        RECT 22.185 148.345 22.585 149.195 ;
        RECT 22.985 148.905 23.255 149.365 ;
        RECT 23.425 148.735 23.710 149.195 ;
        RECT 20.765 147.725 21.320 148.055 ;
        RECT 21.490 147.785 22.585 148.345 ;
        RECT 20.870 147.615 21.320 147.725 ;
        RECT 20.315 146.985 20.700 147.555 ;
        RECT 20.870 147.445 21.995 147.615 ;
        RECT 20.870 146.815 21.195 147.275 ;
        RECT 21.715 146.985 21.995 147.445 ;
        RECT 22.185 146.985 22.585 147.785 ;
        RECT 22.755 148.515 23.710 148.735 ;
        RECT 22.755 147.615 22.965 148.515 ;
        RECT 23.135 147.785 23.825 148.345 ;
        RECT 23.995 148.290 24.265 149.195 ;
        RECT 24.435 148.605 24.765 149.365 ;
        RECT 24.945 148.435 25.115 149.195 ;
        RECT 22.755 147.445 23.710 147.615 ;
        RECT 22.985 146.815 23.255 147.275 ;
        RECT 23.425 146.985 23.710 147.445 ;
        RECT 23.995 147.490 24.165 148.290 ;
        RECT 24.450 148.265 25.115 148.435 ;
        RECT 25.840 148.975 26.175 149.195 ;
        RECT 27.180 148.985 27.535 149.365 ;
        RECT 25.840 148.355 26.095 148.975 ;
        RECT 26.345 148.815 26.575 148.855 ;
        RECT 27.705 148.815 27.955 149.195 ;
        RECT 26.345 148.615 27.955 148.815 ;
        RECT 26.345 148.525 26.530 148.615 ;
        RECT 27.120 148.605 27.955 148.615 ;
        RECT 28.205 148.585 28.455 149.365 ;
        RECT 28.625 148.515 28.885 149.195 ;
        RECT 26.685 148.415 27.015 148.445 ;
        RECT 26.685 148.355 28.485 148.415 ;
        RECT 24.450 148.120 24.620 148.265 ;
        RECT 25.840 148.245 28.545 148.355 ;
        RECT 25.840 148.185 27.015 148.245 ;
        RECT 28.345 148.210 28.545 148.245 ;
        RECT 24.335 147.790 24.620 148.120 ;
        RECT 24.450 147.535 24.620 147.790 ;
        RECT 24.855 147.715 25.185 148.085 ;
        RECT 25.835 147.805 26.325 148.005 ;
        RECT 26.515 147.805 26.990 148.015 ;
        RECT 23.995 146.985 24.255 147.490 ;
        RECT 24.450 147.365 25.115 147.535 ;
        RECT 24.435 146.815 24.765 147.195 ;
        RECT 24.945 146.985 25.115 147.365 ;
        RECT 25.840 146.815 26.295 147.580 ;
        RECT 26.770 147.405 26.990 147.805 ;
        RECT 27.235 147.805 27.565 148.015 ;
        RECT 27.235 147.405 27.445 147.805 ;
        RECT 27.735 147.770 28.145 148.075 ;
        RECT 28.375 147.635 28.545 148.210 ;
        RECT 28.275 147.515 28.545 147.635 ;
        RECT 27.700 147.470 28.545 147.515 ;
        RECT 27.700 147.345 28.455 147.470 ;
        RECT 27.700 147.195 27.870 147.345 ;
        RECT 28.715 147.315 28.885 148.515 ;
        RECT 29.060 148.975 29.395 149.195 ;
        RECT 30.400 148.985 30.755 149.365 ;
        RECT 29.060 148.355 29.315 148.975 ;
        RECT 29.565 148.815 29.795 148.855 ;
        RECT 30.925 148.815 31.175 149.195 ;
        RECT 29.565 148.615 31.175 148.815 ;
        RECT 29.565 148.525 29.750 148.615 ;
        RECT 30.340 148.605 31.175 148.615 ;
        RECT 31.425 148.585 31.675 149.365 ;
        RECT 31.845 148.515 32.105 149.195 ;
        RECT 29.905 148.415 30.235 148.445 ;
        RECT 29.905 148.355 31.705 148.415 ;
        RECT 29.060 148.245 31.765 148.355 ;
        RECT 29.060 148.185 30.235 148.245 ;
        RECT 31.565 148.210 31.765 148.245 ;
        RECT 29.055 147.805 29.545 148.005 ;
        RECT 29.735 147.805 30.210 148.015 ;
        RECT 26.570 146.985 27.870 147.195 ;
        RECT 28.125 146.815 28.455 147.175 ;
        RECT 28.625 146.985 28.885 147.315 ;
        RECT 29.060 146.815 29.515 147.580 ;
        RECT 29.990 147.405 30.210 147.805 ;
        RECT 30.455 147.805 30.785 148.015 ;
        RECT 30.455 147.405 30.665 147.805 ;
        RECT 30.955 147.770 31.365 148.075 ;
        RECT 31.595 147.635 31.765 148.210 ;
        RECT 31.495 147.515 31.765 147.635 ;
        RECT 30.920 147.470 31.765 147.515 ;
        RECT 30.920 147.345 31.675 147.470 ;
        RECT 30.920 147.195 31.090 147.345 ;
        RECT 31.935 147.315 32.105 148.515 ;
        RECT 32.305 148.175 32.555 149.365 ;
        RECT 29.790 146.985 31.090 147.195 ;
        RECT 31.345 146.815 31.675 147.175 ;
        RECT 31.845 146.985 32.105 147.315 ;
        RECT 32.375 146.815 32.545 147.615 ;
        RECT 32.780 147.095 32.995 149.195 ;
        RECT 33.185 148.605 33.985 149.365 ;
        RECT 34.380 148.435 34.765 149.195 ;
        RECT 33.165 148.225 34.765 148.435 ;
        RECT 35.090 148.345 35.290 149.135 ;
        RECT 35.460 148.525 35.780 149.365 ;
        RECT 35.955 148.395 36.225 149.165 ;
        RECT 36.395 148.585 36.725 149.365 ;
        RECT 36.930 148.760 37.115 149.165 ;
        RECT 37.285 148.940 37.620 149.365 ;
        RECT 36.930 148.585 37.595 148.760 ;
        RECT 33.165 147.625 33.445 148.225 ;
        RECT 34.935 148.175 35.290 148.345 ;
        RECT 34.935 148.055 35.115 148.175 ;
        RECT 33.625 147.805 33.980 148.055 ;
        RECT 34.150 147.805 34.615 148.055 ;
        RECT 34.785 147.805 35.115 148.055 ;
        RECT 35.460 148.005 35.780 148.345 ;
        RECT 35.285 147.805 35.780 148.005 ;
        RECT 35.955 148.225 37.085 148.395 ;
        RECT 33.165 147.445 34.405 147.625 ;
        RECT 34.750 147.555 35.780 147.595 ;
        RECT 34.040 147.375 34.405 147.445 ;
        RECT 34.580 147.425 35.780 147.555 ;
        RECT 33.215 146.815 33.395 147.275 ;
        RECT 34.580 147.205 34.920 147.425 ;
        RECT 33.655 147.025 34.920 147.205 ;
        RECT 35.105 146.815 35.275 147.255 ;
        RECT 35.445 147.010 35.780 147.425 ;
        RECT 35.955 147.315 36.125 148.225 ;
        RECT 36.295 147.475 36.655 148.055 ;
        RECT 36.835 147.725 37.085 148.225 ;
        RECT 37.255 147.555 37.595 148.585 ;
        RECT 36.910 147.385 37.595 147.555 ;
        RECT 37.815 148.525 38.070 149.195 ;
        RECT 38.240 148.605 38.570 149.365 ;
        RECT 38.740 148.765 38.990 149.195 ;
        RECT 39.160 148.945 39.515 149.365 ;
        RECT 39.705 149.025 40.875 149.195 ;
        RECT 39.705 148.985 40.035 149.025 ;
        RECT 40.145 148.765 40.375 148.855 ;
        RECT 38.740 148.525 40.375 148.765 ;
        RECT 40.545 148.525 40.875 149.025 ;
        RECT 37.815 147.395 37.985 148.525 ;
        RECT 41.045 148.355 41.215 149.195 ;
        RECT 38.155 148.185 41.215 148.355 ;
        RECT 41.475 148.200 41.765 149.365 ;
        RECT 41.975 149.025 43.115 149.195 ;
        RECT 41.975 148.565 42.275 149.025 ;
        RECT 42.445 148.395 42.775 148.855 ;
        RECT 38.155 147.635 38.325 148.185 ;
        RECT 42.015 148.175 42.775 148.395 ;
        RECT 42.945 148.395 43.115 149.025 ;
        RECT 43.285 148.565 43.615 149.365 ;
        RECT 43.785 148.395 44.060 149.195 ;
        RECT 42.945 148.185 44.060 148.395 ;
        RECT 44.325 148.355 44.495 149.195 ;
        RECT 44.665 149.025 45.835 149.195 ;
        RECT 44.665 148.525 44.995 149.025 ;
        RECT 45.505 148.985 45.835 149.025 ;
        RECT 46.025 148.945 46.380 149.365 ;
        RECT 45.165 148.765 45.395 148.855 ;
        RECT 46.550 148.765 46.800 149.195 ;
        RECT 45.165 148.525 46.800 148.765 ;
        RECT 46.970 148.605 47.300 149.365 ;
        RECT 47.470 148.525 47.725 149.195 ;
        RECT 47.515 148.515 47.725 148.525 ;
        RECT 44.325 148.185 47.385 148.355 ;
        RECT 38.545 147.835 38.920 148.005 ;
        RECT 38.555 147.805 38.920 147.835 ;
        RECT 39.090 147.805 39.420 148.005 ;
        RECT 38.155 147.465 38.955 147.635 ;
        RECT 35.955 146.985 36.215 147.315 ;
        RECT 36.425 146.815 36.700 147.295 ;
        RECT 36.910 146.985 37.115 147.385 ;
        RECT 37.815 147.325 38.000 147.395 ;
        RECT 37.815 147.315 38.025 147.325 ;
        RECT 37.285 146.815 37.620 147.215 ;
        RECT 37.815 146.985 38.070 147.315 ;
        RECT 38.285 146.815 38.615 147.295 ;
        RECT 38.785 147.235 38.955 147.465 ;
        RECT 39.135 147.405 39.420 147.805 ;
        RECT 39.690 147.805 40.165 148.005 ;
        RECT 40.335 147.805 40.780 148.005 ;
        RECT 40.950 147.805 41.300 148.015 ;
        RECT 39.690 147.405 39.970 147.805 ;
        RECT 42.015 147.635 42.230 148.175 ;
        RECT 42.400 147.805 43.170 148.005 ;
        RECT 43.340 147.805 44.060 148.005 ;
        RECT 44.240 147.805 44.590 148.015 ;
        RECT 44.760 147.805 45.205 148.005 ;
        RECT 45.375 147.805 45.850 148.005 ;
        RECT 40.150 147.465 41.215 147.635 ;
        RECT 40.150 147.235 40.320 147.465 ;
        RECT 38.785 146.985 40.320 147.235 ;
        RECT 40.545 146.815 40.875 147.295 ;
        RECT 41.045 146.985 41.215 147.465 ;
        RECT 41.475 146.815 41.765 147.540 ;
        RECT 42.015 147.465 43.615 147.635 ;
        RECT 42.445 147.455 43.615 147.465 ;
        RECT 41.985 146.815 42.275 147.285 ;
        RECT 42.445 146.985 42.775 147.455 ;
        RECT 42.945 146.815 43.115 147.285 ;
        RECT 43.285 146.985 43.615 147.455 ;
        RECT 43.785 146.815 44.060 147.635 ;
        RECT 44.325 147.465 45.390 147.635 ;
        RECT 44.325 146.985 44.495 147.465 ;
        RECT 44.665 146.815 44.995 147.295 ;
        RECT 45.220 147.235 45.390 147.465 ;
        RECT 45.570 147.405 45.850 147.805 ;
        RECT 46.120 147.805 46.450 148.005 ;
        RECT 46.620 147.805 46.985 148.005 ;
        RECT 46.120 147.405 46.405 147.805 ;
        RECT 47.215 147.635 47.385 148.185 ;
        RECT 46.585 147.465 47.385 147.635 ;
        RECT 46.585 147.235 46.755 147.465 ;
        RECT 47.555 147.395 47.725 148.515 ;
        RECT 47.945 148.175 48.195 149.365 ;
        RECT 47.540 147.315 47.725 147.395 ;
        RECT 45.220 146.985 46.755 147.235 ;
        RECT 46.925 146.815 47.255 147.295 ;
        RECT 47.470 146.985 47.725 147.315 ;
        RECT 48.015 146.815 48.185 147.615 ;
        RECT 48.420 147.095 48.635 149.195 ;
        RECT 48.825 148.605 49.625 149.365 ;
        RECT 50.020 148.435 50.405 149.195 ;
        RECT 48.805 148.225 50.405 148.435 ;
        RECT 50.730 148.345 50.930 149.135 ;
        RECT 51.100 148.525 51.420 149.365 ;
        RECT 48.805 147.625 49.085 148.225 ;
        RECT 50.575 148.175 50.930 148.345 ;
        RECT 50.575 148.055 50.755 148.175 ;
        RECT 49.265 147.805 49.620 148.055 ;
        RECT 49.790 147.805 50.255 148.055 ;
        RECT 50.425 147.805 50.755 148.055 ;
        RECT 51.100 148.005 51.420 148.345 ;
        RECT 51.625 148.175 51.875 149.365 ;
        RECT 50.925 147.805 51.420 148.005 ;
        RECT 48.805 147.445 50.045 147.625 ;
        RECT 50.390 147.555 51.420 147.595 ;
        RECT 49.680 147.375 50.045 147.445 ;
        RECT 50.220 147.425 51.420 147.555 ;
        RECT 48.855 146.815 49.035 147.275 ;
        RECT 50.220 147.205 50.560 147.425 ;
        RECT 49.295 147.025 50.560 147.205 ;
        RECT 50.745 146.815 50.915 147.255 ;
        RECT 51.085 147.010 51.420 147.425 ;
        RECT 51.695 146.815 51.865 147.615 ;
        RECT 52.100 147.095 52.315 149.195 ;
        RECT 52.505 148.605 53.305 149.365 ;
        RECT 53.700 148.435 54.085 149.195 ;
        RECT 52.485 148.225 54.085 148.435 ;
        RECT 54.410 148.345 54.610 149.135 ;
        RECT 54.780 148.525 55.100 149.365 ;
        RECT 55.275 148.855 56.465 149.145 ;
        RECT 55.295 148.515 56.465 148.685 ;
        RECT 56.635 148.565 56.915 149.365 ;
        RECT 52.485 147.625 52.765 148.225 ;
        RECT 54.255 148.175 54.610 148.345 ;
        RECT 54.255 148.055 54.435 148.175 ;
        RECT 52.945 147.805 53.300 148.055 ;
        RECT 53.470 147.805 53.935 148.055 ;
        RECT 54.105 147.805 54.435 148.055 ;
        RECT 54.780 148.005 55.100 148.345 ;
        RECT 55.295 148.225 55.620 148.515 ;
        RECT 56.295 148.395 56.465 148.515 ;
        RECT 55.790 148.055 55.985 148.345 ;
        RECT 56.295 148.225 56.955 148.395 ;
        RECT 57.125 148.225 57.400 149.195 ;
        RECT 56.785 148.055 56.955 148.225 ;
        RECT 54.605 147.805 55.100 148.005 ;
        RECT 55.275 147.725 55.620 148.055 ;
        RECT 55.790 147.725 56.615 148.055 ;
        RECT 56.785 147.725 57.060 148.055 ;
        RECT 52.485 147.445 53.725 147.625 ;
        RECT 54.070 147.555 55.100 147.595 ;
        RECT 56.785 147.555 56.955 147.725 ;
        RECT 53.360 147.375 53.725 147.445 ;
        RECT 53.900 147.425 55.100 147.555 ;
        RECT 52.535 146.815 52.715 147.275 ;
        RECT 53.900 147.205 54.240 147.425 ;
        RECT 52.975 147.025 54.240 147.205 ;
        RECT 54.425 146.815 54.595 147.255 ;
        RECT 54.765 147.010 55.100 147.425 ;
        RECT 55.290 147.385 56.955 147.555 ;
        RECT 57.230 147.490 57.400 148.225 ;
        RECT 55.290 147.035 55.545 147.385 ;
        RECT 55.715 146.815 56.045 147.215 ;
        RECT 56.215 147.035 56.385 147.385 ;
        RECT 56.555 146.815 56.935 147.215 ;
        RECT 57.125 147.145 57.400 147.490 ;
        RECT 57.580 148.175 57.835 149.055 ;
        RECT 58.005 148.225 58.310 149.365 ;
        RECT 58.650 148.985 58.980 149.365 ;
        RECT 59.160 148.815 59.330 149.105 ;
        RECT 59.500 148.905 59.750 149.365 ;
        RECT 58.530 148.645 59.330 148.815 ;
        RECT 59.920 148.855 60.790 149.195 ;
        RECT 57.580 147.525 57.790 148.175 ;
        RECT 58.530 148.055 58.700 148.645 ;
        RECT 59.920 148.475 60.090 148.855 ;
        RECT 61.025 148.735 61.195 149.195 ;
        RECT 61.365 148.905 61.735 149.365 ;
        RECT 62.030 148.765 62.200 149.105 ;
        RECT 62.370 148.935 62.700 149.365 ;
        RECT 62.935 148.765 63.105 149.105 ;
        RECT 58.870 148.305 60.090 148.475 ;
        RECT 60.260 148.395 60.720 148.685 ;
        RECT 61.025 148.565 61.585 148.735 ;
        RECT 62.030 148.595 63.105 148.765 ;
        RECT 63.275 148.865 63.955 149.195 ;
        RECT 64.170 148.865 64.420 149.195 ;
        RECT 64.590 148.905 64.840 149.365 ;
        RECT 61.415 148.425 61.585 148.565 ;
        RECT 60.260 148.385 61.225 148.395 ;
        RECT 59.920 148.215 60.090 148.305 ;
        RECT 60.550 148.225 61.225 148.385 ;
        RECT 57.960 148.025 58.700 148.055 ;
        RECT 57.960 147.725 58.875 148.025 ;
        RECT 58.550 147.550 58.875 147.725 ;
        RECT 57.580 146.995 57.835 147.525 ;
        RECT 58.005 146.815 58.310 147.275 ;
        RECT 58.555 147.195 58.875 147.550 ;
        RECT 59.045 147.765 59.585 148.135 ;
        RECT 59.920 148.045 60.325 148.215 ;
        RECT 59.045 147.365 59.285 147.765 ;
        RECT 59.765 147.595 59.985 147.875 ;
        RECT 59.455 147.425 59.985 147.595 ;
        RECT 59.455 147.195 59.625 147.425 ;
        RECT 60.155 147.265 60.325 148.045 ;
        RECT 60.495 147.435 60.845 148.055 ;
        RECT 61.015 147.435 61.225 148.225 ;
        RECT 61.415 148.255 62.915 148.425 ;
        RECT 61.415 147.565 61.585 148.255 ;
        RECT 63.275 148.085 63.445 148.865 ;
        RECT 64.250 148.735 64.420 148.865 ;
        RECT 61.755 147.915 63.445 148.085 ;
        RECT 63.615 148.305 64.080 148.695 ;
        RECT 64.250 148.565 64.645 148.735 ;
        RECT 61.755 147.735 61.925 147.915 ;
        RECT 58.555 147.025 59.625 147.195 ;
        RECT 59.795 146.815 59.985 147.255 ;
        RECT 60.155 146.985 61.105 147.265 ;
        RECT 61.415 147.175 61.675 147.565 ;
        RECT 62.095 147.495 62.885 147.745 ;
        RECT 61.325 147.005 61.675 147.175 ;
        RECT 61.885 146.815 62.215 147.275 ;
        RECT 63.090 147.205 63.260 147.915 ;
        RECT 63.615 147.715 63.785 148.305 ;
        RECT 63.430 147.495 63.785 147.715 ;
        RECT 63.955 147.495 64.305 148.115 ;
        RECT 64.475 147.205 64.645 148.565 ;
        RECT 65.010 148.395 65.335 149.180 ;
        RECT 64.815 147.345 65.275 148.395 ;
        RECT 63.090 147.035 63.945 147.205 ;
        RECT 64.150 147.035 64.645 147.205 ;
        RECT 64.815 146.815 65.145 147.175 ;
        RECT 65.505 147.075 65.675 149.195 ;
        RECT 65.845 148.865 66.175 149.365 ;
        RECT 66.345 148.695 66.600 149.195 ;
        RECT 65.850 148.525 66.600 148.695 ;
        RECT 65.850 147.535 66.080 148.525 ;
        RECT 66.250 147.705 66.600 148.355 ;
        RECT 67.235 148.200 67.525 149.365 ;
        RECT 67.695 148.290 67.965 149.195 ;
        RECT 68.135 148.605 68.465 149.365 ;
        RECT 68.645 148.435 68.815 149.195 ;
        RECT 69.080 148.695 69.335 149.195 ;
        RECT 69.505 148.865 69.835 149.365 ;
        RECT 69.080 148.525 69.830 148.695 ;
        RECT 65.850 147.365 66.600 147.535 ;
        RECT 65.845 146.815 66.175 147.195 ;
        RECT 66.345 147.075 66.600 147.365 ;
        RECT 67.235 146.815 67.525 147.540 ;
        RECT 67.695 147.490 67.865 148.290 ;
        RECT 68.150 148.265 68.815 148.435 ;
        RECT 68.150 148.120 68.320 148.265 ;
        RECT 68.035 147.790 68.320 148.120 ;
        RECT 68.150 147.535 68.320 147.790 ;
        RECT 68.555 147.715 68.885 148.085 ;
        RECT 69.080 147.705 69.430 148.355 ;
        RECT 69.600 147.535 69.830 148.525 ;
        RECT 67.695 146.985 67.955 147.490 ;
        RECT 68.150 147.365 68.815 147.535 ;
        RECT 68.135 146.815 68.465 147.195 ;
        RECT 68.645 146.985 68.815 147.365 ;
        RECT 69.080 147.365 69.830 147.535 ;
        RECT 69.080 147.075 69.335 147.365 ;
        RECT 69.505 146.815 69.835 147.195 ;
        RECT 70.005 147.075 70.175 149.195 ;
        RECT 70.345 148.395 70.670 149.180 ;
        RECT 70.840 148.905 71.090 149.365 ;
        RECT 71.260 148.865 71.510 149.195 ;
        RECT 71.725 148.865 72.405 149.195 ;
        RECT 71.260 148.735 71.430 148.865 ;
        RECT 71.035 148.565 71.430 148.735 ;
        RECT 70.405 147.345 70.865 148.395 ;
        RECT 71.035 147.205 71.205 148.565 ;
        RECT 71.600 148.305 72.065 148.695 ;
        RECT 71.375 147.495 71.725 148.115 ;
        RECT 71.895 147.715 72.065 148.305 ;
        RECT 72.235 148.085 72.405 148.865 ;
        RECT 72.575 148.765 72.745 149.105 ;
        RECT 72.980 148.935 73.310 149.365 ;
        RECT 73.480 148.765 73.650 149.105 ;
        RECT 73.945 148.905 74.315 149.365 ;
        RECT 72.575 148.595 73.650 148.765 ;
        RECT 74.485 148.735 74.655 149.195 ;
        RECT 74.890 148.855 75.760 149.195 ;
        RECT 75.930 148.905 76.180 149.365 ;
        RECT 74.095 148.565 74.655 148.735 ;
        RECT 74.095 148.425 74.265 148.565 ;
        RECT 72.765 148.255 74.265 148.425 ;
        RECT 74.960 148.395 75.420 148.685 ;
        RECT 72.235 147.915 73.925 148.085 ;
        RECT 71.895 147.495 72.250 147.715 ;
        RECT 72.420 147.205 72.590 147.915 ;
        RECT 72.795 147.495 73.585 147.745 ;
        RECT 73.755 147.735 73.925 147.915 ;
        RECT 74.095 147.565 74.265 148.255 ;
        RECT 70.535 146.815 70.865 147.175 ;
        RECT 71.035 147.035 71.530 147.205 ;
        RECT 71.735 147.035 72.590 147.205 ;
        RECT 73.465 146.815 73.795 147.275 ;
        RECT 74.005 147.175 74.265 147.565 ;
        RECT 74.455 148.385 75.420 148.395 ;
        RECT 75.590 148.475 75.760 148.855 ;
        RECT 76.350 148.815 76.520 149.105 ;
        RECT 76.700 148.985 77.030 149.365 ;
        RECT 76.350 148.645 77.150 148.815 ;
        RECT 74.455 148.225 75.130 148.385 ;
        RECT 75.590 148.305 76.810 148.475 ;
        RECT 74.455 147.435 74.665 148.225 ;
        RECT 75.590 148.215 75.760 148.305 ;
        RECT 74.835 147.435 75.185 148.055 ;
        RECT 75.355 148.045 75.760 148.215 ;
        RECT 75.355 147.265 75.525 148.045 ;
        RECT 75.695 147.595 75.915 147.875 ;
        RECT 76.095 147.765 76.635 148.135 ;
        RECT 76.980 148.055 77.150 148.645 ;
        RECT 77.370 148.225 77.675 149.365 ;
        RECT 77.845 148.175 78.100 149.055 ;
        RECT 78.280 148.225 78.535 149.365 ;
        RECT 78.705 148.325 79.015 149.195 ;
        RECT 79.215 148.905 79.505 149.365 ;
        RECT 79.675 148.985 80.985 149.155 ;
        RECT 79.675 148.735 79.845 148.985 ;
        RECT 81.515 148.905 81.735 149.365 ;
        RECT 81.905 148.735 82.240 149.195 ;
        RECT 79.185 148.565 79.845 148.735 ;
        RECT 80.015 148.565 82.240 148.735 ;
        RECT 76.980 148.025 77.720 148.055 ;
        RECT 75.695 147.425 76.225 147.595 ;
        RECT 74.005 147.005 74.355 147.175 ;
        RECT 74.575 146.985 75.525 147.265 ;
        RECT 75.695 146.815 75.885 147.255 ;
        RECT 76.055 147.195 76.225 147.425 ;
        RECT 76.395 147.365 76.635 147.765 ;
        RECT 76.805 147.725 77.720 148.025 ;
        RECT 76.805 147.550 77.130 147.725 ;
        RECT 76.805 147.195 77.125 147.550 ;
        RECT 77.890 147.525 78.100 148.175 ;
        RECT 76.055 147.025 77.125 147.195 ;
        RECT 77.370 146.815 77.675 147.275 ;
        RECT 77.845 146.995 78.100 147.525 ;
        RECT 78.280 146.815 78.535 147.615 ;
        RECT 78.705 147.480 78.875 148.325 ;
        RECT 79.185 148.055 79.355 148.565 ;
        RECT 80.015 148.395 80.185 148.565 ;
        RECT 79.045 147.725 79.355 148.055 ;
        RECT 79.525 148.225 80.185 148.395 ;
        RECT 79.525 147.725 79.695 148.225 ;
        RECT 80.465 148.045 81.280 148.355 ;
        RECT 80.465 148.010 80.635 148.045 ;
        RECT 79.185 147.535 79.355 147.725 ;
        RECT 78.705 146.985 78.955 147.480 ;
        RECT 79.185 147.365 79.795 147.535 ;
        RECT 80.005 147.495 80.635 148.010 ;
        RECT 80.815 147.465 81.280 147.755 ;
        RECT 81.550 147.485 81.740 148.355 ;
        RECT 79.625 147.195 79.795 147.365 ;
        RECT 79.125 146.815 79.455 147.195 ;
        RECT 79.625 147.025 80.920 147.195 ;
        RECT 81.090 147.150 81.280 147.465 ;
        RECT 81.540 146.815 81.740 147.315 ;
        RECT 81.910 146.985 82.240 148.565 ;
        RECT 82.415 148.605 82.930 149.015 ;
        RECT 83.165 148.605 83.335 149.365 ;
        RECT 83.505 149.025 85.535 149.195 ;
        RECT 82.415 147.795 82.755 148.605 ;
        RECT 83.505 148.360 83.675 149.025 ;
        RECT 84.070 148.685 85.195 148.855 ;
        RECT 82.925 148.170 83.675 148.360 ;
        RECT 83.845 148.345 84.855 148.515 ;
        RECT 82.415 147.625 83.645 147.795 ;
        RECT 82.690 147.020 82.935 147.625 ;
        RECT 83.155 146.815 83.665 147.350 ;
        RECT 83.845 146.985 84.035 148.345 ;
        RECT 84.205 147.325 84.480 148.145 ;
        RECT 84.685 147.545 84.855 148.345 ;
        RECT 85.025 147.555 85.195 148.685 ;
        RECT 85.365 148.055 85.535 149.025 ;
        RECT 85.705 148.225 85.875 149.365 ;
        RECT 86.045 148.225 86.380 149.195 ;
        RECT 85.365 147.725 85.560 148.055 ;
        RECT 85.785 147.725 86.040 148.055 ;
        RECT 85.785 147.555 85.955 147.725 ;
        RECT 86.210 147.555 86.380 148.225 ;
        RECT 87.480 148.215 87.740 149.365 ;
        RECT 87.915 148.290 88.170 149.195 ;
        RECT 88.340 148.605 88.670 149.365 ;
        RECT 88.885 148.435 89.055 149.195 ;
        RECT 85.025 147.385 85.955 147.555 ;
        RECT 85.025 147.350 85.200 147.385 ;
        RECT 84.205 147.155 84.485 147.325 ;
        RECT 84.205 146.985 84.480 147.155 ;
        RECT 84.670 146.985 85.200 147.350 ;
        RECT 85.625 146.815 85.955 147.215 ;
        RECT 86.125 146.985 86.380 147.555 ;
        RECT 87.480 146.815 87.740 147.655 ;
        RECT 87.915 147.560 88.085 148.290 ;
        RECT 88.340 148.265 89.055 148.435 ;
        RECT 89.775 148.565 90.215 149.195 ;
        RECT 88.340 148.055 88.510 148.265 ;
        RECT 88.255 147.725 88.510 148.055 ;
        RECT 87.915 146.985 88.170 147.560 ;
        RECT 88.340 147.535 88.510 147.725 ;
        RECT 88.790 147.715 89.145 148.085 ;
        RECT 89.775 147.555 90.085 148.565 ;
        RECT 90.390 148.515 90.705 149.365 ;
        RECT 90.875 149.025 92.305 149.195 ;
        RECT 90.875 148.345 91.045 149.025 ;
        RECT 90.255 148.175 91.045 148.345 ;
        RECT 90.255 147.725 90.425 148.175 ;
        RECT 91.215 148.055 91.415 148.855 ;
        RECT 90.595 147.725 90.985 148.005 ;
        RECT 91.170 147.725 91.415 148.055 ;
        RECT 91.615 147.725 91.865 148.855 ;
        RECT 92.055 148.395 92.305 149.025 ;
        RECT 92.485 148.565 92.815 149.365 ;
        RECT 92.055 148.225 92.825 148.395 ;
        RECT 92.080 147.725 92.485 148.055 ;
        RECT 92.655 147.555 92.825 148.225 ;
        RECT 92.995 148.200 93.285 149.365 ;
        RECT 93.460 148.695 93.715 149.195 ;
        RECT 93.885 148.865 94.215 149.365 ;
        RECT 93.460 148.525 94.210 148.695 ;
        RECT 93.460 147.705 93.810 148.355 ;
        RECT 88.340 147.365 89.055 147.535 ;
        RECT 88.340 146.815 88.670 147.195 ;
        RECT 88.885 146.985 89.055 147.365 ;
        RECT 89.775 146.995 90.215 147.555 ;
        RECT 90.385 146.815 90.835 147.555 ;
        RECT 91.005 147.385 92.165 147.555 ;
        RECT 91.005 146.985 91.175 147.385 ;
        RECT 91.345 146.815 91.765 147.215 ;
        RECT 91.935 146.985 92.165 147.385 ;
        RECT 92.335 146.985 92.825 147.555 ;
        RECT 92.995 146.815 93.285 147.540 ;
        RECT 93.980 147.535 94.210 148.525 ;
        RECT 93.460 147.365 94.210 147.535 ;
        RECT 93.460 147.075 93.715 147.365 ;
        RECT 93.885 146.815 94.215 147.195 ;
        RECT 94.385 147.075 94.555 149.195 ;
        RECT 94.725 148.395 95.050 149.180 ;
        RECT 95.220 148.905 95.470 149.365 ;
        RECT 95.640 148.865 95.890 149.195 ;
        RECT 96.105 148.865 96.785 149.195 ;
        RECT 95.640 148.735 95.810 148.865 ;
        RECT 95.415 148.565 95.810 148.735 ;
        RECT 94.785 147.345 95.245 148.395 ;
        RECT 95.415 147.205 95.585 148.565 ;
        RECT 95.980 148.305 96.445 148.695 ;
        RECT 95.755 147.495 96.105 148.115 ;
        RECT 96.275 147.715 96.445 148.305 ;
        RECT 96.615 148.085 96.785 148.865 ;
        RECT 96.955 148.765 97.125 149.105 ;
        RECT 97.360 148.935 97.690 149.365 ;
        RECT 97.860 148.765 98.030 149.105 ;
        RECT 98.325 148.905 98.695 149.365 ;
        RECT 96.955 148.595 98.030 148.765 ;
        RECT 98.865 148.735 99.035 149.195 ;
        RECT 99.270 148.855 100.140 149.195 ;
        RECT 100.310 148.905 100.560 149.365 ;
        RECT 98.475 148.565 99.035 148.735 ;
        RECT 98.475 148.425 98.645 148.565 ;
        RECT 97.145 148.255 98.645 148.425 ;
        RECT 99.340 148.395 99.800 148.685 ;
        RECT 96.615 147.915 98.305 148.085 ;
        RECT 96.275 147.495 96.630 147.715 ;
        RECT 96.800 147.205 96.970 147.915 ;
        RECT 97.175 147.495 97.965 147.745 ;
        RECT 98.135 147.735 98.305 147.915 ;
        RECT 98.475 147.565 98.645 148.255 ;
        RECT 94.915 146.815 95.245 147.175 ;
        RECT 95.415 147.035 95.910 147.205 ;
        RECT 96.115 147.035 96.970 147.205 ;
        RECT 97.845 146.815 98.175 147.275 ;
        RECT 98.385 147.175 98.645 147.565 ;
        RECT 98.835 148.385 99.800 148.395 ;
        RECT 99.970 148.475 100.140 148.855 ;
        RECT 100.730 148.815 100.900 149.105 ;
        RECT 101.080 148.985 101.410 149.365 ;
        RECT 100.730 148.645 101.530 148.815 ;
        RECT 98.835 148.225 99.510 148.385 ;
        RECT 99.970 148.305 101.190 148.475 ;
        RECT 98.835 147.435 99.045 148.225 ;
        RECT 99.970 148.215 100.140 148.305 ;
        RECT 99.215 147.435 99.565 148.055 ;
        RECT 99.735 148.045 100.140 148.215 ;
        RECT 99.735 147.265 99.905 148.045 ;
        RECT 100.075 147.595 100.295 147.875 ;
        RECT 100.475 147.765 101.015 148.135 ;
        RECT 101.360 148.055 101.530 148.645 ;
        RECT 101.750 148.225 102.055 149.365 ;
        RECT 102.225 148.175 102.480 149.055 ;
        RECT 102.655 148.275 104.325 149.365 ;
        RECT 104.740 148.610 105.070 149.365 ;
        RECT 105.240 148.815 105.430 149.195 ;
        RECT 105.600 148.985 105.930 149.365 ;
        RECT 106.100 148.815 106.310 149.195 ;
        RECT 106.480 148.925 106.760 149.365 ;
        RECT 106.930 149.005 108.910 149.195 ;
        RECT 105.240 148.755 106.310 148.815 ;
        RECT 108.720 148.815 108.910 149.005 ;
        RECT 109.080 148.985 109.410 149.365 ;
        RECT 109.580 148.815 109.815 149.195 ;
        RECT 105.240 148.585 108.550 148.755 ;
        RECT 108.720 148.645 109.815 148.815 ;
        RECT 105.240 148.430 106.455 148.585 ;
        RECT 109.985 148.550 110.270 149.365 ;
        RECT 101.360 148.025 102.100 148.055 ;
        RECT 100.075 147.425 100.605 147.595 ;
        RECT 98.385 147.005 98.735 147.175 ;
        RECT 98.955 146.985 99.905 147.265 ;
        RECT 100.075 146.815 100.265 147.255 ;
        RECT 100.435 147.195 100.605 147.425 ;
        RECT 100.775 147.365 101.015 147.765 ;
        RECT 101.185 147.725 102.100 148.025 ;
        RECT 101.185 147.550 101.510 147.725 ;
        RECT 101.185 147.195 101.505 147.550 ;
        RECT 102.270 147.525 102.480 148.175 ;
        RECT 100.435 147.025 101.505 147.195 ;
        RECT 101.750 146.815 102.055 147.275 ;
        RECT 102.225 146.995 102.480 147.525 ;
        RECT 102.655 147.585 103.405 148.105 ;
        RECT 103.575 147.755 104.325 148.275 ;
        RECT 104.555 148.175 106.455 148.430 ;
        RECT 106.695 148.245 109.815 148.415 ;
        RECT 102.655 146.815 104.325 147.585 ;
        RECT 104.555 147.575 104.965 148.175 ;
        RECT 105.135 147.745 106.485 148.005 ;
        RECT 106.695 147.720 106.945 148.245 ;
        RECT 107.115 147.800 108.405 148.075 ;
        RECT 108.915 148.050 109.815 148.245 ;
        RECT 110.945 148.395 111.275 149.180 ;
        RECT 110.945 148.225 111.625 148.395 ;
        RECT 111.805 148.225 112.135 149.365 ;
        RECT 112.320 148.735 112.655 149.195 ;
        RECT 112.825 148.905 113.045 149.365 ;
        RECT 113.575 148.985 114.885 149.155 ;
        RECT 114.715 148.735 114.885 148.985 ;
        RECT 115.055 148.905 115.345 149.365 ;
        RECT 112.320 148.565 114.545 148.735 ;
        RECT 114.715 148.565 115.375 148.735 ;
        RECT 108.915 147.745 110.265 148.050 ;
        RECT 110.935 147.805 111.285 148.055 ;
        RECT 111.455 147.625 111.625 148.225 ;
        RECT 111.795 147.805 112.145 148.055 ;
        RECT 104.555 147.345 106.360 147.575 ;
        RECT 106.530 147.345 110.270 147.550 ;
        RECT 106.530 147.175 106.760 147.345 ;
        RECT 104.740 146.985 106.760 147.175 ;
        RECT 106.930 146.815 107.260 147.175 ;
        RECT 107.790 146.815 108.120 147.175 ;
        RECT 108.650 146.815 108.980 147.175 ;
        RECT 109.510 146.815 109.840 147.175 ;
        RECT 110.955 146.815 111.195 147.625 ;
        RECT 111.365 146.985 111.695 147.625 ;
        RECT 111.865 146.815 112.135 147.625 ;
        RECT 112.320 146.985 112.650 148.565 ;
        RECT 114.375 148.395 114.545 148.565 ;
        RECT 112.820 147.485 113.010 148.355 ;
        RECT 113.280 148.045 114.095 148.355 ;
        RECT 114.375 148.225 115.035 148.395 ;
        RECT 113.925 148.010 114.095 148.045 ;
        RECT 113.280 147.465 113.745 147.755 ;
        RECT 113.925 147.495 114.555 148.010 ;
        RECT 114.865 147.725 115.035 148.225 ;
        RECT 115.205 148.055 115.375 148.565 ;
        RECT 115.545 148.325 115.855 149.195 ;
        RECT 115.205 147.725 115.515 148.055 ;
        RECT 115.205 147.535 115.375 147.725 ;
        RECT 112.820 146.815 113.020 147.315 ;
        RECT 113.280 147.150 113.470 147.465 ;
        RECT 114.765 147.365 115.375 147.535 ;
        RECT 115.685 147.480 115.855 148.325 ;
        RECT 116.025 148.225 116.280 149.365 ;
        RECT 117.375 148.225 117.635 149.365 ;
        RECT 117.805 148.215 118.135 149.195 ;
        RECT 118.305 148.225 118.585 149.365 ;
        RECT 117.395 147.805 117.730 148.055 ;
        RECT 117.900 147.615 118.070 148.215 ;
        RECT 118.755 148.200 119.045 149.365 ;
        RECT 119.715 148.415 120.005 149.185 ;
        RECT 120.575 148.825 120.835 149.185 ;
        RECT 121.005 148.995 121.335 149.365 ;
        RECT 121.505 148.825 121.765 149.185 ;
        RECT 120.575 148.595 121.765 148.825 ;
        RECT 121.955 148.645 122.285 149.365 ;
        RECT 122.455 148.415 122.720 149.185 ;
        RECT 119.715 148.235 122.210 148.415 ;
        RECT 118.240 147.785 118.575 148.055 ;
        RECT 119.685 147.725 119.955 148.055 ;
        RECT 120.135 147.725 120.570 148.055 ;
        RECT 120.750 147.725 121.325 148.055 ;
        RECT 121.505 147.725 121.785 148.055 ;
        RECT 114.765 147.195 114.935 147.365 ;
        RECT 113.640 147.025 114.935 147.195 ;
        RECT 115.105 146.815 115.435 147.195 ;
        RECT 115.605 146.985 115.855 147.480 ;
        RECT 116.025 146.815 116.280 147.615 ;
        RECT 117.375 146.985 118.070 147.615 ;
        RECT 118.275 146.815 118.585 147.615 ;
        RECT 121.985 147.545 122.210 148.235 ;
        RECT 118.755 146.815 119.045 147.540 ;
        RECT 119.725 147.355 122.210 147.545 ;
        RECT 119.725 146.995 119.950 147.355 ;
        RECT 120.130 146.815 120.460 147.185 ;
        RECT 120.640 146.995 120.895 147.355 ;
        RECT 121.460 146.815 122.205 147.185 ;
        RECT 122.385 146.995 122.720 148.415 ;
        RECT 123.100 148.395 123.430 149.195 ;
        RECT 123.600 148.565 123.930 149.365 ;
        RECT 124.230 148.395 124.560 149.195 ;
        RECT 125.205 148.565 125.455 149.365 ;
        RECT 123.100 148.225 125.535 148.395 ;
        RECT 125.725 148.225 125.895 149.365 ;
        RECT 126.065 148.225 126.405 149.195 ;
        RECT 122.895 147.805 123.245 148.055 ;
        RECT 123.430 147.595 123.600 148.225 ;
        RECT 123.770 147.805 124.100 148.005 ;
        RECT 124.270 147.805 124.600 148.005 ;
        RECT 124.770 147.805 125.190 148.005 ;
        RECT 125.365 147.975 125.535 148.225 ;
        RECT 125.365 147.805 126.060 147.975 ;
        RECT 123.100 146.985 123.600 147.595 ;
        RECT 124.230 147.465 125.455 147.635 ;
        RECT 126.230 147.615 126.405 148.225 ;
        RECT 126.575 148.605 127.090 149.015 ;
        RECT 127.325 148.605 127.495 149.365 ;
        RECT 127.665 149.025 129.695 149.195 ;
        RECT 126.575 147.795 126.915 148.605 ;
        RECT 127.665 148.360 127.835 149.025 ;
        RECT 128.230 148.685 129.355 148.855 ;
        RECT 127.085 148.170 127.835 148.360 ;
        RECT 128.005 148.345 129.015 148.515 ;
        RECT 126.575 147.625 127.805 147.795 ;
        RECT 124.230 146.985 124.560 147.465 ;
        RECT 124.730 146.815 124.955 147.275 ;
        RECT 125.125 146.985 125.455 147.465 ;
        RECT 125.645 146.815 125.895 147.615 ;
        RECT 126.065 146.985 126.405 147.615 ;
        RECT 126.850 147.020 127.095 147.625 ;
        RECT 127.315 146.815 127.825 147.350 ;
        RECT 128.005 146.985 128.195 148.345 ;
        RECT 128.365 147.325 128.640 148.145 ;
        RECT 128.845 147.545 129.015 148.345 ;
        RECT 129.185 147.555 129.355 148.685 ;
        RECT 129.525 148.055 129.695 149.025 ;
        RECT 129.865 148.225 130.035 149.365 ;
        RECT 130.205 148.225 130.540 149.195 ;
        RECT 131.645 148.395 131.975 149.195 ;
        RECT 132.145 148.565 132.375 149.365 ;
        RECT 132.545 148.395 132.875 149.195 ;
        RECT 131.645 148.225 132.875 148.395 ;
        RECT 133.045 148.225 133.300 149.365 ;
        RECT 133.940 148.695 134.195 149.195 ;
        RECT 134.365 148.865 134.695 149.365 ;
        RECT 133.940 148.525 134.690 148.695 ;
        RECT 129.525 147.725 129.720 148.055 ;
        RECT 129.945 147.725 130.200 148.055 ;
        RECT 129.945 147.555 130.115 147.725 ;
        RECT 130.370 147.555 130.540 148.225 ;
        RECT 131.635 147.725 131.945 148.055 ;
        RECT 129.185 147.385 130.115 147.555 ;
        RECT 129.185 147.350 129.360 147.385 ;
        RECT 128.365 147.155 128.645 147.325 ;
        RECT 128.365 146.985 128.640 147.155 ;
        RECT 128.830 146.985 129.360 147.350 ;
        RECT 129.785 146.815 130.115 147.215 ;
        RECT 130.285 146.985 130.540 147.555 ;
        RECT 131.645 147.325 131.975 147.555 ;
        RECT 132.150 147.495 132.525 148.055 ;
        RECT 132.695 147.325 132.875 148.225 ;
        RECT 133.060 147.475 133.280 148.055 ;
        RECT 133.940 147.705 134.290 148.355 ;
        RECT 134.460 147.535 134.690 148.525 ;
        RECT 131.645 146.985 132.875 147.325 ;
        RECT 133.940 147.365 134.690 147.535 ;
        RECT 133.045 146.815 133.300 147.305 ;
        RECT 133.940 147.075 134.195 147.365 ;
        RECT 134.365 146.815 134.695 147.195 ;
        RECT 134.865 147.075 135.035 149.195 ;
        RECT 135.205 148.395 135.530 149.180 ;
        RECT 135.700 148.905 135.950 149.365 ;
        RECT 136.120 148.865 136.370 149.195 ;
        RECT 136.585 148.865 137.265 149.195 ;
        RECT 136.120 148.735 136.290 148.865 ;
        RECT 135.895 148.565 136.290 148.735 ;
        RECT 135.265 147.345 135.725 148.395 ;
        RECT 135.895 147.205 136.065 148.565 ;
        RECT 136.460 148.305 136.925 148.695 ;
        RECT 136.235 147.495 136.585 148.115 ;
        RECT 136.755 147.715 136.925 148.305 ;
        RECT 137.095 148.085 137.265 148.865 ;
        RECT 137.435 148.765 137.605 149.105 ;
        RECT 137.840 148.935 138.170 149.365 ;
        RECT 138.340 148.765 138.510 149.105 ;
        RECT 138.805 148.905 139.175 149.365 ;
        RECT 137.435 148.595 138.510 148.765 ;
        RECT 139.345 148.735 139.515 149.195 ;
        RECT 139.750 148.855 140.620 149.195 ;
        RECT 140.790 148.905 141.040 149.365 ;
        RECT 138.955 148.565 139.515 148.735 ;
        RECT 138.955 148.425 139.125 148.565 ;
        RECT 137.625 148.255 139.125 148.425 ;
        RECT 139.820 148.395 140.280 148.685 ;
        RECT 137.095 147.915 138.785 148.085 ;
        RECT 136.755 147.495 137.110 147.715 ;
        RECT 137.280 147.205 137.450 147.915 ;
        RECT 137.655 147.495 138.445 147.745 ;
        RECT 138.615 147.735 138.785 147.915 ;
        RECT 138.955 147.565 139.125 148.255 ;
        RECT 135.395 146.815 135.725 147.175 ;
        RECT 135.895 147.035 136.390 147.205 ;
        RECT 136.595 147.035 137.450 147.205 ;
        RECT 138.325 146.815 138.655 147.275 ;
        RECT 138.865 147.175 139.125 147.565 ;
        RECT 139.315 148.385 140.280 148.395 ;
        RECT 140.450 148.475 140.620 148.855 ;
        RECT 141.210 148.815 141.380 149.105 ;
        RECT 141.560 148.985 141.890 149.365 ;
        RECT 141.210 148.645 142.010 148.815 ;
        RECT 139.315 148.225 139.990 148.385 ;
        RECT 140.450 148.305 141.670 148.475 ;
        RECT 139.315 147.435 139.525 148.225 ;
        RECT 140.450 148.215 140.620 148.305 ;
        RECT 139.695 147.435 140.045 148.055 ;
        RECT 140.215 148.045 140.620 148.215 ;
        RECT 140.215 147.265 140.385 148.045 ;
        RECT 140.555 147.595 140.775 147.875 ;
        RECT 140.955 147.765 141.495 148.135 ;
        RECT 141.840 148.025 142.010 148.645 ;
        RECT 142.185 148.305 142.355 149.365 ;
        RECT 142.565 148.355 142.855 149.195 ;
        RECT 143.025 148.525 143.195 149.365 ;
        RECT 143.405 148.355 143.655 149.195 ;
        RECT 143.865 148.525 144.035 149.365 ;
        RECT 142.565 148.185 144.290 148.355 ;
        RECT 144.515 148.200 144.805 149.365 ;
        RECT 144.975 148.930 150.320 149.365 ;
        RECT 150.495 148.930 155.840 149.365 ;
        RECT 140.555 147.425 141.085 147.595 ;
        RECT 138.865 147.005 139.215 147.175 ;
        RECT 139.435 146.985 140.385 147.265 ;
        RECT 140.555 146.815 140.745 147.255 ;
        RECT 140.915 147.195 141.085 147.425 ;
        RECT 141.255 147.365 141.495 147.765 ;
        RECT 141.665 148.015 142.010 148.025 ;
        RECT 141.665 147.805 143.695 148.015 ;
        RECT 141.665 147.550 141.990 147.805 ;
        RECT 143.880 147.635 144.290 148.185 ;
        RECT 141.665 147.195 141.985 147.550 ;
        RECT 140.915 147.025 141.985 147.195 ;
        RECT 142.185 146.815 142.355 147.625 ;
        RECT 142.525 147.465 144.290 147.635 ;
        RECT 142.525 146.985 142.855 147.465 ;
        RECT 143.025 146.815 143.195 147.285 ;
        RECT 143.365 146.985 143.695 147.465 ;
        RECT 143.865 146.815 144.035 147.285 ;
        RECT 144.515 146.815 144.805 147.540 ;
        RECT 146.560 147.360 146.900 148.190 ;
        RECT 148.380 147.680 148.730 148.930 ;
        RECT 152.080 147.360 152.420 148.190 ;
        RECT 153.900 147.680 154.250 148.930 ;
        RECT 156.935 148.275 158.145 149.365 ;
        RECT 156.935 147.735 157.455 148.275 ;
        RECT 157.625 147.565 158.145 148.105 ;
        RECT 144.975 146.815 150.320 147.360 ;
        RECT 150.495 146.815 155.840 147.360 ;
        RECT 156.935 146.815 158.145 147.565 ;
        RECT 2.750 146.645 158.230 146.815 ;
        RECT 2.835 145.895 4.045 146.645 ;
        RECT 2.835 145.355 3.355 145.895 ;
        RECT 3.525 145.185 4.045 145.725 ;
        RECT 2.835 144.095 4.045 145.185 ;
        RECT 5.140 145.045 5.475 146.465 ;
        RECT 5.655 146.275 6.400 146.645 ;
        RECT 6.965 146.105 7.220 146.465 ;
        RECT 7.400 146.275 7.730 146.645 ;
        RECT 7.910 146.105 8.135 146.465 ;
        RECT 5.650 145.915 8.135 146.105 ;
        RECT 5.650 145.225 5.875 145.915 ;
        RECT 8.360 145.905 8.615 146.475 ;
        RECT 8.785 146.245 9.115 146.645 ;
        RECT 9.540 146.110 10.070 146.475 ;
        RECT 9.540 146.075 9.715 146.110 ;
        RECT 8.785 145.905 9.715 146.075 ;
        RECT 10.260 145.965 10.535 146.475 ;
        RECT 6.075 145.405 6.355 145.735 ;
        RECT 6.535 145.405 7.110 145.735 ;
        RECT 7.290 145.405 7.725 145.735 ;
        RECT 7.905 145.405 8.175 145.735 ;
        RECT 8.360 145.235 8.530 145.905 ;
        RECT 8.785 145.735 8.955 145.905 ;
        RECT 8.700 145.405 8.955 145.735 ;
        RECT 9.180 145.405 9.375 145.735 ;
        RECT 5.650 145.045 8.145 145.225 ;
        RECT 5.140 144.275 5.405 145.045 ;
        RECT 5.575 144.095 5.905 144.815 ;
        RECT 6.095 144.635 7.285 144.865 ;
        RECT 6.095 144.275 6.355 144.635 ;
        RECT 6.525 144.095 6.855 144.465 ;
        RECT 7.025 144.275 7.285 144.635 ;
        RECT 7.855 144.275 8.145 145.045 ;
        RECT 8.360 144.265 8.695 145.235 ;
        RECT 8.865 144.095 9.035 145.235 ;
        RECT 9.205 144.435 9.375 145.405 ;
        RECT 9.545 144.775 9.715 145.905 ;
        RECT 9.885 145.115 10.055 145.915 ;
        RECT 10.255 145.795 10.535 145.965 ;
        RECT 10.260 145.315 10.535 145.795 ;
        RECT 10.705 145.115 10.895 146.475 ;
        RECT 11.075 146.110 11.585 146.645 ;
        RECT 11.805 145.835 12.050 146.440 ;
        RECT 12.500 145.905 12.755 146.475 ;
        RECT 12.925 146.245 13.255 146.645 ;
        RECT 13.680 146.110 14.210 146.475 ;
        RECT 13.680 146.075 13.855 146.110 ;
        RECT 12.925 145.905 13.855 146.075 ;
        RECT 11.095 145.665 12.325 145.835 ;
        RECT 9.885 144.945 10.895 145.115 ;
        RECT 11.065 145.100 11.815 145.290 ;
        RECT 9.545 144.605 10.670 144.775 ;
        RECT 11.065 144.435 11.235 145.100 ;
        RECT 11.985 144.855 12.325 145.665 ;
        RECT 9.205 144.265 11.235 144.435 ;
        RECT 11.405 144.095 11.575 144.855 ;
        RECT 11.810 144.445 12.325 144.855 ;
        RECT 12.500 145.235 12.670 145.905 ;
        RECT 12.925 145.735 13.095 145.905 ;
        RECT 12.840 145.405 13.095 145.735 ;
        RECT 13.320 145.405 13.515 145.735 ;
        RECT 12.500 144.265 12.835 145.235 ;
        RECT 13.005 144.095 13.175 145.235 ;
        RECT 13.345 144.435 13.515 145.405 ;
        RECT 13.685 144.775 13.855 145.905 ;
        RECT 14.025 145.115 14.195 145.915 ;
        RECT 14.400 145.625 14.675 146.475 ;
        RECT 14.395 145.455 14.675 145.625 ;
        RECT 14.400 145.315 14.675 145.455 ;
        RECT 14.845 145.115 15.035 146.475 ;
        RECT 15.215 146.110 15.725 146.645 ;
        RECT 15.945 145.835 16.190 146.440 ;
        RECT 17.100 145.880 17.555 146.645 ;
        RECT 17.830 146.265 19.130 146.475 ;
        RECT 19.385 146.285 19.715 146.645 ;
        RECT 18.960 146.115 19.130 146.265 ;
        RECT 19.885 146.145 20.145 146.475 ;
        RECT 15.235 145.665 16.465 145.835 ;
        RECT 14.025 144.945 15.035 145.115 ;
        RECT 15.205 145.100 15.955 145.290 ;
        RECT 13.685 144.605 14.810 144.775 ;
        RECT 15.205 144.435 15.375 145.100 ;
        RECT 16.125 144.855 16.465 145.665 ;
        RECT 18.030 145.655 18.250 146.055 ;
        RECT 17.095 145.455 17.585 145.655 ;
        RECT 17.775 145.445 18.250 145.655 ;
        RECT 18.495 145.655 18.705 146.055 ;
        RECT 18.960 145.990 19.715 146.115 ;
        RECT 18.960 145.945 19.805 145.990 ;
        RECT 19.535 145.825 19.805 145.945 ;
        RECT 18.495 145.445 18.825 145.655 ;
        RECT 18.995 145.385 19.405 145.690 ;
        RECT 13.345 144.265 15.375 144.435 ;
        RECT 15.545 144.095 15.715 144.855 ;
        RECT 15.950 144.445 16.465 144.855 ;
        RECT 17.100 145.215 18.275 145.275 ;
        RECT 19.635 145.250 19.805 145.825 ;
        RECT 19.605 145.215 19.805 145.250 ;
        RECT 17.100 145.105 19.805 145.215 ;
        RECT 17.100 144.485 17.355 145.105 ;
        RECT 17.945 145.045 19.745 145.105 ;
        RECT 17.945 145.015 18.275 145.045 ;
        RECT 19.975 144.945 20.145 146.145 ;
        RECT 20.365 146.105 20.590 146.465 ;
        RECT 20.770 146.275 21.100 146.645 ;
        RECT 21.280 146.105 21.535 146.465 ;
        RECT 22.100 146.275 22.845 146.645 ;
        RECT 20.365 145.915 22.850 146.105 ;
        RECT 20.325 145.405 20.595 145.735 ;
        RECT 20.775 145.405 21.210 145.735 ;
        RECT 21.390 145.405 21.965 145.735 ;
        RECT 22.145 145.405 22.425 145.735 ;
        RECT 22.625 145.225 22.850 145.915 ;
        RECT 17.605 144.845 17.790 144.935 ;
        RECT 18.380 144.845 19.215 144.855 ;
        RECT 17.605 144.645 19.215 144.845 ;
        RECT 17.605 144.605 17.835 144.645 ;
        RECT 17.100 144.265 17.435 144.485 ;
        RECT 18.440 144.095 18.795 144.475 ;
        RECT 18.965 144.265 19.215 144.645 ;
        RECT 19.465 144.095 19.715 144.875 ;
        RECT 19.885 144.265 20.145 144.945 ;
        RECT 20.355 145.045 22.850 145.225 ;
        RECT 23.025 145.045 23.360 146.465 ;
        RECT 23.625 146.095 23.795 146.475 ;
        RECT 23.975 146.265 24.305 146.645 ;
        RECT 23.625 145.925 24.290 146.095 ;
        RECT 24.485 145.970 24.745 146.475 ;
        RECT 23.555 145.375 23.885 145.745 ;
        RECT 24.120 145.670 24.290 145.925 ;
        RECT 24.120 145.340 24.405 145.670 ;
        RECT 24.120 145.195 24.290 145.340 ;
        RECT 20.355 144.275 20.645 145.045 ;
        RECT 21.215 144.635 22.405 144.865 ;
        RECT 21.215 144.275 21.475 144.635 ;
        RECT 21.645 144.095 21.975 144.465 ;
        RECT 22.145 144.275 22.405 144.635 ;
        RECT 22.595 144.095 22.925 144.815 ;
        RECT 23.095 144.275 23.360 145.045 ;
        RECT 23.625 145.025 24.290 145.195 ;
        RECT 24.575 145.170 24.745 145.970 ;
        RECT 25.015 145.845 25.185 146.645 ;
        RECT 23.625 144.265 23.795 145.025 ;
        RECT 23.975 144.095 24.305 144.855 ;
        RECT 24.475 144.265 24.745 145.170 ;
        RECT 24.945 144.095 25.195 145.285 ;
        RECT 25.420 144.265 25.635 146.365 ;
        RECT 25.855 146.185 26.035 146.645 ;
        RECT 26.295 146.255 27.560 146.435 ;
        RECT 26.680 146.015 27.045 146.085 ;
        RECT 25.805 145.835 27.045 146.015 ;
        RECT 27.220 146.035 27.560 146.255 ;
        RECT 27.745 146.205 27.915 146.645 ;
        RECT 28.085 146.035 28.420 146.450 ;
        RECT 27.220 145.905 28.420 146.035 ;
        RECT 28.595 145.920 28.885 146.645 ;
        RECT 27.390 145.865 28.420 145.905 ;
        RECT 25.805 145.235 26.085 145.835 ;
        RECT 30.035 145.825 30.245 146.645 ;
        RECT 30.415 145.845 30.745 146.475 ;
        RECT 26.265 145.405 26.620 145.655 ;
        RECT 26.790 145.405 27.255 145.655 ;
        RECT 27.425 145.405 27.755 145.655 ;
        RECT 27.925 145.455 28.420 145.655 ;
        RECT 27.575 145.285 27.755 145.405 ;
        RECT 25.805 145.025 27.405 145.235 ;
        RECT 27.575 145.115 27.930 145.285 ;
        RECT 28.100 145.115 28.420 145.455 ;
        RECT 25.825 144.095 26.625 144.855 ;
        RECT 27.020 144.265 27.405 145.025 ;
        RECT 27.730 144.325 27.930 145.115 ;
        RECT 28.100 144.095 28.420 144.935 ;
        RECT 28.595 144.095 28.885 145.260 ;
        RECT 30.415 145.245 30.665 145.845 ;
        RECT 30.915 145.825 31.145 146.645 ;
        RECT 31.355 145.905 31.740 146.475 ;
        RECT 31.910 146.185 32.235 146.645 ;
        RECT 32.755 146.015 33.035 146.475 ;
        RECT 30.835 145.405 31.165 145.655 ;
        RECT 30.035 144.095 30.245 145.235 ;
        RECT 30.415 144.265 30.745 145.245 ;
        RECT 31.355 145.235 31.635 145.905 ;
        RECT 31.910 145.845 33.035 146.015 ;
        RECT 31.910 145.735 32.360 145.845 ;
        RECT 31.805 145.405 32.360 145.735 ;
        RECT 33.225 145.675 33.625 146.475 ;
        RECT 34.025 146.185 34.295 146.645 ;
        RECT 34.465 146.015 34.750 146.475 ;
        RECT 30.915 144.095 31.145 145.235 ;
        RECT 31.355 144.265 31.740 145.235 ;
        RECT 31.910 144.945 32.360 145.405 ;
        RECT 32.530 145.115 33.625 145.675 ;
        RECT 31.910 144.725 33.035 144.945 ;
        RECT 31.910 144.095 32.235 144.555 ;
        RECT 32.755 144.265 33.035 144.725 ;
        RECT 33.225 144.265 33.625 145.115 ;
        RECT 33.795 145.845 34.750 146.015 ;
        RECT 35.150 146.015 35.435 146.475 ;
        RECT 35.605 146.185 35.875 146.645 ;
        RECT 35.150 145.845 36.105 146.015 ;
        RECT 33.795 144.945 34.005 145.845 ;
        RECT 34.175 145.115 34.865 145.675 ;
        RECT 35.035 145.115 35.725 145.675 ;
        RECT 35.895 144.945 36.105 145.845 ;
        RECT 33.795 144.725 34.750 144.945 ;
        RECT 34.025 144.095 34.295 144.555 ;
        RECT 34.465 144.265 34.750 144.725 ;
        RECT 35.150 144.725 36.105 144.945 ;
        RECT 36.275 145.675 36.675 146.475 ;
        RECT 36.865 146.015 37.145 146.475 ;
        RECT 37.665 146.185 37.990 146.645 ;
        RECT 36.865 145.845 37.990 146.015 ;
        RECT 38.160 145.905 38.545 146.475 ;
        RECT 38.720 146.095 38.975 146.385 ;
        RECT 39.145 146.265 39.475 146.645 ;
        RECT 38.720 145.925 39.470 146.095 ;
        RECT 37.540 145.735 37.990 145.845 ;
        RECT 36.275 145.115 37.370 145.675 ;
        RECT 37.540 145.405 38.095 145.735 ;
        RECT 35.150 144.265 35.435 144.725 ;
        RECT 35.605 144.095 35.875 144.555 ;
        RECT 36.275 144.265 36.675 145.115 ;
        RECT 37.540 144.945 37.990 145.405 ;
        RECT 38.265 145.235 38.545 145.905 ;
        RECT 36.865 144.725 37.990 144.945 ;
        RECT 36.865 144.265 37.145 144.725 ;
        RECT 37.665 144.095 37.990 144.555 ;
        RECT 38.160 144.265 38.545 145.235 ;
        RECT 38.720 145.105 39.070 145.755 ;
        RECT 39.240 144.935 39.470 145.925 ;
        RECT 38.720 144.765 39.470 144.935 ;
        RECT 38.720 144.265 38.975 144.765 ;
        RECT 39.145 144.095 39.475 144.595 ;
        RECT 39.645 144.265 39.815 146.385 ;
        RECT 40.175 146.285 40.505 146.645 ;
        RECT 40.675 146.255 41.170 146.425 ;
        RECT 41.375 146.255 42.230 146.425 ;
        RECT 40.045 145.065 40.505 146.115 ;
        RECT 39.985 144.280 40.310 145.065 ;
        RECT 40.675 144.895 40.845 146.255 ;
        RECT 41.015 145.345 41.365 145.965 ;
        RECT 41.535 145.745 41.890 145.965 ;
        RECT 41.535 145.155 41.705 145.745 ;
        RECT 42.060 145.545 42.230 146.255 ;
        RECT 43.105 146.185 43.435 146.645 ;
        RECT 43.645 146.285 43.995 146.455 ;
        RECT 42.435 145.715 43.225 145.965 ;
        RECT 43.645 145.895 43.905 146.285 ;
        RECT 44.215 146.195 45.165 146.475 ;
        RECT 45.335 146.205 45.525 146.645 ;
        RECT 45.695 146.265 46.765 146.435 ;
        RECT 43.395 145.545 43.565 145.725 ;
        RECT 40.675 144.725 41.070 144.895 ;
        RECT 41.240 144.765 41.705 145.155 ;
        RECT 41.875 145.375 43.565 145.545 ;
        RECT 40.900 144.595 41.070 144.725 ;
        RECT 41.875 144.595 42.045 145.375 ;
        RECT 43.735 145.205 43.905 145.895 ;
        RECT 42.405 145.035 43.905 145.205 ;
        RECT 44.095 145.235 44.305 146.025 ;
        RECT 44.475 145.405 44.825 146.025 ;
        RECT 44.995 145.415 45.165 146.195 ;
        RECT 45.695 146.035 45.865 146.265 ;
        RECT 45.335 145.865 45.865 146.035 ;
        RECT 45.335 145.585 45.555 145.865 ;
        RECT 46.035 145.695 46.275 146.095 ;
        RECT 44.995 145.245 45.400 145.415 ;
        RECT 45.735 145.325 46.275 145.695 ;
        RECT 46.445 145.910 46.765 146.265 ;
        RECT 47.010 146.185 47.315 146.645 ;
        RECT 47.485 145.935 47.740 146.465 ;
        RECT 46.445 145.735 46.770 145.910 ;
        RECT 46.445 145.435 47.360 145.735 ;
        RECT 46.620 145.405 47.360 145.435 ;
        RECT 44.095 145.075 44.770 145.235 ;
        RECT 45.230 145.155 45.400 145.245 ;
        RECT 44.095 145.065 45.060 145.075 ;
        RECT 43.735 144.895 43.905 145.035 ;
        RECT 40.480 144.095 40.730 144.555 ;
        RECT 40.900 144.265 41.150 144.595 ;
        RECT 41.365 144.265 42.045 144.595 ;
        RECT 42.215 144.695 43.290 144.865 ;
        RECT 43.735 144.725 44.295 144.895 ;
        RECT 44.600 144.775 45.060 145.065 ;
        RECT 45.230 144.985 46.450 145.155 ;
        RECT 42.215 144.355 42.385 144.695 ;
        RECT 42.620 144.095 42.950 144.525 ;
        RECT 43.120 144.355 43.290 144.695 ;
        RECT 43.585 144.095 43.955 144.555 ;
        RECT 44.125 144.265 44.295 144.725 ;
        RECT 45.230 144.605 45.400 144.985 ;
        RECT 46.620 144.815 46.790 145.405 ;
        RECT 47.530 145.285 47.740 145.935 ;
        RECT 48.475 145.845 48.645 146.645 ;
        RECT 44.530 144.265 45.400 144.605 ;
        RECT 45.990 144.645 46.790 144.815 ;
        RECT 45.570 144.095 45.820 144.555 ;
        RECT 45.990 144.355 46.160 144.645 ;
        RECT 46.340 144.095 46.670 144.475 ;
        RECT 47.010 144.095 47.315 145.235 ;
        RECT 47.485 144.405 47.740 145.285 ;
        RECT 48.405 144.095 48.655 145.285 ;
        RECT 48.880 144.265 49.095 146.365 ;
        RECT 49.315 146.185 49.495 146.645 ;
        RECT 49.755 146.255 51.020 146.435 ;
        RECT 50.140 146.015 50.505 146.085 ;
        RECT 49.265 145.835 50.505 146.015 ;
        RECT 50.680 146.035 51.020 146.255 ;
        RECT 51.205 146.205 51.375 146.645 ;
        RECT 51.545 146.035 51.880 146.450 ;
        RECT 50.680 145.905 51.880 146.035 ;
        RECT 53.065 146.095 53.235 146.475 ;
        RECT 53.415 146.265 53.745 146.645 ;
        RECT 53.065 145.925 53.730 146.095 ;
        RECT 53.925 145.970 54.185 146.475 ;
        RECT 50.850 145.865 51.880 145.905 ;
        RECT 49.265 145.235 49.545 145.835 ;
        RECT 49.725 145.405 50.080 145.655 ;
        RECT 50.250 145.405 50.715 145.655 ;
        RECT 50.885 145.405 51.215 145.655 ;
        RECT 51.385 145.455 51.880 145.655 ;
        RECT 51.035 145.285 51.215 145.405 ;
        RECT 49.265 145.025 50.865 145.235 ;
        RECT 51.035 145.115 51.390 145.285 ;
        RECT 51.560 145.115 51.880 145.455 ;
        RECT 52.995 145.375 53.325 145.745 ;
        RECT 53.560 145.670 53.730 145.925 ;
        RECT 53.560 145.340 53.845 145.670 ;
        RECT 53.560 145.195 53.730 145.340 ;
        RECT 49.285 144.095 50.085 144.855 ;
        RECT 50.480 144.265 50.865 145.025 ;
        RECT 51.190 144.325 51.390 145.115 ;
        RECT 53.065 145.025 53.730 145.195 ;
        RECT 54.015 145.170 54.185 145.970 ;
        RECT 54.355 145.920 54.645 146.645 ;
        RECT 54.815 145.845 55.510 146.475 ;
        RECT 55.715 145.845 56.025 146.645 ;
        RECT 54.835 145.405 55.170 145.655 ;
        RECT 55.340 145.285 55.510 145.845 ;
        RECT 56.930 145.835 57.175 146.440 ;
        RECT 57.395 146.110 57.905 146.645 ;
        RECT 55.680 145.405 56.015 145.675 ;
        RECT 56.655 145.665 57.885 145.835 ;
        RECT 51.560 144.095 51.880 144.935 ;
        RECT 53.065 144.265 53.235 145.025 ;
        RECT 53.415 144.095 53.745 144.855 ;
        RECT 53.915 144.265 54.185 145.170 ;
        RECT 54.355 144.095 54.645 145.260 ;
        RECT 55.335 145.245 55.510 145.285 ;
        RECT 54.815 144.095 55.075 145.235 ;
        RECT 55.245 144.265 55.575 145.245 ;
        RECT 55.745 144.095 56.025 145.235 ;
        RECT 56.655 144.855 56.995 145.665 ;
        RECT 57.165 145.100 57.915 145.290 ;
        RECT 56.655 144.445 57.170 144.855 ;
        RECT 57.405 144.095 57.575 144.855 ;
        RECT 57.745 144.435 57.915 145.100 ;
        RECT 58.085 145.115 58.275 146.475 ;
        RECT 58.445 146.305 58.720 146.475 ;
        RECT 58.445 146.135 58.725 146.305 ;
        RECT 58.445 145.315 58.720 146.135 ;
        RECT 58.910 146.110 59.440 146.475 ;
        RECT 59.865 146.245 60.195 146.645 ;
        RECT 59.265 146.075 59.440 146.110 ;
        RECT 58.925 145.115 59.095 145.915 ;
        RECT 58.085 144.945 59.095 145.115 ;
        RECT 59.265 145.905 60.195 146.075 ;
        RECT 60.365 145.905 60.620 146.475 ;
        RECT 60.885 146.095 61.055 146.475 ;
        RECT 61.270 146.265 61.600 146.645 ;
        RECT 60.885 145.925 61.600 146.095 ;
        RECT 59.265 144.775 59.435 145.905 ;
        RECT 60.025 145.735 60.195 145.905 ;
        RECT 58.310 144.605 59.435 144.775 ;
        RECT 59.605 145.405 59.800 145.735 ;
        RECT 60.025 145.405 60.280 145.735 ;
        RECT 59.605 144.435 59.775 145.405 ;
        RECT 60.450 145.235 60.620 145.905 ;
        RECT 60.795 145.375 61.150 145.745 ;
        RECT 61.430 145.735 61.600 145.925 ;
        RECT 61.770 145.900 62.025 146.475 ;
        RECT 61.430 145.405 61.685 145.735 ;
        RECT 57.745 144.265 59.775 144.435 ;
        RECT 59.945 144.095 60.115 145.235 ;
        RECT 60.285 144.265 60.620 145.235 ;
        RECT 61.430 145.195 61.600 145.405 ;
        RECT 60.885 145.025 61.600 145.195 ;
        RECT 61.855 145.170 62.025 145.900 ;
        RECT 62.200 145.805 62.460 146.645 ;
        RECT 62.640 146.095 62.895 146.385 ;
        RECT 63.065 146.265 63.395 146.645 ;
        RECT 62.640 145.925 63.390 146.095 ;
        RECT 60.885 144.265 61.055 145.025 ;
        RECT 61.270 144.095 61.600 144.855 ;
        RECT 61.770 144.265 62.025 145.170 ;
        RECT 62.200 144.095 62.460 145.245 ;
        RECT 62.640 145.105 62.990 145.755 ;
        RECT 63.160 144.935 63.390 145.925 ;
        RECT 62.640 144.765 63.390 144.935 ;
        RECT 62.640 144.265 62.895 144.765 ;
        RECT 63.065 144.095 63.395 144.595 ;
        RECT 63.565 144.265 63.735 146.385 ;
        RECT 64.095 146.285 64.425 146.645 ;
        RECT 64.595 146.255 65.090 146.425 ;
        RECT 65.295 146.255 66.150 146.425 ;
        RECT 63.965 145.065 64.425 146.115 ;
        RECT 63.905 144.280 64.230 145.065 ;
        RECT 64.595 144.895 64.765 146.255 ;
        RECT 64.935 145.345 65.285 145.965 ;
        RECT 65.455 145.745 65.810 145.965 ;
        RECT 65.455 145.155 65.625 145.745 ;
        RECT 65.980 145.545 66.150 146.255 ;
        RECT 67.025 146.185 67.355 146.645 ;
        RECT 67.565 146.285 67.915 146.455 ;
        RECT 66.355 145.715 67.145 145.965 ;
        RECT 67.565 145.895 67.825 146.285 ;
        RECT 68.135 146.195 69.085 146.475 ;
        RECT 69.255 146.205 69.445 146.645 ;
        RECT 69.615 146.265 70.685 146.435 ;
        RECT 67.315 145.545 67.485 145.725 ;
        RECT 64.595 144.725 64.990 144.895 ;
        RECT 65.160 144.765 65.625 145.155 ;
        RECT 65.795 145.375 67.485 145.545 ;
        RECT 64.820 144.595 64.990 144.725 ;
        RECT 65.795 144.595 65.965 145.375 ;
        RECT 67.655 145.205 67.825 145.895 ;
        RECT 66.325 145.035 67.825 145.205 ;
        RECT 68.015 145.235 68.225 146.025 ;
        RECT 68.395 145.405 68.745 146.025 ;
        RECT 68.915 145.415 69.085 146.195 ;
        RECT 69.615 146.035 69.785 146.265 ;
        RECT 69.255 145.865 69.785 146.035 ;
        RECT 69.255 145.585 69.475 145.865 ;
        RECT 69.955 145.695 70.195 146.095 ;
        RECT 68.915 145.245 69.320 145.415 ;
        RECT 69.655 145.325 70.195 145.695 ;
        RECT 70.365 145.910 70.685 146.265 ;
        RECT 70.930 146.185 71.235 146.645 ;
        RECT 71.405 145.935 71.660 146.465 ;
        RECT 70.365 145.735 70.690 145.910 ;
        RECT 70.365 145.435 71.280 145.735 ;
        RECT 70.540 145.405 71.280 145.435 ;
        RECT 68.015 145.075 68.690 145.235 ;
        RECT 69.150 145.155 69.320 145.245 ;
        RECT 68.015 145.065 68.980 145.075 ;
        RECT 67.655 144.895 67.825 145.035 ;
        RECT 64.400 144.095 64.650 144.555 ;
        RECT 64.820 144.265 65.070 144.595 ;
        RECT 65.285 144.265 65.965 144.595 ;
        RECT 66.135 144.695 67.210 144.865 ;
        RECT 67.655 144.725 68.215 144.895 ;
        RECT 68.520 144.775 68.980 145.065 ;
        RECT 69.150 144.985 70.370 145.155 ;
        RECT 66.135 144.355 66.305 144.695 ;
        RECT 66.540 144.095 66.870 144.525 ;
        RECT 67.040 144.355 67.210 144.695 ;
        RECT 67.505 144.095 67.875 144.555 ;
        RECT 68.045 144.265 68.215 144.725 ;
        RECT 69.150 144.605 69.320 144.985 ;
        RECT 70.540 144.815 70.710 145.405 ;
        RECT 71.450 145.285 71.660 145.935 ;
        RECT 72.110 145.835 72.355 146.440 ;
        RECT 72.575 146.110 73.085 146.645 ;
        RECT 68.450 144.265 69.320 144.605 ;
        RECT 69.910 144.645 70.710 144.815 ;
        RECT 69.490 144.095 69.740 144.555 ;
        RECT 69.910 144.355 70.080 144.645 ;
        RECT 70.260 144.095 70.590 144.475 ;
        RECT 70.930 144.095 71.235 145.235 ;
        RECT 71.405 144.405 71.660 145.285 ;
        RECT 71.835 145.665 73.065 145.835 ;
        RECT 71.835 144.855 72.175 145.665 ;
        RECT 72.345 145.100 73.095 145.290 ;
        RECT 71.835 144.445 72.350 144.855 ;
        RECT 72.585 144.095 72.755 144.855 ;
        RECT 72.925 144.435 73.095 145.100 ;
        RECT 73.265 145.115 73.455 146.475 ;
        RECT 73.625 146.305 73.900 146.475 ;
        RECT 73.625 146.135 73.905 146.305 ;
        RECT 73.625 145.315 73.900 146.135 ;
        RECT 74.090 146.110 74.620 146.475 ;
        RECT 75.045 146.245 75.375 146.645 ;
        RECT 74.445 146.075 74.620 146.110 ;
        RECT 74.105 145.115 74.275 145.915 ;
        RECT 73.265 144.945 74.275 145.115 ;
        RECT 74.445 145.905 75.375 146.075 ;
        RECT 75.545 145.905 75.800 146.475 ;
        RECT 74.445 144.775 74.615 145.905 ;
        RECT 75.205 145.735 75.375 145.905 ;
        RECT 73.490 144.605 74.615 144.775 ;
        RECT 74.785 145.405 74.980 145.735 ;
        RECT 75.205 145.405 75.460 145.735 ;
        RECT 74.785 144.435 74.955 145.405 ;
        RECT 75.630 145.235 75.800 145.905 ;
        RECT 72.925 144.265 74.955 144.435 ;
        RECT 75.125 144.095 75.295 145.235 ;
        RECT 75.465 144.265 75.800 145.235 ;
        RECT 75.980 144.895 76.310 146.475 ;
        RECT 76.480 146.145 76.680 146.645 ;
        RECT 76.940 145.995 77.130 146.310 ;
        RECT 77.300 146.265 78.595 146.435 ;
        RECT 78.765 146.265 79.095 146.645 ;
        RECT 78.425 146.095 78.595 146.265 ;
        RECT 76.480 145.105 76.670 145.975 ;
        RECT 76.940 145.705 77.405 145.995 ;
        RECT 77.585 145.450 78.215 145.965 ;
        RECT 78.425 145.925 79.035 146.095 ;
        RECT 79.265 145.980 79.515 146.475 ;
        RECT 78.865 145.735 79.035 145.925 ;
        RECT 77.585 145.415 77.755 145.450 ;
        RECT 76.940 145.105 77.755 145.415 ;
        RECT 78.525 145.235 78.695 145.735 ;
        RECT 78.035 145.065 78.695 145.235 ;
        RECT 78.865 145.405 79.175 145.735 ;
        RECT 78.035 144.895 78.205 145.065 ;
        RECT 78.865 144.895 79.035 145.405 ;
        RECT 79.345 145.135 79.515 145.980 ;
        RECT 79.685 145.845 79.940 146.645 ;
        RECT 80.115 145.920 80.405 146.645 ;
        RECT 80.850 145.835 81.095 146.440 ;
        RECT 81.315 146.110 81.825 146.645 ;
        RECT 80.575 145.665 81.805 145.835 ;
        RECT 75.980 144.725 78.205 144.895 ;
        RECT 78.375 144.725 79.035 144.895 ;
        RECT 75.980 144.265 76.315 144.725 ;
        RECT 76.485 144.095 76.705 144.555 ;
        RECT 78.375 144.475 78.545 144.725 ;
        RECT 77.235 144.305 78.545 144.475 ;
        RECT 78.715 144.095 79.005 144.555 ;
        RECT 79.205 144.265 79.515 145.135 ;
        RECT 79.685 144.095 79.940 145.235 ;
        RECT 80.115 144.095 80.405 145.260 ;
        RECT 80.575 144.855 80.915 145.665 ;
        RECT 81.085 145.100 81.835 145.290 ;
        RECT 80.575 144.445 81.090 144.855 ;
        RECT 81.325 144.095 81.495 144.855 ;
        RECT 81.665 144.435 81.835 145.100 ;
        RECT 82.005 145.115 82.195 146.475 ;
        RECT 82.365 146.305 82.640 146.475 ;
        RECT 82.365 146.135 82.645 146.305 ;
        RECT 82.365 145.315 82.640 146.135 ;
        RECT 82.830 146.110 83.360 146.475 ;
        RECT 83.785 146.245 84.115 146.645 ;
        RECT 83.185 146.075 83.360 146.110 ;
        RECT 82.845 145.115 83.015 145.915 ;
        RECT 82.005 144.945 83.015 145.115 ;
        RECT 83.185 145.905 84.115 146.075 ;
        RECT 84.285 145.905 84.540 146.475 ;
        RECT 83.185 144.775 83.355 145.905 ;
        RECT 83.945 145.735 84.115 145.905 ;
        RECT 82.230 144.605 83.355 144.775 ;
        RECT 83.525 145.405 83.720 145.735 ;
        RECT 83.945 145.405 84.200 145.735 ;
        RECT 83.525 144.435 83.695 145.405 ;
        RECT 84.370 145.235 84.540 145.905 ;
        RECT 84.715 145.875 86.385 146.645 ;
        RECT 87.180 146.135 87.420 146.645 ;
        RECT 87.600 146.135 87.880 146.465 ;
        RECT 88.110 146.135 88.325 146.645 ;
        RECT 84.715 145.355 85.465 145.875 ;
        RECT 81.665 144.265 83.695 144.435 ;
        RECT 83.865 144.095 84.035 145.235 ;
        RECT 84.205 144.265 84.540 145.235 ;
        RECT 85.635 145.185 86.385 145.705 ;
        RECT 87.075 145.405 87.430 145.965 ;
        RECT 87.600 145.235 87.770 146.135 ;
        RECT 87.940 145.405 88.205 145.965 ;
        RECT 88.495 145.905 89.110 146.475 ;
        RECT 89.775 146.135 90.115 146.645 ;
        RECT 88.455 145.235 88.625 145.735 ;
        RECT 84.715 144.095 86.385 145.185 ;
        RECT 87.200 145.065 88.625 145.235 ;
        RECT 87.200 144.890 87.590 145.065 ;
        RECT 88.075 144.095 88.405 144.895 ;
        RECT 88.795 144.885 89.110 145.905 ;
        RECT 89.785 145.405 90.125 145.965 ;
        RECT 90.295 145.735 90.545 146.465 ;
        RECT 90.870 146.105 91.055 146.465 ;
        RECT 91.235 146.275 91.565 146.645 ;
        RECT 91.745 146.105 91.970 146.465 ;
        RECT 90.870 145.915 92.350 146.105 ;
        RECT 90.295 145.405 90.935 145.735 ;
        RECT 91.115 145.405 91.445 145.735 ;
        RECT 88.575 144.265 89.110 144.885 ;
        RECT 89.940 145.005 91.045 145.205 ;
        RECT 89.940 144.275 90.190 145.005 ;
        RECT 90.360 144.095 90.690 144.825 ;
        RECT 90.860 144.275 91.045 145.005 ;
        RECT 91.215 144.275 91.445 145.405 ;
        RECT 91.625 145.115 91.925 145.735 ;
        RECT 92.135 144.945 92.350 145.915 ;
        RECT 91.625 144.275 92.350 144.945 ;
        RECT 92.995 145.700 93.335 146.475 ;
        RECT 93.505 146.185 93.675 146.645 ;
        RECT 93.915 146.210 94.275 146.475 ;
        RECT 93.915 146.205 94.270 146.210 ;
        RECT 93.915 146.195 94.265 146.205 ;
        RECT 93.915 146.190 94.260 146.195 ;
        RECT 93.915 146.180 94.255 146.190 ;
        RECT 94.905 146.185 95.075 146.645 ;
        RECT 93.915 146.175 94.250 146.180 ;
        RECT 93.915 146.165 94.240 146.175 ;
        RECT 93.915 146.155 94.230 146.165 ;
        RECT 93.915 146.015 94.215 146.155 ;
        RECT 93.505 145.825 94.215 146.015 ;
        RECT 94.405 146.015 94.735 146.095 ;
        RECT 95.245 146.015 95.585 146.475 ;
        RECT 94.405 145.825 95.585 146.015 ;
        RECT 92.995 144.265 93.275 145.700 ;
        RECT 93.505 145.255 93.790 145.825 ;
        RECT 93.975 145.425 94.445 145.655 ;
        RECT 94.615 145.635 94.945 145.655 ;
        RECT 94.615 145.455 95.065 145.635 ;
        RECT 95.255 145.455 95.585 145.655 ;
        RECT 93.505 145.040 94.655 145.255 ;
        RECT 93.445 144.095 94.155 144.870 ;
        RECT 94.325 144.265 94.655 145.040 ;
        RECT 94.850 144.340 95.065 145.455 ;
        RECT 95.355 145.115 95.585 145.455 ;
        RECT 95.245 144.095 95.575 144.815 ;
        RECT 96.675 144.265 97.425 146.475 ;
        RECT 98.550 145.905 99.165 146.475 ;
        RECT 99.335 146.135 99.550 146.645 ;
        RECT 99.780 146.135 100.060 146.465 ;
        RECT 100.240 146.135 100.480 146.645 ;
        RECT 100.980 146.135 101.220 146.645 ;
        RECT 101.400 146.135 101.680 146.465 ;
        RECT 101.910 146.135 102.125 146.645 ;
        RECT 98.550 144.885 98.865 145.905 ;
        RECT 99.035 145.235 99.205 145.735 ;
        RECT 99.455 145.405 99.720 145.965 ;
        RECT 99.890 145.235 100.060 146.135 ;
        RECT 100.230 145.405 100.585 145.965 ;
        RECT 100.875 145.405 101.230 145.965 ;
        RECT 101.400 145.235 101.570 146.135 ;
        RECT 101.740 145.405 102.005 145.965 ;
        RECT 102.295 145.905 102.910 146.475 ;
        RECT 102.255 145.235 102.425 145.735 ;
        RECT 99.035 145.065 100.460 145.235 ;
        RECT 98.550 144.265 99.085 144.885 ;
        RECT 99.255 144.095 99.585 144.895 ;
        RECT 100.070 144.890 100.460 145.065 ;
        RECT 101.000 145.065 102.425 145.235 ;
        RECT 101.000 144.890 101.390 145.065 ;
        RECT 101.875 144.095 102.205 144.895 ;
        RECT 102.595 144.885 102.910 145.905 ;
        RECT 102.375 144.265 102.910 144.885 ;
        RECT 104.035 144.265 104.785 146.475 ;
        RECT 105.875 145.920 106.165 146.645 ;
        RECT 106.580 146.285 108.600 146.475 ;
        RECT 108.770 146.285 109.100 146.645 ;
        RECT 109.630 146.285 109.960 146.645 ;
        RECT 110.490 146.285 110.820 146.645 ;
        RECT 111.350 146.285 111.680 146.645 ;
        RECT 108.370 146.115 108.600 146.285 ;
        RECT 106.395 145.885 108.200 146.115 ;
        RECT 108.370 145.910 112.110 146.115 ;
        RECT 106.395 145.285 106.805 145.885 ;
        RECT 106.975 145.455 108.325 145.715 ;
        RECT 105.875 144.095 106.165 145.260 ;
        RECT 106.395 145.030 108.295 145.285 ;
        RECT 108.535 145.215 108.785 145.740 ;
        RECT 108.955 145.385 110.245 145.660 ;
        RECT 110.755 145.410 112.105 145.715 ;
        RECT 110.755 145.215 111.655 145.410 ;
        RECT 108.535 145.045 111.655 145.215 ;
        RECT 107.080 144.875 108.295 145.030 ;
        RECT 106.580 144.095 106.910 144.850 ;
        RECT 107.080 144.705 110.390 144.875 ;
        RECT 107.080 144.645 108.150 144.705 ;
        RECT 107.080 144.265 107.270 144.645 ;
        RECT 107.440 144.095 107.770 144.475 ;
        RECT 107.940 144.265 108.150 144.645 ;
        RECT 110.560 144.645 111.655 144.815 ;
        RECT 108.320 144.095 108.600 144.535 ;
        RECT 110.560 144.455 110.750 144.645 ;
        RECT 108.770 144.265 110.750 144.455 ;
        RECT 110.920 144.095 111.250 144.475 ;
        RECT 111.420 144.265 111.655 144.645 ;
        RECT 111.825 144.095 112.110 144.910 ;
        RECT 112.320 144.895 112.650 146.475 ;
        RECT 112.820 146.145 113.020 146.645 ;
        RECT 113.280 145.995 113.470 146.310 ;
        RECT 113.640 146.265 114.935 146.435 ;
        RECT 115.105 146.265 115.435 146.645 ;
        RECT 114.765 146.095 114.935 146.265 ;
        RECT 112.820 145.105 113.010 145.975 ;
        RECT 113.280 145.705 113.745 145.995 ;
        RECT 113.925 145.450 114.555 145.965 ;
        RECT 114.765 145.925 115.375 146.095 ;
        RECT 115.605 145.980 115.855 146.475 ;
        RECT 115.205 145.735 115.375 145.925 ;
        RECT 113.925 145.415 114.095 145.450 ;
        RECT 113.280 145.105 114.095 145.415 ;
        RECT 114.865 145.235 115.035 145.735 ;
        RECT 114.375 145.065 115.035 145.235 ;
        RECT 115.205 145.405 115.515 145.735 ;
        RECT 114.375 144.895 114.545 145.065 ;
        RECT 115.205 144.895 115.375 145.405 ;
        RECT 115.685 145.135 115.855 145.980 ;
        RECT 116.025 145.845 116.280 146.645 ;
        RECT 117.385 146.255 119.315 146.445 ;
        RECT 119.485 146.285 122.855 146.475 ;
        RECT 119.145 146.115 119.315 146.255 ;
        RECT 123.390 146.245 123.720 146.645 ;
        RECT 124.250 146.245 124.580 146.645 ;
        RECT 125.115 146.245 125.445 146.645 ;
        RECT 125.955 146.245 126.285 146.645 ;
        RECT 117.375 145.915 118.975 146.085 ;
        RECT 112.320 144.725 114.545 144.895 ;
        RECT 114.715 144.725 115.375 144.895 ;
        RECT 112.320 144.265 112.655 144.725 ;
        RECT 112.825 144.095 113.045 144.555 ;
        RECT 114.715 144.475 114.885 144.725 ;
        RECT 113.575 144.305 114.885 144.475 ;
        RECT 115.055 144.095 115.345 144.555 ;
        RECT 115.545 144.265 115.855 145.135 ;
        RECT 116.025 144.095 116.280 145.235 ;
        RECT 117.375 145.215 117.665 145.915 ;
        RECT 119.145 145.905 121.075 146.115 ;
        RECT 121.265 145.825 126.730 146.075 ;
        RECT 127.770 145.835 128.015 146.440 ;
        RECT 128.235 146.110 128.745 146.645 ;
        RECT 127.495 145.665 128.725 145.835 ;
        RECT 117.835 145.385 119.045 145.655 ;
        RECT 119.230 145.385 120.840 145.655 ;
        RECT 121.105 145.385 122.745 145.655 ;
        RECT 123.400 145.385 124.615 145.655 ;
        RECT 125.110 145.390 126.865 145.655 ;
        RECT 122.955 145.215 123.125 145.285 ;
        RECT 117.375 145.045 124.680 145.215 ;
        RECT 117.375 144.265 117.650 145.045 ;
        RECT 117.820 144.095 118.135 144.875 ;
        RECT 118.305 144.265 118.485 145.045 ;
        RECT 118.680 144.095 118.965 144.875 ;
        RECT 119.135 144.265 119.325 145.045 ;
        RECT 119.495 144.095 119.805 144.875 ;
        RECT 119.975 144.265 120.165 145.045 ;
        RECT 120.335 144.095 120.645 144.875 ;
        RECT 120.815 144.265 121.005 145.045 ;
        RECT 121.365 144.095 121.690 144.875 ;
        RECT 121.860 144.265 122.050 145.045 ;
        RECT 122.220 144.095 122.510 144.875 ;
        RECT 122.700 144.265 122.890 145.045 ;
        RECT 123.075 144.460 123.405 144.875 ;
        RECT 123.575 144.630 123.770 145.045 ;
        RECT 124.335 145.010 124.680 145.045 ;
        RECT 125.335 145.045 126.370 145.215 ;
        RECT 125.335 144.840 125.525 145.045 ;
        RECT 123.995 144.670 125.525 144.840 ;
        RECT 123.995 144.460 124.295 144.670 ;
        RECT 123.075 144.265 124.295 144.460 ;
        RECT 124.845 144.095 125.175 144.500 ;
        RECT 125.345 144.265 125.525 144.670 ;
        RECT 125.700 144.095 126.010 144.875 ;
        RECT 126.180 144.265 126.370 145.045 ;
        RECT 126.555 144.095 126.865 145.195 ;
        RECT 127.495 144.855 127.835 145.665 ;
        RECT 128.005 145.100 128.755 145.290 ;
        RECT 127.495 144.445 128.010 144.855 ;
        RECT 128.245 144.095 128.415 144.855 ;
        RECT 128.585 144.435 128.755 145.100 ;
        RECT 128.925 145.115 129.115 146.475 ;
        RECT 129.285 146.305 129.560 146.475 ;
        RECT 129.285 146.135 129.565 146.305 ;
        RECT 129.285 145.315 129.560 146.135 ;
        RECT 129.750 146.110 130.280 146.475 ;
        RECT 130.705 146.245 131.035 146.645 ;
        RECT 130.105 146.075 130.280 146.110 ;
        RECT 129.765 145.115 129.935 145.915 ;
        RECT 128.925 144.945 129.935 145.115 ;
        RECT 130.105 145.905 131.035 146.075 ;
        RECT 131.205 145.905 131.460 146.475 ;
        RECT 131.635 145.920 131.925 146.645 ;
        RECT 132.120 146.255 132.450 146.645 ;
        RECT 132.620 146.085 132.845 146.465 ;
        RECT 130.105 144.775 130.275 145.905 ;
        RECT 130.865 145.735 131.035 145.905 ;
        RECT 129.150 144.605 130.275 144.775 ;
        RECT 130.445 145.405 130.640 145.735 ;
        RECT 130.865 145.405 131.120 145.735 ;
        RECT 130.445 144.435 130.615 145.405 ;
        RECT 131.290 145.235 131.460 145.905 ;
        RECT 132.105 145.405 132.345 146.055 ;
        RECT 132.515 145.905 132.845 146.085 ;
        RECT 128.585 144.265 130.615 144.435 ;
        RECT 130.785 144.095 130.955 145.235 ;
        RECT 131.125 144.265 131.460 145.235 ;
        RECT 131.635 144.095 131.925 145.260 ;
        RECT 132.515 145.235 132.690 145.905 ;
        RECT 133.045 145.735 133.275 146.355 ;
        RECT 133.455 145.915 133.755 146.645 ;
        RECT 134.400 146.095 134.655 146.385 ;
        RECT 134.825 146.265 135.155 146.645 ;
        RECT 134.400 145.925 135.150 146.095 ;
        RECT 132.860 145.405 133.275 145.735 ;
        RECT 133.455 145.405 133.750 145.735 ;
        RECT 132.105 145.045 132.690 145.235 ;
        RECT 132.105 144.275 132.380 145.045 ;
        RECT 132.860 144.875 133.755 145.205 ;
        RECT 134.400 145.105 134.750 145.755 ;
        RECT 134.920 144.935 135.150 145.925 ;
        RECT 132.550 144.705 133.755 144.875 ;
        RECT 132.550 144.275 132.880 144.705 ;
        RECT 133.050 144.095 133.245 144.535 ;
        RECT 133.425 144.275 133.755 144.705 ;
        RECT 134.400 144.765 135.150 144.935 ;
        RECT 134.400 144.265 134.655 144.765 ;
        RECT 134.825 144.095 135.155 144.595 ;
        RECT 135.325 144.265 135.495 146.385 ;
        RECT 135.855 146.285 136.185 146.645 ;
        RECT 136.355 146.255 136.850 146.425 ;
        RECT 137.055 146.255 137.910 146.425 ;
        RECT 135.725 145.065 136.185 146.115 ;
        RECT 135.665 144.280 135.990 145.065 ;
        RECT 136.355 144.895 136.525 146.255 ;
        RECT 136.695 145.345 137.045 145.965 ;
        RECT 137.215 145.745 137.570 145.965 ;
        RECT 137.215 145.155 137.385 145.745 ;
        RECT 137.740 145.545 137.910 146.255 ;
        RECT 138.785 146.185 139.115 146.645 ;
        RECT 139.325 146.285 139.675 146.455 ;
        RECT 138.115 145.715 138.905 145.965 ;
        RECT 139.325 145.895 139.585 146.285 ;
        RECT 139.895 146.195 140.845 146.475 ;
        RECT 141.015 146.205 141.205 146.645 ;
        RECT 141.375 146.265 142.445 146.435 ;
        RECT 139.075 145.545 139.245 145.725 ;
        RECT 136.355 144.725 136.750 144.895 ;
        RECT 136.920 144.765 137.385 145.155 ;
        RECT 137.555 145.375 139.245 145.545 ;
        RECT 136.580 144.595 136.750 144.725 ;
        RECT 137.555 144.595 137.725 145.375 ;
        RECT 139.415 145.205 139.585 145.895 ;
        RECT 138.085 145.035 139.585 145.205 ;
        RECT 139.775 145.235 139.985 146.025 ;
        RECT 140.155 145.405 140.505 146.025 ;
        RECT 140.675 145.415 140.845 146.195 ;
        RECT 141.375 146.035 141.545 146.265 ;
        RECT 141.015 145.865 141.545 146.035 ;
        RECT 141.015 145.585 141.235 145.865 ;
        RECT 141.715 145.695 141.955 146.095 ;
        RECT 140.675 145.245 141.080 145.415 ;
        RECT 141.415 145.325 141.955 145.695 ;
        RECT 142.125 145.910 142.445 146.265 ;
        RECT 142.690 146.185 142.995 146.645 ;
        RECT 143.165 145.935 143.420 146.465 ;
        RECT 142.125 145.735 142.450 145.910 ;
        RECT 142.125 145.435 143.040 145.735 ;
        RECT 142.300 145.405 143.040 145.435 ;
        RECT 139.775 145.075 140.450 145.235 ;
        RECT 140.910 145.155 141.080 145.245 ;
        RECT 139.775 145.065 140.740 145.075 ;
        RECT 139.415 144.895 139.585 145.035 ;
        RECT 136.160 144.095 136.410 144.555 ;
        RECT 136.580 144.265 136.830 144.595 ;
        RECT 137.045 144.265 137.725 144.595 ;
        RECT 137.895 144.695 138.970 144.865 ;
        RECT 139.415 144.725 139.975 144.895 ;
        RECT 140.280 144.775 140.740 145.065 ;
        RECT 140.910 144.985 142.130 145.155 ;
        RECT 137.895 144.355 138.065 144.695 ;
        RECT 138.300 144.095 138.630 144.525 ;
        RECT 138.800 144.355 138.970 144.695 ;
        RECT 139.265 144.095 139.635 144.555 ;
        RECT 139.805 144.265 139.975 144.725 ;
        RECT 140.910 144.605 141.080 144.985 ;
        RECT 142.300 144.815 142.470 145.405 ;
        RECT 143.210 145.285 143.420 145.935 ;
        RECT 140.210 144.265 141.080 144.605 ;
        RECT 141.670 144.645 142.470 144.815 ;
        RECT 141.250 144.095 141.500 144.555 ;
        RECT 141.670 144.355 141.840 144.645 ;
        RECT 142.020 144.095 142.350 144.475 ;
        RECT 142.690 144.095 142.995 145.235 ;
        RECT 143.165 144.405 143.420 145.285 ;
        RECT 143.595 145.970 143.855 146.475 ;
        RECT 144.035 146.265 144.365 146.645 ;
        RECT 144.545 146.095 144.715 146.475 ;
        RECT 143.595 145.170 143.765 145.970 ;
        RECT 144.050 145.925 144.715 146.095 ;
        RECT 144.975 145.970 145.235 146.475 ;
        RECT 145.415 146.265 145.745 146.645 ;
        RECT 145.925 146.095 146.095 146.475 ;
        RECT 146.355 146.100 151.700 146.645 ;
        RECT 144.050 145.670 144.220 145.925 ;
        RECT 143.935 145.340 144.220 145.670 ;
        RECT 144.455 145.375 144.785 145.745 ;
        RECT 144.050 145.195 144.220 145.340 ;
        RECT 143.595 144.265 143.865 145.170 ;
        RECT 144.050 145.025 144.715 145.195 ;
        RECT 144.035 144.095 144.365 144.855 ;
        RECT 144.545 144.265 144.715 145.025 ;
        RECT 144.975 145.170 145.145 145.970 ;
        RECT 145.430 145.925 146.095 146.095 ;
        RECT 145.430 145.670 145.600 145.925 ;
        RECT 145.315 145.340 145.600 145.670 ;
        RECT 145.835 145.375 146.165 145.745 ;
        RECT 145.430 145.195 145.600 145.340 ;
        RECT 147.940 145.270 148.280 146.100 ;
        RECT 151.875 145.875 155.385 146.645 ;
        RECT 155.555 145.895 156.765 146.645 ;
        RECT 156.935 145.895 158.145 146.645 ;
        RECT 144.975 144.265 145.245 145.170 ;
        RECT 145.430 145.025 146.095 145.195 ;
        RECT 145.415 144.095 145.745 144.855 ;
        RECT 145.925 144.265 146.095 145.025 ;
        RECT 149.760 144.530 150.110 145.780 ;
        RECT 151.875 145.355 153.525 145.875 ;
        RECT 153.695 145.185 155.385 145.705 ;
        RECT 155.555 145.355 156.075 145.895 ;
        RECT 156.245 145.185 156.765 145.725 ;
        RECT 146.355 144.095 151.700 144.530 ;
        RECT 151.875 144.095 155.385 145.185 ;
        RECT 155.555 144.095 156.765 145.185 ;
        RECT 156.935 145.185 157.455 145.725 ;
        RECT 157.625 145.355 158.145 145.895 ;
        RECT 156.935 144.095 158.145 145.185 ;
        RECT 2.750 143.925 158.230 144.095 ;
        RECT 2.835 142.835 4.045 143.925 ;
        RECT 4.305 143.255 4.475 143.755 ;
        RECT 4.645 143.425 4.975 143.925 ;
        RECT 4.305 143.085 4.970 143.255 ;
        RECT 2.835 142.125 3.355 142.665 ;
        RECT 3.525 142.295 4.045 142.835 ;
        RECT 4.220 142.265 4.570 142.915 ;
        RECT 2.835 141.375 4.045 142.125 ;
        RECT 4.740 142.095 4.970 143.085 ;
        RECT 4.305 141.925 4.970 142.095 ;
        RECT 4.305 141.635 4.475 141.925 ;
        RECT 4.645 141.375 4.975 141.755 ;
        RECT 5.145 141.635 5.370 143.755 ;
        RECT 5.585 143.425 5.915 143.925 ;
        RECT 6.085 143.255 6.255 143.755 ;
        RECT 6.490 143.540 7.320 143.710 ;
        RECT 7.560 143.545 7.940 143.925 ;
        RECT 5.560 143.085 6.255 143.255 ;
        RECT 5.560 142.115 5.730 143.085 ;
        RECT 5.900 142.295 6.310 142.915 ;
        RECT 6.480 142.865 6.980 143.245 ;
        RECT 5.560 141.925 6.255 142.115 ;
        RECT 6.480 141.995 6.700 142.865 ;
        RECT 7.150 142.695 7.320 143.540 ;
        RECT 8.120 143.375 8.290 143.665 ;
        RECT 8.460 143.545 8.790 143.925 ;
        RECT 9.260 143.455 9.890 143.705 ;
        RECT 10.070 143.545 10.490 143.925 ;
        RECT 9.720 143.375 9.890 143.455 ;
        RECT 10.690 143.375 10.930 143.665 ;
        RECT 7.490 143.125 8.860 143.375 ;
        RECT 7.490 142.865 7.740 143.125 ;
        RECT 8.250 142.695 8.500 142.855 ;
        RECT 7.150 142.525 8.500 142.695 ;
        RECT 7.150 142.485 7.570 142.525 ;
        RECT 6.880 141.935 7.230 142.305 ;
        RECT 5.585 141.375 5.915 141.755 ;
        RECT 6.085 141.595 6.255 141.925 ;
        RECT 7.400 141.755 7.570 142.485 ;
        RECT 8.670 142.355 8.860 143.125 ;
        RECT 7.740 142.025 8.150 142.355 ;
        RECT 8.440 142.015 8.860 142.355 ;
        RECT 9.030 142.945 9.550 143.255 ;
        RECT 9.720 143.205 10.930 143.375 ;
        RECT 11.160 143.235 11.490 143.925 ;
        RECT 9.030 142.185 9.200 142.945 ;
        RECT 9.370 142.355 9.550 142.765 ;
        RECT 9.720 142.695 9.890 143.205 ;
        RECT 11.660 143.055 11.830 143.665 ;
        RECT 12.100 143.205 12.430 143.715 ;
        RECT 11.660 143.035 11.980 143.055 ;
        RECT 10.060 142.865 11.980 143.035 ;
        RECT 9.720 142.525 11.620 142.695 ;
        RECT 9.950 142.185 10.280 142.305 ;
        RECT 9.030 142.015 10.280 142.185 ;
        RECT 6.555 141.555 7.570 141.755 ;
        RECT 7.740 141.375 8.150 141.815 ;
        RECT 8.440 141.585 8.690 142.015 ;
        RECT 8.890 141.375 9.210 141.835 ;
        RECT 10.450 141.765 10.620 142.525 ;
        RECT 11.290 142.465 11.620 142.525 ;
        RECT 10.810 142.295 11.140 142.355 ;
        RECT 10.810 142.025 11.470 142.295 ;
        RECT 11.790 141.970 11.980 142.865 ;
        RECT 9.770 141.595 10.620 141.765 ;
        RECT 10.820 141.375 11.480 141.855 ;
        RECT 11.660 141.640 11.980 141.970 ;
        RECT 12.180 142.615 12.430 143.205 ;
        RECT 12.610 143.125 12.895 143.925 ;
        RECT 13.075 143.585 13.330 143.615 ;
        RECT 13.075 143.415 13.415 143.585 ;
        RECT 13.075 142.945 13.330 143.415 ;
        RECT 12.180 142.285 12.980 142.615 ;
        RECT 12.180 141.635 12.430 142.285 ;
        RECT 13.150 142.085 13.330 142.945 ;
        RECT 12.610 141.375 12.895 141.835 ;
        RECT 13.075 141.555 13.330 142.085 ;
        RECT 13.875 142.850 14.145 143.755 ;
        RECT 14.315 143.165 14.645 143.925 ;
        RECT 14.825 142.995 14.995 143.755 ;
        RECT 13.875 142.050 14.045 142.850 ;
        RECT 14.330 142.825 14.995 142.995 ;
        RECT 14.330 142.680 14.500 142.825 ;
        RECT 15.715 142.760 16.005 143.925 ;
        RECT 16.180 142.785 16.515 143.755 ;
        RECT 16.685 142.785 16.855 143.925 ;
        RECT 17.025 143.585 19.055 143.755 ;
        RECT 14.215 142.350 14.500 142.680 ;
        RECT 14.330 142.095 14.500 142.350 ;
        RECT 14.735 142.275 15.065 142.645 ;
        RECT 16.180 142.115 16.350 142.785 ;
        RECT 17.025 142.615 17.195 143.585 ;
        RECT 16.520 142.285 16.775 142.615 ;
        RECT 17.000 142.285 17.195 142.615 ;
        RECT 17.365 143.245 18.490 143.415 ;
        RECT 16.605 142.115 16.775 142.285 ;
        RECT 17.365 142.115 17.535 143.245 ;
        RECT 13.875 141.545 14.135 142.050 ;
        RECT 14.330 141.925 14.995 142.095 ;
        RECT 14.315 141.375 14.645 141.755 ;
        RECT 14.825 141.545 14.995 141.925 ;
        RECT 15.715 141.375 16.005 142.100 ;
        RECT 16.180 141.545 16.435 142.115 ;
        RECT 16.605 141.945 17.535 142.115 ;
        RECT 17.705 142.905 18.715 143.075 ;
        RECT 17.705 142.105 17.875 142.905 ;
        RECT 18.080 142.225 18.355 142.705 ;
        RECT 18.075 142.055 18.355 142.225 ;
        RECT 17.360 141.910 17.535 141.945 ;
        RECT 16.605 141.375 16.935 141.775 ;
        RECT 17.360 141.545 17.890 141.910 ;
        RECT 18.080 141.545 18.355 142.055 ;
        RECT 18.525 141.545 18.715 142.905 ;
        RECT 18.885 142.920 19.055 143.585 ;
        RECT 19.225 143.165 19.395 143.925 ;
        RECT 19.630 143.165 20.145 143.575 ;
        RECT 18.885 142.730 19.635 142.920 ;
        RECT 19.805 142.355 20.145 143.165 ;
        RECT 20.815 142.975 21.105 143.745 ;
        RECT 21.675 143.385 21.935 143.745 ;
        RECT 22.105 143.555 22.435 143.925 ;
        RECT 22.605 143.385 22.865 143.745 ;
        RECT 21.675 143.155 22.865 143.385 ;
        RECT 23.055 143.205 23.385 143.925 ;
        RECT 23.555 142.975 23.820 143.745 ;
        RECT 20.815 142.795 23.310 142.975 ;
        RECT 18.915 142.185 20.145 142.355 ;
        RECT 20.785 142.285 21.055 142.615 ;
        RECT 21.235 142.285 21.670 142.615 ;
        RECT 21.850 142.285 22.425 142.615 ;
        RECT 22.605 142.285 22.885 142.615 ;
        RECT 18.895 141.375 19.405 141.910 ;
        RECT 19.625 141.580 19.870 142.185 ;
        RECT 23.085 142.105 23.310 142.795 ;
        RECT 20.825 141.915 23.310 142.105 ;
        RECT 20.825 141.555 21.050 141.915 ;
        RECT 21.230 141.375 21.560 141.745 ;
        RECT 21.740 141.555 21.995 141.915 ;
        RECT 22.560 141.375 23.305 141.745 ;
        RECT 23.485 141.555 23.820 142.975 ;
        RECT 24.085 142.995 24.255 143.755 ;
        RECT 24.435 143.165 24.765 143.925 ;
        RECT 24.085 142.825 24.750 142.995 ;
        RECT 24.935 142.850 25.205 143.755 ;
        RECT 24.580 142.680 24.750 142.825 ;
        RECT 24.015 142.275 24.345 142.645 ;
        RECT 24.580 142.350 24.865 142.680 ;
        RECT 24.580 142.095 24.750 142.350 ;
        RECT 24.085 141.925 24.750 142.095 ;
        RECT 25.035 142.050 25.205 142.850 ;
        RECT 24.085 141.545 24.255 141.925 ;
        RECT 24.435 141.375 24.765 141.755 ;
        RECT 24.945 141.545 25.205 142.050 ;
        RECT 25.835 142.785 26.220 143.755 ;
        RECT 26.390 143.465 26.715 143.925 ;
        RECT 27.235 143.295 27.515 143.755 ;
        RECT 26.390 143.075 27.515 143.295 ;
        RECT 25.835 142.115 26.115 142.785 ;
        RECT 26.390 142.615 26.840 143.075 ;
        RECT 27.705 142.905 28.105 143.755 ;
        RECT 28.505 143.465 28.775 143.925 ;
        RECT 28.945 143.295 29.230 143.755 ;
        RECT 26.285 142.285 26.840 142.615 ;
        RECT 27.010 142.345 28.105 142.905 ;
        RECT 26.390 142.175 26.840 142.285 ;
        RECT 25.835 141.545 26.220 142.115 ;
        RECT 26.390 142.005 27.515 142.175 ;
        RECT 26.390 141.375 26.715 141.835 ;
        RECT 27.235 141.545 27.515 142.005 ;
        RECT 27.705 141.545 28.105 142.345 ;
        RECT 28.275 143.075 29.230 143.295 ;
        RECT 29.520 143.255 29.775 143.755 ;
        RECT 29.945 143.425 30.275 143.925 ;
        RECT 29.520 143.085 30.270 143.255 ;
        RECT 28.275 142.175 28.485 143.075 ;
        RECT 28.655 142.345 29.345 142.905 ;
        RECT 29.520 142.265 29.870 142.915 ;
        RECT 28.275 142.005 29.230 142.175 ;
        RECT 30.040 142.095 30.270 143.085 ;
        RECT 28.505 141.375 28.775 141.835 ;
        RECT 28.945 141.545 29.230 142.005 ;
        RECT 29.520 141.925 30.270 142.095 ;
        RECT 29.520 141.635 29.775 141.925 ;
        RECT 29.945 141.375 30.275 141.755 ;
        RECT 30.445 141.635 30.615 143.755 ;
        RECT 30.785 142.955 31.110 143.740 ;
        RECT 31.280 143.465 31.530 143.925 ;
        RECT 31.700 143.425 31.950 143.755 ;
        RECT 32.165 143.425 32.845 143.755 ;
        RECT 31.700 143.295 31.870 143.425 ;
        RECT 31.475 143.125 31.870 143.295 ;
        RECT 30.845 141.905 31.305 142.955 ;
        RECT 31.475 141.765 31.645 143.125 ;
        RECT 32.040 142.865 32.505 143.255 ;
        RECT 31.815 142.055 32.165 142.675 ;
        RECT 32.335 142.275 32.505 142.865 ;
        RECT 32.675 142.645 32.845 143.425 ;
        RECT 33.015 143.325 33.185 143.665 ;
        RECT 33.420 143.495 33.750 143.925 ;
        RECT 33.920 143.325 34.090 143.665 ;
        RECT 34.385 143.465 34.755 143.925 ;
        RECT 33.015 143.155 34.090 143.325 ;
        RECT 34.925 143.295 35.095 143.755 ;
        RECT 35.330 143.415 36.200 143.755 ;
        RECT 36.370 143.465 36.620 143.925 ;
        RECT 34.535 143.125 35.095 143.295 ;
        RECT 34.535 142.985 34.705 143.125 ;
        RECT 33.205 142.815 34.705 142.985 ;
        RECT 35.400 142.955 35.860 143.245 ;
        RECT 32.675 142.475 34.365 142.645 ;
        RECT 32.335 142.055 32.690 142.275 ;
        RECT 32.860 141.765 33.030 142.475 ;
        RECT 33.235 142.055 34.025 142.305 ;
        RECT 34.195 142.295 34.365 142.475 ;
        RECT 34.535 142.125 34.705 142.815 ;
        RECT 30.975 141.375 31.305 141.735 ;
        RECT 31.475 141.595 31.970 141.765 ;
        RECT 32.175 141.595 33.030 141.765 ;
        RECT 33.905 141.375 34.235 141.835 ;
        RECT 34.445 141.735 34.705 142.125 ;
        RECT 34.895 142.945 35.860 142.955 ;
        RECT 36.030 143.035 36.200 143.415 ;
        RECT 36.790 143.375 36.960 143.665 ;
        RECT 37.140 143.545 37.470 143.925 ;
        RECT 36.790 143.205 37.590 143.375 ;
        RECT 34.895 142.785 35.570 142.945 ;
        RECT 36.030 142.865 37.250 143.035 ;
        RECT 34.895 141.995 35.105 142.785 ;
        RECT 36.030 142.775 36.200 142.865 ;
        RECT 35.275 141.995 35.625 142.615 ;
        RECT 35.795 142.605 36.200 142.775 ;
        RECT 35.795 141.825 35.965 142.605 ;
        RECT 36.135 142.155 36.355 142.435 ;
        RECT 36.535 142.325 37.075 142.695 ;
        RECT 37.420 142.615 37.590 143.205 ;
        RECT 37.810 142.785 38.115 143.925 ;
        RECT 38.285 142.735 38.540 143.615 ;
        RECT 38.735 143.035 38.995 143.745 ;
        RECT 39.165 143.215 39.495 143.925 ;
        RECT 39.665 143.035 39.895 143.745 ;
        RECT 38.735 142.795 39.895 143.035 ;
        RECT 40.075 143.015 40.345 143.745 ;
        RECT 40.525 143.195 40.865 143.925 ;
        RECT 40.075 142.795 40.845 143.015 ;
        RECT 37.420 142.585 38.160 142.615 ;
        RECT 36.135 141.985 36.665 142.155 ;
        RECT 34.445 141.565 34.795 141.735 ;
        RECT 35.015 141.545 35.965 141.825 ;
        RECT 36.135 141.375 36.325 141.815 ;
        RECT 36.495 141.755 36.665 141.985 ;
        RECT 36.835 141.925 37.075 142.325 ;
        RECT 37.245 142.285 38.160 142.585 ;
        RECT 37.245 142.110 37.570 142.285 ;
        RECT 37.245 141.755 37.565 142.110 ;
        RECT 38.330 142.085 38.540 142.735 ;
        RECT 38.725 142.285 39.025 142.615 ;
        RECT 39.205 142.305 39.730 142.615 ;
        RECT 39.910 142.305 40.375 142.615 ;
        RECT 36.495 141.585 37.565 141.755 ;
        RECT 37.810 141.375 38.115 141.835 ;
        RECT 38.285 141.555 38.540 142.085 ;
        RECT 38.735 141.375 39.025 142.105 ;
        RECT 39.205 141.665 39.435 142.305 ;
        RECT 40.555 142.125 40.845 142.795 ;
        RECT 39.615 141.925 40.845 142.125 ;
        RECT 39.615 141.555 39.925 141.925 ;
        RECT 40.105 141.375 40.775 141.745 ;
        RECT 41.035 141.555 41.295 143.745 ;
        RECT 41.475 142.760 41.765 143.925 ;
        RECT 41.940 142.785 42.275 143.755 ;
        RECT 42.445 142.785 42.615 143.925 ;
        RECT 42.785 143.585 44.815 143.755 ;
        RECT 41.940 142.115 42.110 142.785 ;
        RECT 42.785 142.615 42.955 143.585 ;
        RECT 42.280 142.285 42.535 142.615 ;
        RECT 42.760 142.285 42.955 142.615 ;
        RECT 43.125 143.245 44.250 143.415 ;
        RECT 42.365 142.115 42.535 142.285 ;
        RECT 43.125 142.115 43.295 143.245 ;
        RECT 41.475 141.375 41.765 142.100 ;
        RECT 41.940 141.545 42.195 142.115 ;
        RECT 42.365 141.945 43.295 142.115 ;
        RECT 43.465 142.905 44.475 143.075 ;
        RECT 43.465 142.105 43.635 142.905 ;
        RECT 43.120 141.910 43.295 141.945 ;
        RECT 42.365 141.375 42.695 141.775 ;
        RECT 43.120 141.545 43.650 141.910 ;
        RECT 43.840 141.885 44.115 142.705 ;
        RECT 43.835 141.715 44.115 141.885 ;
        RECT 43.840 141.545 44.115 141.715 ;
        RECT 44.285 141.545 44.475 142.905 ;
        RECT 44.645 142.920 44.815 143.585 ;
        RECT 44.985 143.165 45.155 143.925 ;
        RECT 45.390 143.165 45.905 143.575 ;
        RECT 44.645 142.730 45.395 142.920 ;
        RECT 45.565 142.355 45.905 143.165 ;
        RECT 44.675 142.185 45.905 142.355 ;
        RECT 46.075 142.785 46.460 143.755 ;
        RECT 46.630 143.465 46.955 143.925 ;
        RECT 47.475 143.295 47.755 143.755 ;
        RECT 46.630 143.075 47.755 143.295 ;
        RECT 44.655 141.375 45.165 141.910 ;
        RECT 45.385 141.580 45.630 142.185 ;
        RECT 46.075 142.115 46.355 142.785 ;
        RECT 46.630 142.615 47.080 143.075 ;
        RECT 47.945 142.905 48.345 143.755 ;
        RECT 48.745 143.465 49.015 143.925 ;
        RECT 49.185 143.295 49.470 143.755 ;
        RECT 46.525 142.285 47.080 142.615 ;
        RECT 47.250 142.345 48.345 142.905 ;
        RECT 46.630 142.175 47.080 142.285 ;
        RECT 46.075 141.545 46.460 142.115 ;
        RECT 46.630 142.005 47.755 142.175 ;
        RECT 46.630 141.375 46.955 141.835 ;
        RECT 47.475 141.545 47.755 142.005 ;
        RECT 47.945 141.545 48.345 142.345 ;
        RECT 48.515 143.075 49.470 143.295 ;
        RECT 48.515 142.175 48.725 143.075 ;
        RECT 49.845 142.915 50.015 143.755 ;
        RECT 50.185 143.585 51.355 143.755 ;
        RECT 50.185 143.085 50.515 143.585 ;
        RECT 51.025 143.545 51.355 143.585 ;
        RECT 51.545 143.505 51.900 143.925 ;
        RECT 50.685 143.325 50.915 143.415 ;
        RECT 52.070 143.325 52.320 143.755 ;
        RECT 50.685 143.085 52.320 143.325 ;
        RECT 52.490 143.165 52.820 143.925 ;
        RECT 52.990 143.085 53.245 143.755 ;
        RECT 48.895 142.345 49.585 142.905 ;
        RECT 49.845 142.745 52.905 142.915 ;
        RECT 49.760 142.365 50.110 142.575 ;
        RECT 50.280 142.365 50.725 142.565 ;
        RECT 50.895 142.365 51.370 142.565 ;
        RECT 48.515 142.005 49.470 142.175 ;
        RECT 48.745 141.375 49.015 141.835 ;
        RECT 49.185 141.545 49.470 142.005 ;
        RECT 49.845 142.025 50.910 142.195 ;
        RECT 49.845 141.545 50.015 142.025 ;
        RECT 50.185 141.375 50.515 141.855 ;
        RECT 50.740 141.795 50.910 142.025 ;
        RECT 51.090 141.965 51.370 142.365 ;
        RECT 51.640 142.365 51.970 142.565 ;
        RECT 52.140 142.365 52.505 142.565 ;
        RECT 51.640 141.965 51.925 142.365 ;
        RECT 52.735 142.195 52.905 142.745 ;
        RECT 52.105 142.025 52.905 142.195 ;
        RECT 52.105 141.795 52.275 142.025 ;
        RECT 53.075 141.955 53.245 143.085 ;
        RECT 53.435 143.165 53.950 143.575 ;
        RECT 54.185 143.165 54.355 143.925 ;
        RECT 54.525 143.585 56.555 143.755 ;
        RECT 53.435 142.355 53.775 143.165 ;
        RECT 54.525 142.920 54.695 143.585 ;
        RECT 55.090 143.245 56.215 143.415 ;
        RECT 53.945 142.730 54.695 142.920 ;
        RECT 54.865 142.905 55.875 143.075 ;
        RECT 53.435 142.185 54.665 142.355 ;
        RECT 53.060 141.875 53.245 141.955 ;
        RECT 50.740 141.545 52.275 141.795 ;
        RECT 52.445 141.375 52.775 141.855 ;
        RECT 52.990 141.545 53.245 141.875 ;
        RECT 53.710 141.580 53.955 142.185 ;
        RECT 54.175 141.375 54.685 141.910 ;
        RECT 54.865 141.545 55.055 142.905 ;
        RECT 55.225 142.225 55.500 142.705 ;
        RECT 55.225 142.055 55.505 142.225 ;
        RECT 55.705 142.105 55.875 142.905 ;
        RECT 56.045 142.115 56.215 143.245 ;
        RECT 56.385 142.615 56.555 143.585 ;
        RECT 56.725 142.785 56.895 143.925 ;
        RECT 57.065 142.785 57.400 143.755 ;
        RECT 57.950 142.945 58.205 143.615 ;
        RECT 58.385 143.125 58.670 143.925 ;
        RECT 58.850 143.205 59.180 143.715 ;
        RECT 57.950 142.905 58.130 142.945 ;
        RECT 56.385 142.285 56.580 142.615 ;
        RECT 56.805 142.285 57.060 142.615 ;
        RECT 56.805 142.115 56.975 142.285 ;
        RECT 57.230 142.115 57.400 142.785 ;
        RECT 57.865 142.735 58.130 142.905 ;
        RECT 55.225 141.545 55.500 142.055 ;
        RECT 56.045 141.945 56.975 142.115 ;
        RECT 56.045 141.910 56.220 141.945 ;
        RECT 55.690 141.545 56.220 141.910 ;
        RECT 56.645 141.375 56.975 141.775 ;
        RECT 57.145 141.545 57.400 142.115 ;
        RECT 57.950 142.085 58.130 142.735 ;
        RECT 58.850 142.615 59.100 143.205 ;
        RECT 59.450 143.055 59.620 143.665 ;
        RECT 59.790 143.235 60.120 143.925 ;
        RECT 60.350 143.375 60.590 143.665 ;
        RECT 60.790 143.545 61.210 143.925 ;
        RECT 61.390 143.455 62.020 143.705 ;
        RECT 62.490 143.545 62.820 143.925 ;
        RECT 61.390 143.375 61.560 143.455 ;
        RECT 62.990 143.375 63.160 143.665 ;
        RECT 63.340 143.545 63.720 143.925 ;
        RECT 63.960 143.540 64.790 143.710 ;
        RECT 60.350 143.205 61.560 143.375 ;
        RECT 58.300 142.285 59.100 142.615 ;
        RECT 57.950 141.555 58.205 142.085 ;
        RECT 58.385 141.375 58.670 141.835 ;
        RECT 58.850 141.635 59.100 142.285 ;
        RECT 59.300 143.035 59.620 143.055 ;
        RECT 59.300 142.865 61.220 143.035 ;
        RECT 59.300 141.970 59.490 142.865 ;
        RECT 61.390 142.695 61.560 143.205 ;
        RECT 61.730 142.945 62.250 143.255 ;
        RECT 59.660 142.525 61.560 142.695 ;
        RECT 59.660 142.465 59.990 142.525 ;
        RECT 60.140 142.295 60.470 142.355 ;
        RECT 59.810 142.025 60.470 142.295 ;
        RECT 59.300 141.640 59.620 141.970 ;
        RECT 59.800 141.375 60.460 141.855 ;
        RECT 60.660 141.765 60.830 142.525 ;
        RECT 61.730 142.355 61.910 142.765 ;
        RECT 61.000 142.185 61.330 142.305 ;
        RECT 62.080 142.185 62.250 142.945 ;
        RECT 61.000 142.015 62.250 142.185 ;
        RECT 62.420 143.125 63.790 143.375 ;
        RECT 62.420 142.355 62.610 143.125 ;
        RECT 63.540 142.865 63.790 143.125 ;
        RECT 62.780 142.695 63.030 142.855 ;
        RECT 63.960 142.695 64.130 143.540 ;
        RECT 65.025 143.255 65.195 143.755 ;
        RECT 65.365 143.425 65.695 143.925 ;
        RECT 64.300 142.865 64.800 143.245 ;
        RECT 65.025 143.085 65.720 143.255 ;
        RECT 62.780 142.525 64.130 142.695 ;
        RECT 63.710 142.485 64.130 142.525 ;
        RECT 62.420 142.015 62.840 142.355 ;
        RECT 63.130 142.025 63.540 142.355 ;
        RECT 60.660 141.595 61.510 141.765 ;
        RECT 62.070 141.375 62.390 141.835 ;
        RECT 62.590 141.585 62.840 142.015 ;
        RECT 63.130 141.375 63.540 141.815 ;
        RECT 63.710 141.755 63.880 142.485 ;
        RECT 64.050 141.935 64.400 142.305 ;
        RECT 64.580 141.995 64.800 142.865 ;
        RECT 64.970 142.295 65.380 142.915 ;
        RECT 65.550 142.115 65.720 143.085 ;
        RECT 65.025 141.925 65.720 142.115 ;
        RECT 63.710 141.555 64.725 141.755 ;
        RECT 65.025 141.595 65.195 141.925 ;
        RECT 65.365 141.375 65.695 141.755 ;
        RECT 65.910 141.635 66.135 143.755 ;
        RECT 66.305 143.425 66.635 143.925 ;
        RECT 66.805 143.255 66.975 143.755 ;
        RECT 66.310 143.085 66.975 143.255 ;
        RECT 66.310 142.095 66.540 143.085 ;
        RECT 66.710 142.265 67.060 142.915 ;
        RECT 67.235 142.760 67.525 143.925 ;
        RECT 67.870 142.785 68.200 143.925 ;
        RECT 68.500 142.705 68.840 143.645 ;
        RECT 67.750 142.365 68.330 142.615 ;
        RECT 68.500 142.365 68.830 142.705 ;
        RECT 69.010 142.535 69.330 143.645 ;
        RECT 69.000 142.365 69.330 142.535 ;
        RECT 69.510 142.535 69.815 143.645 ;
        RECT 69.985 142.775 70.315 143.755 ;
        RECT 69.510 142.365 69.840 142.535 ;
        RECT 70.050 142.195 70.220 142.775 ;
        RECT 70.485 142.735 70.745 143.925 ;
        RECT 71.835 142.785 72.095 143.925 ;
        RECT 72.335 143.415 73.950 143.745 ;
        RECT 72.345 142.615 72.515 143.175 ;
        RECT 72.775 143.075 73.950 143.245 ;
        RECT 74.120 143.125 74.400 143.925 ;
        RECT 72.775 142.785 73.105 143.075 ;
        RECT 73.780 142.955 73.950 143.075 ;
        RECT 73.275 142.615 73.520 142.905 ;
        RECT 73.780 142.785 74.440 142.955 ;
        RECT 74.610 142.785 74.885 143.755 ;
        RECT 74.270 142.615 74.440 142.785 ;
        RECT 70.390 142.365 70.725 142.565 ;
        RECT 71.840 142.365 72.175 142.615 ;
        RECT 72.345 142.285 73.060 142.615 ;
        RECT 73.275 142.285 74.100 142.615 ;
        RECT 74.270 142.285 74.545 142.615 ;
        RECT 72.345 142.195 72.595 142.285 ;
        RECT 66.310 141.925 66.975 142.095 ;
        RECT 66.305 141.375 66.635 141.755 ;
        RECT 66.805 141.635 66.975 141.925 ;
        RECT 67.235 141.375 67.525 142.100 ;
        RECT 67.870 142.025 69.880 142.195 ;
        RECT 70.050 142.025 70.745 142.195 ;
        RECT 67.870 141.545 68.200 142.025 ;
        RECT 68.370 141.375 68.620 141.855 ;
        RECT 68.790 141.545 69.120 142.025 ;
        RECT 69.710 141.855 69.880 142.025 ;
        RECT 69.290 141.375 69.540 141.855 ;
        RECT 69.710 141.545 70.040 141.855 ;
        RECT 70.405 141.545 70.745 142.025 ;
        RECT 71.835 141.375 72.095 142.195 ;
        RECT 72.265 141.775 72.595 142.195 ;
        RECT 74.270 142.115 74.440 142.285 ;
        RECT 72.775 141.945 74.440 142.115 ;
        RECT 74.715 142.050 74.885 142.785 ;
        RECT 72.775 141.545 73.035 141.945 ;
        RECT 73.205 141.375 73.535 141.775 ;
        RECT 73.705 141.595 73.875 141.945 ;
        RECT 74.045 141.375 74.420 141.775 ;
        RECT 74.610 141.705 74.885 142.050 ;
        RECT 75.980 143.295 76.315 143.755 ;
        RECT 76.485 143.465 76.705 143.925 ;
        RECT 77.235 143.545 78.545 143.715 ;
        RECT 78.375 143.295 78.545 143.545 ;
        RECT 78.715 143.465 79.005 143.925 ;
        RECT 75.980 143.125 78.205 143.295 ;
        RECT 78.375 143.125 79.035 143.295 ;
        RECT 75.980 141.545 76.310 143.125 ;
        RECT 78.035 142.955 78.205 143.125 ;
        RECT 76.480 142.045 76.670 142.915 ;
        RECT 76.940 142.605 77.755 142.915 ;
        RECT 78.035 142.785 78.695 142.955 ;
        RECT 77.585 142.570 77.755 142.605 ;
        RECT 76.940 142.025 77.405 142.315 ;
        RECT 77.585 142.055 78.215 142.570 ;
        RECT 78.525 142.285 78.695 142.785 ;
        RECT 78.865 142.615 79.035 143.125 ;
        RECT 79.205 142.885 79.515 143.755 ;
        RECT 78.865 142.285 79.175 142.615 ;
        RECT 78.865 142.095 79.035 142.285 ;
        RECT 76.480 141.375 76.680 141.875 ;
        RECT 76.940 141.710 77.130 142.025 ;
        RECT 78.425 141.925 79.035 142.095 ;
        RECT 79.345 142.040 79.515 142.885 ;
        RECT 79.685 142.785 79.940 143.925 ;
        RECT 80.115 142.835 81.325 143.925 ;
        RECT 78.425 141.755 78.595 141.925 ;
        RECT 77.300 141.585 78.595 141.755 ;
        RECT 78.765 141.375 79.095 141.755 ;
        RECT 79.265 141.545 79.515 142.040 ;
        RECT 79.685 141.375 79.940 142.175 ;
        RECT 80.115 142.125 80.635 142.665 ;
        RECT 80.805 142.295 81.325 142.835 ;
        RECT 81.500 142.785 81.755 143.925 ;
        RECT 81.950 143.375 83.145 143.705 ;
        RECT 82.005 142.615 82.175 143.175 ;
        RECT 82.400 142.955 82.820 143.205 ;
        RECT 83.325 143.125 83.605 143.925 ;
        RECT 82.400 142.785 83.645 142.955 ;
        RECT 83.815 142.785 84.085 143.755 ;
        RECT 84.255 142.835 86.845 143.925 ;
        RECT 87.120 143.125 87.375 143.925 ;
        RECT 87.545 142.955 87.875 143.755 ;
        RECT 88.045 143.125 88.215 143.925 ;
        RECT 88.385 142.955 88.715 143.755 ;
        RECT 83.475 142.615 83.645 142.785 ;
        RECT 81.500 142.365 81.835 142.615 ;
        RECT 82.005 142.285 82.745 142.615 ;
        RECT 83.475 142.285 83.705 142.615 ;
        RECT 82.005 142.195 82.255 142.285 ;
        RECT 80.115 141.375 81.325 142.125 ;
        RECT 81.520 142.025 82.255 142.195 ;
        RECT 83.475 142.115 83.645 142.285 ;
        RECT 81.520 141.555 81.830 142.025 ;
        RECT 82.905 141.945 83.645 142.115 ;
        RECT 83.915 142.050 84.085 142.785 ;
        RECT 82.000 141.375 82.735 141.855 ;
        RECT 82.905 141.595 83.075 141.945 ;
        RECT 83.245 141.375 83.625 141.775 ;
        RECT 83.815 141.705 84.085 142.050 ;
        RECT 84.255 142.145 85.465 142.665 ;
        RECT 85.635 142.315 86.845 142.835 ;
        RECT 87.015 142.785 88.715 142.955 ;
        RECT 88.885 142.785 89.145 143.925 ;
        RECT 89.315 143.075 89.575 143.755 ;
        RECT 89.745 143.145 89.995 143.925 ;
        RECT 90.245 143.375 90.495 143.755 ;
        RECT 90.665 143.545 91.020 143.925 ;
        RECT 92.025 143.535 92.360 143.755 ;
        RECT 91.625 143.375 91.855 143.415 ;
        RECT 90.245 143.175 91.855 143.375 ;
        RECT 90.245 143.165 91.080 143.175 ;
        RECT 91.670 143.085 91.855 143.175 ;
        RECT 87.015 142.195 87.295 142.785 ;
        RECT 87.465 142.365 88.215 142.615 ;
        RECT 88.385 142.365 89.145 142.615 ;
        RECT 84.255 141.375 86.845 142.145 ;
        RECT 87.015 141.945 87.875 142.195 ;
        RECT 88.045 142.005 89.145 142.175 ;
        RECT 87.125 141.755 87.455 141.775 ;
        RECT 88.045 141.755 88.295 142.005 ;
        RECT 87.125 141.545 88.295 141.755 ;
        RECT 88.465 141.375 88.635 141.835 ;
        RECT 88.805 141.545 89.145 142.005 ;
        RECT 89.315 141.875 89.485 143.075 ;
        RECT 91.185 142.975 91.515 143.005 ;
        RECT 89.715 142.915 91.515 142.975 ;
        RECT 92.105 142.915 92.360 143.535 ;
        RECT 89.655 142.805 92.360 142.915 ;
        RECT 89.655 142.770 89.855 142.805 ;
        RECT 89.655 142.195 89.825 142.770 ;
        RECT 91.185 142.745 92.360 142.805 ;
        RECT 92.995 142.760 93.285 143.925 ;
        RECT 93.455 142.835 96.965 143.925 ;
        RECT 90.055 142.330 90.465 142.635 ;
        RECT 90.635 142.365 90.965 142.575 ;
        RECT 89.655 142.075 89.925 142.195 ;
        RECT 89.655 142.030 90.500 142.075 ;
        RECT 89.745 141.905 90.500 142.030 ;
        RECT 90.755 141.965 90.965 142.365 ;
        RECT 91.210 142.365 91.685 142.575 ;
        RECT 91.875 142.365 92.365 142.565 ;
        RECT 91.210 141.965 91.430 142.365 ;
        RECT 93.455 142.145 95.105 142.665 ;
        RECT 95.275 142.315 96.965 142.835 ;
        RECT 98.055 142.320 98.335 143.755 ;
        RECT 98.505 143.150 99.215 143.925 ;
        RECT 99.385 142.980 99.715 143.755 ;
        RECT 98.565 142.765 99.715 142.980 ;
        RECT 89.315 141.545 89.575 141.875 ;
        RECT 90.330 141.755 90.500 141.905 ;
        RECT 89.745 141.375 90.075 141.735 ;
        RECT 90.330 141.545 91.630 141.755 ;
        RECT 91.905 141.375 92.360 142.140 ;
        RECT 92.995 141.375 93.285 142.100 ;
        RECT 93.455 141.375 96.965 142.145 ;
        RECT 98.055 141.545 98.395 142.320 ;
        RECT 98.565 142.195 98.850 142.765 ;
        RECT 99.035 142.365 99.505 142.595 ;
        RECT 99.910 142.565 100.125 143.680 ;
        RECT 100.305 143.205 100.635 143.925 ;
        RECT 100.415 142.565 100.645 142.905 ;
        RECT 100.815 142.785 101.095 143.925 ;
        RECT 101.265 142.775 101.595 143.755 ;
        RECT 101.765 142.785 102.025 143.925 ;
        RECT 102.855 143.085 103.105 143.925 ;
        RECT 103.275 142.915 103.525 143.755 ;
        RECT 103.695 143.085 103.945 143.925 ;
        RECT 104.115 142.915 104.365 143.755 ;
        RECT 104.575 143.125 105.275 143.925 ;
        RECT 105.445 143.585 106.625 143.755 ;
        RECT 105.445 142.955 105.710 143.585 ;
        RECT 99.675 142.385 100.125 142.565 ;
        RECT 99.675 142.365 100.005 142.385 ;
        RECT 100.315 142.365 100.645 142.565 ;
        RECT 100.825 142.345 101.160 142.615 ;
        RECT 101.330 142.225 101.500 142.775 ;
        RECT 102.655 142.745 104.365 142.915 ;
        RECT 104.620 142.785 105.710 142.955 ;
        RECT 101.670 142.365 102.005 142.615 ;
        RECT 98.565 142.005 99.275 142.195 ;
        RECT 98.975 141.865 99.275 142.005 ;
        RECT 99.465 142.005 100.645 142.195 ;
        RECT 101.330 142.175 101.505 142.225 ;
        RECT 102.655 142.195 102.945 142.745 ;
        RECT 104.620 142.535 104.840 142.785 ;
        RECT 105.880 142.615 106.115 143.340 ;
        RECT 106.285 142.785 106.625 143.585 ;
        RECT 106.820 142.915 107.115 143.755 ;
        RECT 107.285 143.085 107.535 143.925 ;
        RECT 107.705 143.255 107.955 143.755 ;
        RECT 108.125 143.425 108.375 143.925 ;
        RECT 108.545 143.255 108.795 143.755 ;
        RECT 108.965 143.425 109.215 143.925 ;
        RECT 109.485 143.585 113.095 143.755 ;
        RECT 109.485 143.425 109.735 143.585 ;
        RECT 110.325 143.425 110.575 143.585 ;
        RECT 109.905 143.255 110.155 143.415 ;
        RECT 110.745 143.255 110.995 143.415 ;
        RECT 107.705 143.085 110.995 143.255 ;
        RECT 111.165 143.085 111.415 143.585 ;
        RECT 111.585 142.915 111.835 143.415 ;
        RECT 112.005 143.085 112.255 143.585 ;
        RECT 112.425 142.915 112.675 143.415 ;
        RECT 112.845 143.085 113.095 143.585 ;
        RECT 113.265 142.915 113.470 143.705 ;
        RECT 106.820 142.745 111.415 142.915 ;
        RECT 111.585 142.745 113.470 142.915 ;
        RECT 103.115 142.365 104.840 142.535 ;
        RECT 105.010 142.365 105.485 142.615 ;
        RECT 105.655 142.365 106.115 142.615 ;
        RECT 106.285 142.365 106.625 142.615 ;
        RECT 106.820 142.365 107.155 142.575 ;
        RECT 104.620 142.195 104.840 142.365 ;
        RECT 107.325 142.195 107.495 142.745 ;
        RECT 111.245 142.575 111.415 142.745 ;
        RECT 107.745 142.365 109.400 142.575 ;
        RECT 109.745 142.365 111.010 142.575 ;
        RECT 111.245 142.365 112.835 142.575 ;
        RECT 113.130 142.195 113.470 142.745 ;
        RECT 99.465 141.925 99.795 142.005 ;
        RECT 98.975 141.855 99.290 141.865 ;
        RECT 98.975 141.845 99.300 141.855 ;
        RECT 98.975 141.840 99.310 141.845 ;
        RECT 98.565 141.375 98.735 141.835 ;
        RECT 98.975 141.830 99.315 141.840 ;
        RECT 98.975 141.825 99.320 141.830 ;
        RECT 98.975 141.815 99.325 141.825 ;
        RECT 98.975 141.810 99.330 141.815 ;
        RECT 98.975 141.545 99.335 141.810 ;
        RECT 99.965 141.375 100.135 141.835 ;
        RECT 100.305 141.545 100.645 142.005 ;
        RECT 100.815 141.375 101.125 142.175 ;
        RECT 101.330 141.545 102.025 142.175 ;
        RECT 102.655 142.025 104.405 142.195 ;
        RECT 102.895 141.375 103.065 141.845 ;
        RECT 103.235 141.555 103.565 142.025 ;
        RECT 103.735 141.375 103.905 141.845 ;
        RECT 104.075 141.555 104.405 142.025 ;
        RECT 104.620 142.015 106.625 142.195 ;
        RECT 104.575 141.375 105.275 141.845 ;
        RECT 105.445 141.545 105.775 142.015 ;
        RECT 105.945 141.375 106.115 141.845 ;
        RECT 106.285 141.545 106.625 142.015 ;
        RECT 106.820 142.025 107.495 142.195 ;
        RECT 106.820 141.545 107.155 142.025 ;
        RECT 107.665 142.015 113.470 142.195 ;
        RECT 107.325 141.375 107.495 141.845 ;
        RECT 107.665 141.545 107.995 142.015 ;
        RECT 108.165 141.375 108.335 141.845 ;
        RECT 108.505 141.545 108.835 142.015 ;
        RECT 109.005 141.375 109.695 141.845 ;
        RECT 109.865 141.545 110.195 142.015 ;
        RECT 110.365 141.375 110.535 141.845 ;
        RECT 110.705 141.545 111.035 142.015 ;
        RECT 111.205 141.375 111.375 141.845 ;
        RECT 111.545 141.545 111.875 142.015 ;
        RECT 112.045 141.375 112.215 141.845 ;
        RECT 112.385 141.545 112.715 142.015 ;
        RECT 112.885 141.375 113.055 141.845 ;
        RECT 113.225 141.605 113.470 142.015 ;
        RECT 113.700 143.295 114.035 143.755 ;
        RECT 114.205 143.465 114.425 143.925 ;
        RECT 114.955 143.545 116.265 143.715 ;
        RECT 116.095 143.295 116.265 143.545 ;
        RECT 116.435 143.465 116.725 143.925 ;
        RECT 113.700 143.125 115.925 143.295 ;
        RECT 116.095 143.125 116.755 143.295 ;
        RECT 113.700 141.545 114.030 143.125 ;
        RECT 115.755 142.955 115.925 143.125 ;
        RECT 114.200 142.045 114.390 142.915 ;
        RECT 114.660 142.605 115.475 142.915 ;
        RECT 115.755 142.785 116.415 142.955 ;
        RECT 115.305 142.570 115.475 142.605 ;
        RECT 114.660 142.025 115.125 142.315 ;
        RECT 115.305 142.055 115.935 142.570 ;
        RECT 116.245 142.285 116.415 142.785 ;
        RECT 116.585 142.615 116.755 143.125 ;
        RECT 116.925 142.885 117.235 143.755 ;
        RECT 116.585 142.285 116.895 142.615 ;
        RECT 116.585 142.095 116.755 142.285 ;
        RECT 114.200 141.375 114.400 141.875 ;
        RECT 114.660 141.710 114.850 142.025 ;
        RECT 116.145 141.925 116.755 142.095 ;
        RECT 117.065 142.040 117.235 142.885 ;
        RECT 117.405 142.785 117.660 143.925 ;
        RECT 118.755 142.760 119.045 143.925 ;
        RECT 119.235 143.085 119.490 143.755 ;
        RECT 119.660 143.165 119.990 143.925 ;
        RECT 120.160 143.325 120.410 143.755 ;
        RECT 120.580 143.505 120.935 143.925 ;
        RECT 121.125 143.585 122.295 143.755 ;
        RECT 121.125 143.545 121.455 143.585 ;
        RECT 121.565 143.325 121.795 143.415 ;
        RECT 120.160 143.085 121.795 143.325 ;
        RECT 121.965 143.085 122.295 143.585 ;
        RECT 116.145 141.755 116.315 141.925 ;
        RECT 115.020 141.585 116.315 141.755 ;
        RECT 116.485 141.375 116.815 141.755 ;
        RECT 116.985 141.545 117.235 142.040 ;
        RECT 117.405 141.375 117.660 142.175 ;
        RECT 118.755 141.375 119.045 142.100 ;
        RECT 119.235 141.955 119.405 143.085 ;
        RECT 122.465 142.915 122.635 143.755 ;
        RECT 119.575 142.745 122.635 142.915 ;
        RECT 122.895 142.785 123.235 143.755 ;
        RECT 123.405 142.785 123.575 143.925 ;
        RECT 123.845 143.125 124.095 143.925 ;
        RECT 124.740 142.955 125.070 143.755 ;
        RECT 125.370 143.125 125.700 143.925 ;
        RECT 125.870 142.955 126.200 143.755 ;
        RECT 123.765 142.785 126.200 142.955 ;
        RECT 126.585 142.865 126.915 143.715 ;
        RECT 119.575 142.195 119.745 142.745 ;
        RECT 122.895 142.735 123.125 142.785 ;
        RECT 119.975 142.365 120.340 142.565 ;
        RECT 120.510 142.365 120.840 142.565 ;
        RECT 119.575 142.025 120.375 142.195 ;
        RECT 119.235 141.885 119.420 141.955 ;
        RECT 119.235 141.875 119.445 141.885 ;
        RECT 119.235 141.545 119.490 141.875 ;
        RECT 119.705 141.375 120.035 141.855 ;
        RECT 120.205 141.795 120.375 142.025 ;
        RECT 120.555 141.965 120.840 142.365 ;
        RECT 121.110 142.365 121.585 142.565 ;
        RECT 121.755 142.365 122.200 142.565 ;
        RECT 122.370 142.365 122.720 142.575 ;
        RECT 121.110 141.965 121.390 142.365 ;
        RECT 121.570 142.025 122.635 142.195 ;
        RECT 121.570 141.795 121.740 142.025 ;
        RECT 120.205 141.545 121.740 141.795 ;
        RECT 121.965 141.375 122.295 141.855 ;
        RECT 122.465 141.545 122.635 142.025 ;
        RECT 122.895 142.175 123.070 142.735 ;
        RECT 123.765 142.535 123.935 142.785 ;
        RECT 123.240 142.365 123.935 142.535 ;
        RECT 124.110 142.365 124.530 142.565 ;
        RECT 124.700 142.365 125.030 142.565 ;
        RECT 125.200 142.365 125.530 142.565 ;
        RECT 122.895 141.545 123.235 142.175 ;
        RECT 123.405 141.375 123.655 142.175 ;
        RECT 123.845 142.025 125.070 142.195 ;
        RECT 123.845 141.545 124.175 142.025 ;
        RECT 124.345 141.375 124.570 141.835 ;
        RECT 124.740 141.545 125.070 142.025 ;
        RECT 125.700 142.155 125.870 142.785 ;
        RECT 126.055 142.365 126.405 142.615 ;
        RECT 125.700 141.545 126.200 142.155 ;
        RECT 126.585 142.100 126.775 142.865 ;
        RECT 127.085 142.785 127.335 143.925 ;
        RECT 127.525 143.285 127.775 143.705 ;
        RECT 128.005 143.455 128.335 143.925 ;
        RECT 128.565 143.285 128.815 143.705 ;
        RECT 127.525 143.115 128.815 143.285 ;
        RECT 128.995 143.285 129.325 143.715 ;
        RECT 128.995 143.115 129.450 143.285 ;
        RECT 127.515 142.615 127.730 142.945 ;
        RECT 126.945 142.285 127.255 142.615 ;
        RECT 127.425 142.285 127.730 142.615 ;
        RECT 127.905 142.285 128.190 142.945 ;
        RECT 128.385 142.285 128.650 142.945 ;
        RECT 128.865 142.285 129.110 142.945 ;
        RECT 127.085 142.115 127.255 142.285 ;
        RECT 129.280 142.115 129.450 143.115 ;
        RECT 126.585 141.590 126.915 142.100 ;
        RECT 127.085 141.945 129.450 142.115 ;
        RECT 127.085 141.375 127.415 141.775 ;
        RECT 128.465 141.605 128.795 141.945 ;
        RECT 128.965 141.375 129.295 141.775 ;
        RECT 129.805 141.555 130.065 143.745 ;
        RECT 130.235 143.195 130.575 143.925 ;
        RECT 130.755 143.015 131.025 143.745 ;
        RECT 130.255 142.795 131.025 143.015 ;
        RECT 131.205 143.035 131.435 143.745 ;
        RECT 131.605 143.215 131.935 143.925 ;
        RECT 132.105 143.035 132.365 143.745 ;
        RECT 131.205 142.795 132.365 143.035 ;
        RECT 133.500 142.915 133.795 143.755 ;
        RECT 133.965 143.085 134.215 143.925 ;
        RECT 134.385 143.255 134.635 143.755 ;
        RECT 134.805 143.425 135.055 143.925 ;
        RECT 135.225 143.255 135.475 143.755 ;
        RECT 135.645 143.425 135.895 143.925 ;
        RECT 136.165 143.585 139.775 143.755 ;
        RECT 136.165 143.425 136.415 143.585 ;
        RECT 137.005 143.425 137.255 143.585 ;
        RECT 136.585 143.255 136.835 143.415 ;
        RECT 137.425 143.255 137.675 143.415 ;
        RECT 134.385 143.085 137.675 143.255 ;
        RECT 137.845 143.085 138.095 143.585 ;
        RECT 138.265 142.915 138.515 143.415 ;
        RECT 138.685 143.085 138.935 143.585 ;
        RECT 139.105 142.915 139.355 143.415 ;
        RECT 139.525 143.085 139.775 143.585 ;
        RECT 139.945 142.915 140.150 143.705 ;
        RECT 130.255 142.125 130.545 142.795 ;
        RECT 133.500 142.745 138.095 142.915 ;
        RECT 138.265 142.745 140.150 142.915 ;
        RECT 140.385 142.945 140.715 143.755 ;
        RECT 140.885 143.125 141.125 143.925 ;
        RECT 140.385 142.775 141.100 142.945 ;
        RECT 130.725 142.305 131.190 142.615 ;
        RECT 131.370 142.305 131.895 142.615 ;
        RECT 130.255 141.925 131.485 142.125 ;
        RECT 130.325 141.375 130.995 141.745 ;
        RECT 131.175 141.555 131.485 141.925 ;
        RECT 131.665 141.665 131.895 142.305 ;
        RECT 132.075 142.285 132.375 142.615 ;
        RECT 133.500 142.365 133.835 142.575 ;
        RECT 134.005 142.195 134.175 142.745 ;
        RECT 137.925 142.575 138.095 142.745 ;
        RECT 134.425 142.365 136.080 142.575 ;
        RECT 136.425 142.365 137.690 142.575 ;
        RECT 137.925 142.365 139.515 142.575 ;
        RECT 139.810 142.195 140.150 142.745 ;
        RECT 140.380 142.365 140.760 142.605 ;
        RECT 140.930 142.535 141.100 142.775 ;
        RECT 141.305 142.905 141.475 143.755 ;
        RECT 141.645 143.125 141.975 143.925 ;
        RECT 142.145 142.905 142.315 143.755 ;
        RECT 141.305 142.735 142.315 142.905 ;
        RECT 142.485 142.775 142.815 143.925 ;
        RECT 143.145 142.955 143.475 143.740 ;
        RECT 143.145 142.785 143.825 142.955 ;
        RECT 144.005 142.785 144.335 143.925 ;
        RECT 140.930 142.365 141.430 142.535 ;
        RECT 140.930 142.195 141.100 142.365 ;
        RECT 141.820 142.225 142.315 142.735 ;
        RECT 143.135 142.365 143.485 142.615 ;
        RECT 141.815 142.195 142.315 142.225 ;
        RECT 132.075 141.375 132.365 142.105 ;
        RECT 133.500 142.025 134.175 142.195 ;
        RECT 133.500 141.545 133.835 142.025 ;
        RECT 134.345 142.015 140.150 142.195 ;
        RECT 134.005 141.375 134.175 141.845 ;
        RECT 134.345 141.545 134.675 142.015 ;
        RECT 134.845 141.375 135.015 141.845 ;
        RECT 135.185 141.545 135.515 142.015 ;
        RECT 135.685 141.375 136.375 141.845 ;
        RECT 136.545 141.545 136.875 142.015 ;
        RECT 137.045 141.375 137.215 141.845 ;
        RECT 137.385 141.545 137.715 142.015 ;
        RECT 137.885 141.375 138.055 141.845 ;
        RECT 138.225 141.545 138.555 142.015 ;
        RECT 138.725 141.375 138.895 141.845 ;
        RECT 139.065 141.545 139.395 142.015 ;
        RECT 139.565 141.375 139.735 141.845 ;
        RECT 139.905 141.605 140.150 142.015 ;
        RECT 140.465 142.025 141.100 142.195 ;
        RECT 141.305 142.025 142.315 142.195 ;
        RECT 143.655 142.185 143.825 142.785 ;
        RECT 144.515 142.760 144.805 143.925 ;
        RECT 145.030 143.055 145.315 143.925 ;
        RECT 145.485 143.295 145.745 143.755 ;
        RECT 145.920 143.465 146.175 143.925 ;
        RECT 146.345 143.295 146.605 143.755 ;
        RECT 145.485 143.125 146.605 143.295 ;
        RECT 146.775 143.125 147.085 143.925 ;
        RECT 145.485 142.875 145.745 143.125 ;
        RECT 147.255 142.955 147.565 143.755 ;
        RECT 147.735 143.490 153.080 143.925 ;
        RECT 144.990 142.705 145.745 142.875 ;
        RECT 146.535 142.785 147.565 142.955 ;
        RECT 143.995 142.365 144.345 142.615 ;
        RECT 144.990 142.195 145.395 142.705 ;
        RECT 146.535 142.535 146.705 142.785 ;
        RECT 145.565 142.365 146.705 142.535 ;
        RECT 140.465 141.545 140.635 142.025 ;
        RECT 140.815 141.375 141.055 141.855 ;
        RECT 141.305 141.545 141.475 142.025 ;
        RECT 141.645 141.375 141.975 141.855 ;
        RECT 142.145 141.545 142.315 142.025 ;
        RECT 142.485 141.375 142.815 142.175 ;
        RECT 143.155 141.375 143.395 142.185 ;
        RECT 143.565 141.545 143.895 142.185 ;
        RECT 144.065 141.375 144.335 142.185 ;
        RECT 144.515 141.375 144.805 142.100 ;
        RECT 144.990 142.025 146.640 142.195 ;
        RECT 146.875 142.045 147.225 142.615 ;
        RECT 145.035 141.375 145.315 141.855 ;
        RECT 145.485 141.635 145.745 142.025 ;
        RECT 145.920 141.375 146.175 141.855 ;
        RECT 146.345 141.635 146.640 142.025 ;
        RECT 147.395 141.875 147.565 142.785 ;
        RECT 149.320 141.920 149.660 142.750 ;
        RECT 151.140 142.240 151.490 143.490 ;
        RECT 153.255 142.835 156.765 143.925 ;
        RECT 153.255 142.145 154.905 142.665 ;
        RECT 155.075 142.315 156.765 142.835 ;
        RECT 156.935 142.835 158.145 143.925 ;
        RECT 156.935 142.295 157.455 142.835 ;
        RECT 146.820 141.375 147.095 141.855 ;
        RECT 147.265 141.545 147.565 141.875 ;
        RECT 147.735 141.375 153.080 141.920 ;
        RECT 153.255 141.375 156.765 142.145 ;
        RECT 157.625 142.125 158.145 142.665 ;
        RECT 156.935 141.375 158.145 142.125 ;
        RECT 2.750 141.205 158.230 141.375 ;
        RECT 2.835 140.455 4.045 141.205 ;
        RECT 2.835 139.915 3.355 140.455 ;
        RECT 4.680 140.440 5.135 141.205 ;
        RECT 5.410 140.825 6.710 141.035 ;
        RECT 6.965 140.845 7.295 141.205 ;
        RECT 6.540 140.675 6.710 140.825 ;
        RECT 7.465 140.705 7.725 141.035 ;
        RECT 7.495 140.695 7.725 140.705 ;
        RECT 3.525 139.745 4.045 140.285 ;
        RECT 5.610 140.215 5.830 140.615 ;
        RECT 4.675 140.015 5.165 140.215 ;
        RECT 5.355 140.005 5.830 140.215 ;
        RECT 6.075 140.215 6.285 140.615 ;
        RECT 6.540 140.550 7.295 140.675 ;
        RECT 6.540 140.505 7.385 140.550 ;
        RECT 7.115 140.385 7.385 140.505 ;
        RECT 6.075 140.005 6.405 140.215 ;
        RECT 6.575 139.945 6.985 140.250 ;
        RECT 2.835 138.655 4.045 139.745 ;
        RECT 4.680 139.775 5.855 139.835 ;
        RECT 7.215 139.810 7.385 140.385 ;
        RECT 7.185 139.775 7.385 139.810 ;
        RECT 4.680 139.665 7.385 139.775 ;
        RECT 4.680 139.045 4.935 139.665 ;
        RECT 5.525 139.605 7.325 139.665 ;
        RECT 5.525 139.575 5.855 139.605 ;
        RECT 7.555 139.505 7.725 140.695 ;
        RECT 5.185 139.405 5.370 139.495 ;
        RECT 5.960 139.405 6.795 139.415 ;
        RECT 5.185 139.205 6.795 139.405 ;
        RECT 5.185 139.165 5.415 139.205 ;
        RECT 4.680 138.825 5.015 139.045 ;
        RECT 6.020 138.655 6.375 139.035 ;
        RECT 6.545 138.825 6.795 139.205 ;
        RECT 7.045 138.655 7.295 139.435 ;
        RECT 7.465 138.825 7.725 139.505 ;
        RECT 7.895 140.705 8.155 141.035 ;
        RECT 8.325 140.845 8.655 141.205 ;
        RECT 8.910 140.825 10.210 141.035 ;
        RECT 7.895 139.505 8.065 140.705 ;
        RECT 8.910 140.675 9.080 140.825 ;
        RECT 8.325 140.550 9.080 140.675 ;
        RECT 8.235 140.505 9.080 140.550 ;
        RECT 8.235 140.385 8.505 140.505 ;
        RECT 8.235 139.810 8.405 140.385 ;
        RECT 8.635 139.945 9.045 140.250 ;
        RECT 9.335 140.215 9.545 140.615 ;
        RECT 9.215 140.005 9.545 140.215 ;
        RECT 9.790 140.215 10.010 140.615 ;
        RECT 10.485 140.440 10.940 141.205 ;
        RECT 11.205 140.655 11.375 140.945 ;
        RECT 11.545 140.825 11.875 141.205 ;
        RECT 11.205 140.485 11.870 140.655 ;
        RECT 9.790 140.005 10.265 140.215 ;
        RECT 10.455 140.015 10.945 140.215 ;
        RECT 8.235 139.775 8.435 139.810 ;
        RECT 9.765 139.775 10.940 139.835 ;
        RECT 8.235 139.665 10.940 139.775 ;
        RECT 11.120 139.665 11.470 140.315 ;
        RECT 8.295 139.605 10.095 139.665 ;
        RECT 9.765 139.575 10.095 139.605 ;
        RECT 7.895 138.825 8.155 139.505 ;
        RECT 8.325 138.655 8.575 139.435 ;
        RECT 8.825 139.405 9.660 139.415 ;
        RECT 10.250 139.405 10.435 139.495 ;
        RECT 8.825 139.205 10.435 139.405 ;
        RECT 8.825 138.825 9.075 139.205 ;
        RECT 10.205 139.165 10.435 139.205 ;
        RECT 10.685 139.045 10.940 139.665 ;
        RECT 11.640 139.495 11.870 140.485 ;
        RECT 9.245 138.655 9.600 139.035 ;
        RECT 10.605 138.825 10.940 139.045 ;
        RECT 11.205 139.325 11.870 139.495 ;
        RECT 11.205 138.825 11.375 139.325 ;
        RECT 11.545 138.655 11.875 139.155 ;
        RECT 12.045 138.825 12.270 140.945 ;
        RECT 12.485 140.825 12.815 141.205 ;
        RECT 12.985 140.655 13.155 140.985 ;
        RECT 13.455 140.825 14.470 141.025 ;
        RECT 12.460 140.465 13.155 140.655 ;
        RECT 12.460 139.495 12.630 140.465 ;
        RECT 12.800 139.665 13.210 140.285 ;
        RECT 13.380 139.715 13.600 140.585 ;
        RECT 13.780 140.275 14.130 140.645 ;
        RECT 14.300 140.095 14.470 140.825 ;
        RECT 14.640 140.765 15.050 141.205 ;
        RECT 15.340 140.565 15.590 140.995 ;
        RECT 15.790 140.745 16.110 141.205 ;
        RECT 16.670 140.815 17.520 140.985 ;
        RECT 14.640 140.225 15.050 140.555 ;
        RECT 15.340 140.225 15.760 140.565 ;
        RECT 14.050 140.055 14.470 140.095 ;
        RECT 14.050 139.885 15.400 140.055 ;
        RECT 12.460 139.325 13.155 139.495 ;
        RECT 13.380 139.335 13.880 139.715 ;
        RECT 12.485 138.655 12.815 139.155 ;
        RECT 12.985 138.825 13.155 139.325 ;
        RECT 14.050 139.040 14.220 139.885 ;
        RECT 15.150 139.725 15.400 139.885 ;
        RECT 14.390 139.455 14.640 139.715 ;
        RECT 15.570 139.455 15.760 140.225 ;
        RECT 14.390 139.205 15.760 139.455 ;
        RECT 15.930 140.395 17.180 140.565 ;
        RECT 15.930 139.635 16.100 140.395 ;
        RECT 16.850 140.275 17.180 140.395 ;
        RECT 16.270 139.815 16.450 140.225 ;
        RECT 17.350 140.055 17.520 140.815 ;
        RECT 17.720 140.725 18.380 141.205 ;
        RECT 18.560 140.610 18.880 140.940 ;
        RECT 17.710 140.285 18.370 140.555 ;
        RECT 17.710 140.225 18.040 140.285 ;
        RECT 18.190 140.055 18.520 140.115 ;
        RECT 16.620 139.885 18.520 140.055 ;
        RECT 15.930 139.325 16.450 139.635 ;
        RECT 16.620 139.375 16.790 139.885 ;
        RECT 18.690 139.715 18.880 140.610 ;
        RECT 16.960 139.545 18.880 139.715 ;
        RECT 18.560 139.525 18.880 139.545 ;
        RECT 19.080 140.295 19.330 140.945 ;
        RECT 19.510 140.745 19.795 141.205 ;
        RECT 19.975 140.865 20.230 141.025 ;
        RECT 19.975 140.695 20.315 140.865 ;
        RECT 19.975 140.495 20.230 140.695 ;
        RECT 19.080 139.965 19.880 140.295 ;
        RECT 16.620 139.205 17.830 139.375 ;
        RECT 13.390 138.870 14.220 139.040 ;
        RECT 14.460 138.655 14.840 139.035 ;
        RECT 15.020 138.915 15.190 139.205 ;
        RECT 16.620 139.125 16.790 139.205 ;
        RECT 15.360 138.655 15.690 139.035 ;
        RECT 16.160 138.875 16.790 139.125 ;
        RECT 16.970 138.655 17.390 139.035 ;
        RECT 17.590 138.915 17.830 139.205 ;
        RECT 18.060 138.655 18.390 139.345 ;
        RECT 18.560 138.915 18.730 139.525 ;
        RECT 19.080 139.375 19.330 139.965 ;
        RECT 20.050 139.635 20.230 140.495 ;
        RECT 19.000 138.865 19.330 139.375 ;
        RECT 19.510 138.655 19.795 139.455 ;
        RECT 19.975 138.965 20.230 139.635 ;
        RECT 20.775 140.465 21.160 141.035 ;
        RECT 21.330 140.745 21.655 141.205 ;
        RECT 22.175 140.575 22.455 141.035 ;
        RECT 20.775 139.795 21.055 140.465 ;
        RECT 21.330 140.405 22.455 140.575 ;
        RECT 21.330 140.295 21.780 140.405 ;
        RECT 21.225 139.965 21.780 140.295 ;
        RECT 22.645 140.235 23.045 141.035 ;
        RECT 23.445 140.745 23.715 141.205 ;
        RECT 23.885 140.575 24.170 141.035 ;
        RECT 20.775 138.825 21.160 139.795 ;
        RECT 21.330 139.505 21.780 139.965 ;
        RECT 21.950 139.675 23.045 140.235 ;
        RECT 21.330 139.285 22.455 139.505 ;
        RECT 21.330 138.655 21.655 139.115 ;
        RECT 22.175 138.825 22.455 139.285 ;
        RECT 22.645 138.825 23.045 139.675 ;
        RECT 23.215 140.405 24.170 140.575 ;
        RECT 24.460 140.465 24.715 141.035 ;
        RECT 24.885 140.805 25.215 141.205 ;
        RECT 25.640 140.670 26.170 141.035 ;
        RECT 25.640 140.635 25.815 140.670 ;
        RECT 24.885 140.465 25.815 140.635 ;
        RECT 23.215 139.505 23.425 140.405 ;
        RECT 23.595 139.675 24.285 140.235 ;
        RECT 24.460 139.795 24.630 140.465 ;
        RECT 24.885 140.295 25.055 140.465 ;
        RECT 24.800 139.965 25.055 140.295 ;
        RECT 25.280 139.965 25.475 140.295 ;
        RECT 23.215 139.285 24.170 139.505 ;
        RECT 23.445 138.655 23.715 139.115 ;
        RECT 23.885 138.825 24.170 139.285 ;
        RECT 24.460 138.825 24.795 139.795 ;
        RECT 24.965 138.655 25.135 139.795 ;
        RECT 25.305 138.995 25.475 139.965 ;
        RECT 25.645 139.335 25.815 140.465 ;
        RECT 25.985 139.675 26.155 140.475 ;
        RECT 26.360 140.185 26.635 141.035 ;
        RECT 26.355 140.015 26.635 140.185 ;
        RECT 26.360 139.875 26.635 140.015 ;
        RECT 26.805 139.675 26.995 141.035 ;
        RECT 27.175 140.670 27.685 141.205 ;
        RECT 27.905 140.395 28.150 141.000 ;
        RECT 28.595 140.480 28.885 141.205 ;
        RECT 29.060 140.465 29.315 141.035 ;
        RECT 29.485 140.805 29.815 141.205 ;
        RECT 30.240 140.670 30.770 141.035 ;
        RECT 30.960 140.865 31.235 141.035 ;
        RECT 30.955 140.695 31.235 140.865 ;
        RECT 30.240 140.635 30.415 140.670 ;
        RECT 29.485 140.465 30.415 140.635 ;
        RECT 27.195 140.225 28.425 140.395 ;
        RECT 25.985 139.505 26.995 139.675 ;
        RECT 27.165 139.660 27.915 139.850 ;
        RECT 25.645 139.165 26.770 139.335 ;
        RECT 27.165 138.995 27.335 139.660 ;
        RECT 28.085 139.415 28.425 140.225 ;
        RECT 25.305 138.825 27.335 138.995 ;
        RECT 27.505 138.655 27.675 139.415 ;
        RECT 27.910 139.005 28.425 139.415 ;
        RECT 28.595 138.655 28.885 139.820 ;
        RECT 29.060 139.795 29.230 140.465 ;
        RECT 29.485 140.295 29.655 140.465 ;
        RECT 29.400 139.965 29.655 140.295 ;
        RECT 29.880 139.965 30.075 140.295 ;
        RECT 29.060 138.825 29.395 139.795 ;
        RECT 29.565 138.655 29.735 139.795 ;
        RECT 29.905 138.995 30.075 139.965 ;
        RECT 30.245 139.335 30.415 140.465 ;
        RECT 30.585 139.675 30.755 140.475 ;
        RECT 30.960 139.875 31.235 140.695 ;
        RECT 31.405 139.675 31.595 141.035 ;
        RECT 31.775 140.670 32.285 141.205 ;
        RECT 32.505 140.395 32.750 141.000 ;
        RECT 33.200 140.465 33.455 141.035 ;
        RECT 33.625 140.805 33.955 141.205 ;
        RECT 34.380 140.670 34.910 141.035 ;
        RECT 34.380 140.635 34.555 140.670 ;
        RECT 33.625 140.465 34.555 140.635 ;
        RECT 31.795 140.225 33.025 140.395 ;
        RECT 30.585 139.505 31.595 139.675 ;
        RECT 31.765 139.660 32.515 139.850 ;
        RECT 30.245 139.165 31.370 139.335 ;
        RECT 31.765 138.995 31.935 139.660 ;
        RECT 32.685 139.415 33.025 140.225 ;
        RECT 29.905 138.825 31.935 138.995 ;
        RECT 32.105 138.655 32.275 139.415 ;
        RECT 32.510 139.005 33.025 139.415 ;
        RECT 33.200 139.795 33.370 140.465 ;
        RECT 33.625 140.295 33.795 140.465 ;
        RECT 33.540 139.965 33.795 140.295 ;
        RECT 34.020 139.965 34.215 140.295 ;
        RECT 33.200 138.825 33.535 139.795 ;
        RECT 33.705 138.655 33.875 139.795 ;
        RECT 34.045 138.995 34.215 139.965 ;
        RECT 34.385 139.335 34.555 140.465 ;
        RECT 34.725 139.675 34.895 140.475 ;
        RECT 35.100 140.185 35.375 141.035 ;
        RECT 35.095 140.015 35.375 140.185 ;
        RECT 35.100 139.875 35.375 140.015 ;
        RECT 35.545 139.675 35.735 141.035 ;
        RECT 35.915 140.670 36.425 141.205 ;
        RECT 36.645 140.395 36.890 141.000 ;
        RECT 37.610 140.395 37.855 141.000 ;
        RECT 38.075 140.670 38.585 141.205 ;
        RECT 35.935 140.225 37.165 140.395 ;
        RECT 34.725 139.505 35.735 139.675 ;
        RECT 35.905 139.660 36.655 139.850 ;
        RECT 34.385 139.165 35.510 139.335 ;
        RECT 35.905 138.995 36.075 139.660 ;
        RECT 36.825 139.415 37.165 140.225 ;
        RECT 34.045 138.825 36.075 138.995 ;
        RECT 36.245 138.655 36.415 139.415 ;
        RECT 36.650 139.005 37.165 139.415 ;
        RECT 37.335 140.225 38.565 140.395 ;
        RECT 37.335 139.415 37.675 140.225 ;
        RECT 37.845 139.660 38.595 139.850 ;
        RECT 37.335 139.005 37.850 139.415 ;
        RECT 38.085 138.655 38.255 139.415 ;
        RECT 38.425 138.995 38.595 139.660 ;
        RECT 38.765 139.675 38.955 141.035 ;
        RECT 39.125 140.185 39.400 141.035 ;
        RECT 39.590 140.670 40.120 141.035 ;
        RECT 40.545 140.805 40.875 141.205 ;
        RECT 39.945 140.635 40.120 140.670 ;
        RECT 39.125 140.015 39.405 140.185 ;
        RECT 39.125 139.875 39.400 140.015 ;
        RECT 39.605 139.675 39.775 140.475 ;
        RECT 38.765 139.505 39.775 139.675 ;
        RECT 39.945 140.465 40.875 140.635 ;
        RECT 41.045 140.465 41.300 141.035 ;
        RECT 41.535 140.725 41.815 141.205 ;
        RECT 41.985 140.555 42.245 140.945 ;
        RECT 42.420 140.725 42.675 141.205 ;
        RECT 42.845 140.555 43.140 140.945 ;
        RECT 43.320 140.725 43.595 141.205 ;
        RECT 43.765 140.705 44.065 141.035 ;
        RECT 39.945 139.335 40.115 140.465 ;
        RECT 40.705 140.295 40.875 140.465 ;
        RECT 38.990 139.165 40.115 139.335 ;
        RECT 40.285 139.965 40.480 140.295 ;
        RECT 40.705 139.965 40.960 140.295 ;
        RECT 40.285 138.995 40.455 139.965 ;
        RECT 41.130 139.795 41.300 140.465 ;
        RECT 38.425 138.825 40.455 138.995 ;
        RECT 40.625 138.655 40.795 139.795 ;
        RECT 40.965 138.825 41.300 139.795 ;
        RECT 41.490 140.385 43.140 140.555 ;
        RECT 41.490 139.875 41.895 140.385 ;
        RECT 42.065 140.045 43.205 140.215 ;
        RECT 41.490 139.705 42.245 139.875 ;
        RECT 41.530 138.655 41.815 139.525 ;
        RECT 41.985 139.455 42.245 139.705 ;
        RECT 43.035 139.795 43.205 140.045 ;
        RECT 43.375 139.965 43.725 140.535 ;
        RECT 43.895 139.795 44.065 140.705 ;
        RECT 43.035 139.625 44.065 139.795 ;
        RECT 41.985 139.285 43.105 139.455 ;
        RECT 41.985 138.825 42.245 139.285 ;
        RECT 42.420 138.655 42.675 139.115 ;
        RECT 42.845 138.825 43.105 139.285 ;
        RECT 43.275 138.655 43.585 139.455 ;
        RECT 43.755 138.825 44.065 139.625 ;
        RECT 44.240 140.465 44.495 141.035 ;
        RECT 44.665 140.805 44.995 141.205 ;
        RECT 45.420 140.670 45.950 141.035 ;
        RECT 46.140 140.865 46.415 141.035 ;
        RECT 46.135 140.695 46.415 140.865 ;
        RECT 45.420 140.635 45.595 140.670 ;
        RECT 44.665 140.465 45.595 140.635 ;
        RECT 44.240 139.795 44.410 140.465 ;
        RECT 44.665 140.295 44.835 140.465 ;
        RECT 44.580 139.965 44.835 140.295 ;
        RECT 45.060 139.965 45.255 140.295 ;
        RECT 44.240 138.825 44.575 139.795 ;
        RECT 44.745 138.655 44.915 139.795 ;
        RECT 45.085 138.995 45.255 139.965 ;
        RECT 45.425 139.335 45.595 140.465 ;
        RECT 45.765 139.675 45.935 140.475 ;
        RECT 46.140 139.875 46.415 140.695 ;
        RECT 46.585 139.675 46.775 141.035 ;
        RECT 46.955 140.670 47.465 141.205 ;
        RECT 47.685 140.395 47.930 141.000 ;
        RECT 48.925 140.655 49.095 141.035 ;
        RECT 49.275 140.825 49.605 141.205 ;
        RECT 48.925 140.485 49.590 140.655 ;
        RECT 49.785 140.530 50.045 141.035 ;
        RECT 46.975 140.225 48.205 140.395 ;
        RECT 45.765 139.505 46.775 139.675 ;
        RECT 46.945 139.660 47.695 139.850 ;
        RECT 45.425 139.165 46.550 139.335 ;
        RECT 46.945 138.995 47.115 139.660 ;
        RECT 47.865 139.415 48.205 140.225 ;
        RECT 48.855 139.935 49.185 140.305 ;
        RECT 49.420 140.230 49.590 140.485 ;
        RECT 49.420 139.900 49.705 140.230 ;
        RECT 49.420 139.755 49.590 139.900 ;
        RECT 45.085 138.825 47.115 138.995 ;
        RECT 47.285 138.655 47.455 139.415 ;
        RECT 47.690 139.005 48.205 139.415 ;
        RECT 48.925 139.585 49.590 139.755 ;
        RECT 49.875 139.730 50.045 140.530 ;
        RECT 50.490 140.395 50.735 141.000 ;
        RECT 50.955 140.670 51.465 141.205 ;
        RECT 48.925 138.825 49.095 139.585 ;
        RECT 49.275 138.655 49.605 139.415 ;
        RECT 49.775 138.825 50.045 139.730 ;
        RECT 50.215 140.225 51.445 140.395 ;
        RECT 50.215 139.415 50.555 140.225 ;
        RECT 50.725 139.660 51.475 139.850 ;
        RECT 50.215 139.005 50.730 139.415 ;
        RECT 50.965 138.655 51.135 139.415 ;
        RECT 51.305 138.995 51.475 139.660 ;
        RECT 51.645 139.675 51.835 141.035 ;
        RECT 52.005 140.185 52.280 141.035 ;
        RECT 52.470 140.670 53.000 141.035 ;
        RECT 53.425 140.805 53.755 141.205 ;
        RECT 52.825 140.635 53.000 140.670 ;
        RECT 52.005 140.015 52.285 140.185 ;
        RECT 52.005 139.875 52.280 140.015 ;
        RECT 52.485 139.675 52.655 140.475 ;
        RECT 51.645 139.505 52.655 139.675 ;
        RECT 52.825 140.465 53.755 140.635 ;
        RECT 53.925 140.465 54.180 141.035 ;
        RECT 54.355 140.480 54.645 141.205 ;
        RECT 54.820 140.655 55.075 140.945 ;
        RECT 55.245 140.825 55.575 141.205 ;
        RECT 54.820 140.485 55.570 140.655 ;
        RECT 52.825 139.335 52.995 140.465 ;
        RECT 53.585 140.295 53.755 140.465 ;
        RECT 51.870 139.165 52.995 139.335 ;
        RECT 53.165 139.965 53.360 140.295 ;
        RECT 53.585 139.965 53.840 140.295 ;
        RECT 53.165 138.995 53.335 139.965 ;
        RECT 54.010 139.795 54.180 140.465 ;
        RECT 51.305 138.825 53.335 138.995 ;
        RECT 53.505 138.655 53.675 139.795 ;
        RECT 53.845 138.825 54.180 139.795 ;
        RECT 54.355 138.655 54.645 139.820 ;
        RECT 54.820 139.665 55.170 140.315 ;
        RECT 55.340 139.495 55.570 140.485 ;
        RECT 54.820 139.325 55.570 139.495 ;
        RECT 54.820 138.825 55.075 139.325 ;
        RECT 55.245 138.655 55.575 139.155 ;
        RECT 55.745 138.825 55.915 140.945 ;
        RECT 56.275 140.845 56.605 141.205 ;
        RECT 56.775 140.815 57.270 140.985 ;
        RECT 57.475 140.815 58.330 140.985 ;
        RECT 56.145 139.625 56.605 140.675 ;
        RECT 56.085 138.840 56.410 139.625 ;
        RECT 56.775 139.455 56.945 140.815 ;
        RECT 57.115 139.905 57.465 140.525 ;
        RECT 57.635 140.305 57.990 140.525 ;
        RECT 57.635 139.715 57.805 140.305 ;
        RECT 58.160 140.105 58.330 140.815 ;
        RECT 59.205 140.745 59.535 141.205 ;
        RECT 59.745 140.845 60.095 141.015 ;
        RECT 58.535 140.275 59.325 140.525 ;
        RECT 59.745 140.455 60.005 140.845 ;
        RECT 60.315 140.755 61.265 141.035 ;
        RECT 61.435 140.765 61.625 141.205 ;
        RECT 61.795 140.825 62.865 140.995 ;
        RECT 59.495 140.105 59.665 140.285 ;
        RECT 56.775 139.285 57.170 139.455 ;
        RECT 57.340 139.325 57.805 139.715 ;
        RECT 57.975 139.935 59.665 140.105 ;
        RECT 57.000 139.155 57.170 139.285 ;
        RECT 57.975 139.155 58.145 139.935 ;
        RECT 59.835 139.765 60.005 140.455 ;
        RECT 58.505 139.595 60.005 139.765 ;
        RECT 60.195 139.795 60.405 140.585 ;
        RECT 60.575 139.965 60.925 140.585 ;
        RECT 61.095 139.975 61.265 140.755 ;
        RECT 61.795 140.595 61.965 140.825 ;
        RECT 61.435 140.425 61.965 140.595 ;
        RECT 61.435 140.145 61.655 140.425 ;
        RECT 62.135 140.255 62.375 140.655 ;
        RECT 61.095 139.805 61.500 139.975 ;
        RECT 61.835 139.885 62.375 140.255 ;
        RECT 62.545 140.470 62.865 140.825 ;
        RECT 63.110 140.745 63.415 141.205 ;
        RECT 63.585 140.495 63.840 141.025 ;
        RECT 62.545 140.295 62.870 140.470 ;
        RECT 62.545 139.995 63.460 140.295 ;
        RECT 62.720 139.965 63.460 139.995 ;
        RECT 60.195 139.635 60.870 139.795 ;
        RECT 61.330 139.715 61.500 139.805 ;
        RECT 60.195 139.625 61.160 139.635 ;
        RECT 59.835 139.455 60.005 139.595 ;
        RECT 56.580 138.655 56.830 139.115 ;
        RECT 57.000 138.825 57.250 139.155 ;
        RECT 57.465 138.825 58.145 139.155 ;
        RECT 58.315 139.255 59.390 139.425 ;
        RECT 59.835 139.285 60.395 139.455 ;
        RECT 60.700 139.335 61.160 139.625 ;
        RECT 61.330 139.545 62.550 139.715 ;
        RECT 58.315 138.915 58.485 139.255 ;
        RECT 58.720 138.655 59.050 139.085 ;
        RECT 59.220 138.915 59.390 139.255 ;
        RECT 59.685 138.655 60.055 139.115 ;
        RECT 60.225 138.825 60.395 139.285 ;
        RECT 61.330 139.165 61.500 139.545 ;
        RECT 62.720 139.375 62.890 139.965 ;
        RECT 63.630 139.845 63.840 140.495 ;
        RECT 60.630 138.825 61.500 139.165 ;
        RECT 62.090 139.205 62.890 139.375 ;
        RECT 61.670 138.655 61.920 139.115 ;
        RECT 62.090 138.915 62.260 139.205 ;
        RECT 62.440 138.655 62.770 139.035 ;
        RECT 63.110 138.655 63.415 139.795 ;
        RECT 63.585 138.965 63.840 139.845 ;
        RECT 64.015 140.465 64.400 141.035 ;
        RECT 64.570 140.745 64.895 141.205 ;
        RECT 65.415 140.575 65.695 141.035 ;
        RECT 64.015 139.795 64.295 140.465 ;
        RECT 64.570 140.405 65.695 140.575 ;
        RECT 64.570 140.295 65.020 140.405 ;
        RECT 64.465 139.965 65.020 140.295 ;
        RECT 65.885 140.235 66.285 141.035 ;
        RECT 66.685 140.745 66.955 141.205 ;
        RECT 67.125 140.575 67.410 141.035 ;
        RECT 68.205 140.685 68.460 140.985 ;
        RECT 68.630 140.805 68.960 141.205 ;
        RECT 64.015 138.825 64.400 139.795 ;
        RECT 64.570 139.505 65.020 139.965 ;
        RECT 65.190 139.675 66.285 140.235 ;
        RECT 64.570 139.285 65.695 139.505 ;
        RECT 64.570 138.655 64.895 139.115 ;
        RECT 65.415 138.825 65.695 139.285 ;
        RECT 65.885 138.825 66.285 139.675 ;
        RECT 66.455 140.405 67.410 140.575 ;
        RECT 68.155 140.635 68.460 140.685 ;
        RECT 69.130 140.635 69.300 140.985 ;
        RECT 69.600 140.725 69.770 141.205 ;
        RECT 70.005 140.695 70.355 141.025 ;
        RECT 70.525 140.725 70.695 141.205 ;
        RECT 68.155 140.555 69.300 140.635 ;
        RECT 68.155 140.525 69.865 140.555 ;
        RECT 68.155 140.465 70.015 140.525 ;
        RECT 66.455 139.505 66.665 140.405 ;
        RECT 66.835 139.675 67.525 140.235 ;
        RECT 68.155 139.795 68.325 140.465 ;
        RECT 69.130 140.385 70.015 140.465 ;
        RECT 69.695 140.355 70.015 140.385 ;
        RECT 68.500 139.965 68.800 140.295 ;
        RECT 66.455 139.285 67.410 139.505 ;
        RECT 68.155 139.365 68.460 139.795 ;
        RECT 68.630 139.505 68.800 139.965 ;
        RECT 69.060 139.675 69.595 140.215 ;
        RECT 69.845 139.965 70.015 140.355 ;
        RECT 70.185 139.795 70.355 140.695 ;
        RECT 70.945 140.555 71.205 141.000 ;
        RECT 71.420 140.845 71.750 141.205 ;
        RECT 71.920 140.675 72.250 141.035 ;
        RECT 72.420 140.765 72.655 141.205 ;
        RECT 73.245 140.825 73.580 141.205 ;
        RECT 74.540 140.865 74.875 141.035 ;
        RECT 69.960 139.590 70.355 139.795 ;
        RECT 70.525 140.385 71.205 140.555 ;
        RECT 71.430 140.505 72.250 140.675 ;
        RECT 68.630 139.420 69.740 139.505 ;
        RECT 70.525 139.480 70.695 140.385 ;
        RECT 70.865 139.650 71.205 140.215 ;
        RECT 70.525 139.420 71.205 139.480 ;
        RECT 68.630 139.335 71.205 139.420 ;
        RECT 66.685 138.655 66.955 139.115 ;
        RECT 67.125 138.825 67.410 139.285 ;
        RECT 69.570 139.250 71.205 139.335 ;
        RECT 68.155 138.925 69.355 139.165 ;
        RECT 69.535 138.655 69.865 139.080 ;
        RECT 70.380 138.655 70.740 139.080 ;
        RECT 70.945 139.070 71.205 139.250 ;
        RECT 71.430 139.385 71.625 140.505 ;
        RECT 72.820 140.465 74.090 140.655 ;
        RECT 74.260 140.465 74.875 140.865 ;
        RECT 75.325 140.825 77.335 141.035 ;
        RECT 71.795 139.965 72.475 140.295 ;
        RECT 72.645 139.965 72.980 140.295 ;
        RECT 73.150 140.185 73.440 140.295 ;
        RECT 73.150 140.015 73.445 140.185 ;
        RECT 73.150 139.965 73.440 140.015 ;
        RECT 73.730 139.965 74.090 140.295 ;
        RECT 72.305 139.780 72.475 139.965 ;
        RECT 74.260 139.780 74.440 140.465 ;
        RECT 75.325 140.405 75.575 140.825 ;
        RECT 75.745 140.485 76.915 140.655 ;
        RECT 74.610 139.965 74.885 140.295 ;
        RECT 76.665 140.215 76.915 140.485 ;
        RECT 77.085 140.575 77.335 140.825 ;
        RECT 77.505 140.745 77.675 141.205 ;
        RECT 77.845 140.575 78.175 141.035 ;
        RECT 78.345 140.745 78.515 141.205 ;
        RECT 78.685 140.575 79.020 141.035 ;
        RECT 77.085 140.385 79.020 140.575 ;
        RECT 80.115 140.480 80.405 141.205 ;
        RECT 80.575 140.815 81.885 140.985 ;
        RECT 75.055 139.965 76.495 140.215 ;
        RECT 76.665 139.795 77.200 140.215 ;
        RECT 77.380 139.965 79.000 140.215 ;
        RECT 80.575 139.875 80.965 140.815 ;
        RECT 82.155 140.735 82.325 141.205 ;
        RECT 81.135 140.565 81.465 140.645 ;
        RECT 82.495 140.565 82.860 141.035 ;
        RECT 83.030 140.735 83.200 141.205 ;
        RECT 83.370 140.565 83.700 141.035 ;
        RECT 81.135 140.385 83.700 140.565 ;
        RECT 83.870 140.385 84.040 141.205 ;
        RECT 84.350 140.565 84.680 141.035 ;
        RECT 84.850 140.735 85.020 141.205 ;
        RECT 85.190 140.815 86.365 141.035 ;
        RECT 85.190 140.565 85.440 140.815 ;
        RECT 84.350 140.385 85.440 140.565 ;
        RECT 85.610 140.395 86.385 140.645 ;
        RECT 81.175 140.045 81.835 140.215 ;
        RECT 72.305 139.525 74.880 139.780 ;
        RECT 71.430 139.215 72.160 139.385 ;
        RECT 71.470 138.655 71.800 139.035 ;
        RECT 71.970 138.825 72.160 139.215 ;
        RECT 72.340 138.655 72.770 139.355 ;
        RECT 73.275 138.825 73.945 139.525 ;
        RECT 74.115 138.655 74.445 139.355 ;
        RECT 74.615 138.825 74.880 139.525 ;
        RECT 75.745 139.625 78.595 139.795 ;
        RECT 75.325 138.655 75.575 139.455 ;
        RECT 75.745 138.825 76.075 139.625 ;
        RECT 76.245 138.655 76.415 139.455 ;
        RECT 76.585 138.825 76.915 139.625 ;
        RECT 77.085 138.655 77.255 139.455 ;
        RECT 77.425 138.825 77.755 139.625 ;
        RECT 77.925 138.655 78.095 139.455 ;
        RECT 78.265 138.825 78.595 139.625 ;
        RECT 78.765 138.655 79.020 139.795 ;
        RECT 80.115 138.655 80.405 139.820 ;
        RECT 80.575 139.665 81.425 139.875 ;
        RECT 81.665 139.835 81.835 140.045 ;
        RECT 82.515 140.005 83.540 140.215 ;
        RECT 83.765 140.015 85.215 140.215 ;
        RECT 83.370 139.845 83.540 140.005 ;
        RECT 85.510 140.005 85.985 140.215 ;
        RECT 85.510 139.845 85.680 140.005 ;
        RECT 81.665 139.665 83.160 139.835 ;
        RECT 83.370 139.675 85.680 139.845 ;
        RECT 81.175 139.495 81.425 139.665 ;
        RECT 82.990 139.505 83.160 139.665 ;
        RECT 86.155 139.505 86.385 140.395 ;
        RECT 86.555 140.455 87.765 141.205 ;
        RECT 86.555 139.915 87.075 140.455 ;
        RECT 87.940 140.440 88.395 141.205 ;
        RECT 88.670 140.825 89.970 141.035 ;
        RECT 90.225 140.845 90.555 141.205 ;
        RECT 89.800 140.675 89.970 140.825 ;
        RECT 90.725 140.705 90.985 141.035 ;
        RECT 90.755 140.695 90.985 140.705 ;
        RECT 87.245 139.745 87.765 140.285 ;
        RECT 88.870 140.215 89.090 140.615 ;
        RECT 87.935 140.015 88.425 140.215 ;
        RECT 88.615 140.005 89.090 140.215 ;
        RECT 89.335 140.215 89.545 140.615 ;
        RECT 89.800 140.550 90.555 140.675 ;
        RECT 89.800 140.505 90.645 140.550 ;
        RECT 90.375 140.385 90.645 140.505 ;
        RECT 89.335 140.005 89.665 140.215 ;
        RECT 89.835 139.945 90.245 140.250 ;
        RECT 80.575 138.655 81.005 139.495 ;
        RECT 81.175 139.325 82.745 139.495 ;
        RECT 82.990 139.335 86.385 139.505 ;
        RECT 81.175 139.165 81.425 139.325 ;
        RECT 82.535 139.165 82.745 139.325 ;
        RECT 84.390 139.325 86.385 139.335 ;
        RECT 81.595 138.655 81.845 139.155 ;
        RECT 82.115 138.995 82.365 139.155 ;
        RECT 82.915 138.995 83.240 139.165 ;
        RECT 82.115 138.825 83.240 138.995 ;
        RECT 83.410 138.655 83.660 139.155 ;
        RECT 83.830 138.825 84.080 139.165 ;
        RECT 84.390 138.825 84.640 139.325 ;
        RECT 84.810 138.655 85.060 139.155 ;
        RECT 85.230 138.825 85.480 139.325 ;
        RECT 85.650 138.655 85.900 139.155 ;
        RECT 86.070 138.825 86.385 139.325 ;
        RECT 86.555 138.655 87.765 139.745 ;
        RECT 87.940 139.775 89.115 139.835 ;
        RECT 90.475 139.810 90.645 140.385 ;
        RECT 90.445 139.775 90.645 139.810 ;
        RECT 87.940 139.665 90.645 139.775 ;
        RECT 87.940 139.045 88.195 139.665 ;
        RECT 88.785 139.605 90.585 139.665 ;
        RECT 88.785 139.575 89.115 139.605 ;
        RECT 90.815 139.505 90.985 140.695 ;
        RECT 91.215 140.385 91.425 141.205 ;
        RECT 91.595 140.405 91.925 141.035 ;
        RECT 91.595 139.805 91.845 140.405 ;
        RECT 92.095 140.385 92.325 141.205 ;
        RECT 92.535 140.435 96.045 141.205 ;
        RECT 97.135 140.465 97.475 141.035 ;
        RECT 97.670 140.540 97.840 141.205 ;
        RECT 98.120 140.865 98.340 140.910 ;
        RECT 98.115 140.695 98.340 140.865 ;
        RECT 98.510 140.725 98.955 140.895 ;
        RECT 98.120 140.555 98.340 140.695 ;
        RECT 92.015 139.965 92.345 140.215 ;
        RECT 92.535 139.915 94.185 140.435 ;
        RECT 88.445 139.405 88.630 139.495 ;
        RECT 89.220 139.405 90.055 139.415 ;
        RECT 88.445 139.205 90.055 139.405 ;
        RECT 88.445 139.165 88.675 139.205 ;
        RECT 87.940 138.825 88.275 139.045 ;
        RECT 89.280 138.655 89.635 139.035 ;
        RECT 89.805 138.825 90.055 139.205 ;
        RECT 90.305 138.655 90.555 139.435 ;
        RECT 90.725 138.825 90.985 139.505 ;
        RECT 91.215 138.655 91.425 139.795 ;
        RECT 91.595 138.825 91.925 139.805 ;
        RECT 92.095 138.655 92.325 139.795 ;
        RECT 94.355 139.745 96.045 140.265 ;
        RECT 92.535 138.655 96.045 139.745 ;
        RECT 97.135 139.495 97.310 140.465 ;
        RECT 98.120 140.385 98.615 140.555 ;
        RECT 97.480 139.845 97.650 140.295 ;
        RECT 97.820 140.015 98.270 140.215 ;
        RECT 98.440 140.190 98.615 140.385 ;
        RECT 98.785 139.935 98.955 140.725 ;
        RECT 99.125 140.600 99.375 140.970 ;
        RECT 99.205 140.215 99.375 140.600 ;
        RECT 99.545 140.565 99.795 140.970 ;
        RECT 99.965 140.735 100.135 141.205 ;
        RECT 100.305 140.565 100.645 140.970 ;
        RECT 99.545 140.385 100.645 140.565 ;
        RECT 100.835 140.705 101.090 141.035 ;
        RECT 101.305 140.725 101.635 141.205 ;
        RECT 101.805 140.785 103.340 141.035 ;
        RECT 100.835 140.695 101.045 140.705 ;
        RECT 100.835 140.625 101.020 140.695 ;
        RECT 99.205 140.045 99.400 140.215 ;
        RECT 97.480 139.675 97.875 139.845 ;
        RECT 98.785 139.795 99.060 139.935 ;
        RECT 97.135 138.825 97.395 139.495 ;
        RECT 97.705 139.405 97.875 139.675 ;
        RECT 98.045 139.575 99.060 139.795 ;
        RECT 99.230 139.795 99.400 140.045 ;
        RECT 99.570 139.965 100.130 140.215 ;
        RECT 99.230 139.405 99.785 139.795 ;
        RECT 97.705 139.235 99.785 139.405 ;
        RECT 97.565 138.655 97.895 139.055 ;
        RECT 98.765 138.655 99.165 139.055 ;
        RECT 99.455 139.000 99.785 139.235 ;
        RECT 99.955 138.865 100.130 139.965 ;
        RECT 100.300 139.645 100.645 140.215 ;
        RECT 100.835 139.495 101.005 140.625 ;
        RECT 101.805 140.555 101.975 140.785 ;
        RECT 101.175 140.385 101.975 140.555 ;
        RECT 101.175 139.835 101.345 140.385 ;
        RECT 102.155 140.215 102.440 140.615 ;
        RECT 101.575 140.185 101.940 140.215 ;
        RECT 101.565 140.015 101.940 140.185 ;
        RECT 102.110 140.015 102.440 140.215 ;
        RECT 102.710 140.215 102.990 140.615 ;
        RECT 103.170 140.555 103.340 140.785 ;
        RECT 103.565 140.725 103.895 141.205 ;
        RECT 104.065 140.555 104.235 141.035 ;
        RECT 103.170 140.385 104.235 140.555 ;
        RECT 104.495 140.455 105.705 141.205 ;
        RECT 105.875 140.480 106.165 141.205 ;
        RECT 106.340 140.635 106.660 141.035 ;
        RECT 102.710 140.015 103.185 140.215 ;
        RECT 103.355 140.015 103.800 140.215 ;
        RECT 103.970 140.005 104.320 140.215 ;
        RECT 104.495 139.915 105.015 140.455 ;
        RECT 101.175 139.665 104.235 139.835 ;
        RECT 105.185 139.745 105.705 140.285 ;
        RECT 106.340 139.845 106.510 140.635 ;
        RECT 106.830 140.385 107.140 141.205 ;
        RECT 107.310 140.575 107.640 141.035 ;
        RECT 107.810 140.745 108.060 141.205 ;
        RECT 108.250 140.825 110.300 141.035 ;
        RECT 108.250 140.575 109.000 140.655 ;
        RECT 107.310 140.385 109.000 140.575 ;
        RECT 109.170 140.385 109.340 140.825 ;
        RECT 109.510 140.385 110.300 140.655 ;
        RECT 110.475 140.575 110.815 141.035 ;
        RECT 110.985 140.745 111.155 141.205 ;
        RECT 111.325 140.825 112.495 141.035 ;
        RECT 111.325 140.575 111.575 140.825 ;
        RECT 112.165 140.805 112.495 140.825 ;
        RECT 110.475 140.405 111.575 140.575 ;
        RECT 111.745 140.385 112.605 140.635 ;
        RECT 112.775 140.385 113.035 141.205 ;
        RECT 113.205 140.385 113.535 140.805 ;
        RECT 113.715 140.720 114.505 140.985 ;
        RECT 106.680 140.015 107.030 140.215 ;
        RECT 107.310 140.015 107.990 140.215 ;
        RECT 108.200 140.015 109.390 140.215 ;
        RECT 109.570 139.845 109.900 140.215 ;
        RECT 100.300 138.655 100.645 139.475 ;
        RECT 100.835 138.825 101.090 139.495 ;
        RECT 101.260 138.655 101.590 139.415 ;
        RECT 101.760 139.255 103.395 139.495 ;
        RECT 101.760 138.825 102.010 139.255 ;
        RECT 103.165 139.165 103.395 139.255 ;
        RECT 102.180 138.655 102.535 139.075 ;
        RECT 102.725 138.995 103.055 139.035 ;
        RECT 103.565 138.995 103.895 139.495 ;
        RECT 102.725 138.825 103.895 138.995 ;
        RECT 104.065 138.825 104.235 139.665 ;
        RECT 104.495 138.655 105.705 139.745 ;
        RECT 105.875 138.655 106.165 139.820 ;
        RECT 106.340 139.675 109.900 139.845 ;
        RECT 106.340 139.225 106.510 139.675 ;
        RECT 110.100 139.505 110.300 140.385 ;
        RECT 110.475 139.965 111.235 140.215 ;
        RECT 111.405 139.965 112.155 140.215 ;
        RECT 112.325 139.795 112.605 140.385 ;
        RECT 113.285 140.295 113.535 140.385 ;
        RECT 106.340 138.825 106.660 139.225 ;
        RECT 106.830 138.655 107.140 139.455 ;
        RECT 107.310 139.335 110.300 139.505 ;
        RECT 107.310 139.285 108.480 139.335 ;
        RECT 107.310 138.825 107.640 139.285 ;
        RECT 107.810 138.655 107.980 139.115 ;
        RECT 108.150 138.825 108.480 139.285 ;
        RECT 109.510 139.285 110.300 139.335 ;
        RECT 108.650 138.655 108.900 139.115 ;
        RECT 109.090 138.655 109.340 139.115 ;
        RECT 109.510 138.825 109.760 139.285 ;
        RECT 110.010 138.655 110.300 139.115 ;
        RECT 110.475 138.655 110.735 139.795 ;
        RECT 110.905 139.625 112.605 139.795 ;
        RECT 110.905 138.825 111.235 139.625 ;
        RECT 111.405 138.655 111.575 139.455 ;
        RECT 111.745 138.825 112.075 139.625 ;
        RECT 112.245 138.655 112.500 139.455 ;
        RECT 112.775 139.335 113.115 140.215 ;
        RECT 113.285 140.045 114.080 140.295 ;
        RECT 112.775 138.655 113.035 139.165 ;
        RECT 113.285 138.825 113.455 140.045 ;
        RECT 114.250 139.865 114.505 140.720 ;
        RECT 114.675 140.565 114.875 140.985 ;
        RECT 115.065 140.745 115.395 141.205 ;
        RECT 114.675 140.045 115.085 140.565 ;
        RECT 115.565 140.555 115.825 141.035 ;
        RECT 116.045 140.815 116.375 141.205 ;
        RECT 116.545 140.635 116.715 140.955 ;
        RECT 116.885 140.815 117.215 141.205 ;
        RECT 117.630 140.805 118.585 140.975 ;
        RECT 115.255 139.865 115.485 140.295 ;
        RECT 113.695 139.695 115.485 139.865 ;
        RECT 113.695 139.330 113.945 139.695 ;
        RECT 114.115 139.335 114.445 139.525 ;
        RECT 114.665 139.400 115.380 139.695 ;
        RECT 115.655 139.525 115.825 140.555 ;
        RECT 114.115 139.160 114.310 139.335 ;
        RECT 113.695 138.655 114.310 139.160 ;
        RECT 114.480 138.825 114.955 139.165 ;
        RECT 115.125 138.655 115.340 139.200 ;
        RECT 115.550 138.825 115.825 139.525 ;
        RECT 115.995 140.465 118.245 140.635 ;
        RECT 115.995 139.505 116.165 140.465 ;
        RECT 116.335 139.845 116.580 140.295 ;
        RECT 116.750 140.015 117.300 140.215 ;
        RECT 117.470 140.045 117.845 140.215 ;
        RECT 117.470 139.845 117.640 140.045 ;
        RECT 118.015 139.965 118.245 140.465 ;
        RECT 116.335 139.675 117.640 139.845 ;
        RECT 118.415 139.925 118.585 140.805 ;
        RECT 118.755 140.370 119.045 141.205 ;
        RECT 119.215 140.260 119.555 141.035 ;
        RECT 119.725 140.745 119.895 141.205 ;
        RECT 120.135 140.770 120.495 141.035 ;
        RECT 120.135 140.765 120.490 140.770 ;
        RECT 120.135 140.755 120.485 140.765 ;
        RECT 120.135 140.750 120.480 140.755 ;
        RECT 120.135 140.740 120.475 140.750 ;
        RECT 121.125 140.745 121.295 141.205 ;
        RECT 120.135 140.735 120.470 140.740 ;
        RECT 120.135 140.725 120.460 140.735 ;
        RECT 120.135 140.715 120.450 140.725 ;
        RECT 120.135 140.575 120.435 140.715 ;
        RECT 119.725 140.385 120.435 140.575 ;
        RECT 120.625 140.575 120.955 140.655 ;
        RECT 121.465 140.575 121.805 141.035 ;
        RECT 120.625 140.385 121.805 140.575 ;
        RECT 121.975 140.465 122.705 141.030 ;
        RECT 118.415 139.755 119.045 139.925 ;
        RECT 115.995 138.825 116.375 139.505 ;
        RECT 116.965 138.655 117.135 139.505 ;
        RECT 117.305 139.335 118.545 139.505 ;
        RECT 117.305 138.825 117.635 139.335 ;
        RECT 117.805 138.655 117.975 139.165 ;
        RECT 118.145 138.825 118.545 139.335 ;
        RECT 118.725 138.825 119.045 139.755 ;
        RECT 119.215 138.825 119.495 140.260 ;
        RECT 119.725 139.815 120.010 140.385 ;
        RECT 120.195 139.985 120.665 140.215 ;
        RECT 120.835 140.195 121.165 140.215 ;
        RECT 120.835 140.015 121.285 140.195 ;
        RECT 121.475 140.015 121.805 140.215 ;
        RECT 119.725 139.600 120.875 139.815 ;
        RECT 119.665 138.655 120.375 139.430 ;
        RECT 120.545 138.825 120.875 139.600 ;
        RECT 121.070 138.900 121.285 140.015 ;
        RECT 121.575 139.675 121.805 140.015 ;
        RECT 121.975 139.965 122.320 140.295 ;
        RECT 121.465 138.655 121.795 139.375 ;
        RECT 121.975 138.655 122.320 139.795 ;
        RECT 122.490 138.825 122.705 140.465 ;
        RECT 122.950 140.555 123.280 141.035 ;
        RECT 123.465 140.725 123.635 141.205 ;
        RECT 123.805 140.555 124.135 141.035 ;
        RECT 122.950 140.385 124.135 140.555 ;
        RECT 124.305 140.385 124.475 141.205 ;
        RECT 125.285 140.555 125.455 141.035 ;
        RECT 125.625 140.725 125.955 141.205 ;
        RECT 126.180 140.785 127.715 141.035 ;
        RECT 126.180 140.555 126.350 140.785 ;
        RECT 125.285 140.385 126.350 140.555 ;
        RECT 126.530 140.215 126.810 140.615 ;
        RECT 122.950 139.965 123.425 140.215 ;
        RECT 122.950 138.885 123.190 139.965 ;
        RECT 123.595 138.825 124.040 140.215 ;
        RECT 124.210 139.965 124.560 140.215 ;
        RECT 125.200 140.005 125.550 140.215 ;
        RECT 125.720 140.015 126.165 140.215 ;
        RECT 126.335 140.015 126.810 140.215 ;
        RECT 127.080 140.215 127.365 140.615 ;
        RECT 127.545 140.555 127.715 140.785 ;
        RECT 127.885 140.725 128.215 141.205 ;
        RECT 128.430 140.705 128.685 141.035 ;
        RECT 128.500 140.625 128.685 140.705 ;
        RECT 127.545 140.385 128.345 140.555 ;
        RECT 127.080 140.015 127.410 140.215 ;
        RECT 127.580 140.185 127.945 140.215 ;
        RECT 127.580 140.015 127.955 140.185 ;
        RECT 128.175 139.835 128.345 140.385 ;
        RECT 124.210 138.655 124.560 139.795 ;
        RECT 125.285 139.665 128.345 139.835 ;
        RECT 125.285 138.825 125.455 139.665 ;
        RECT 128.515 139.505 128.685 140.625 ;
        RECT 128.895 140.475 129.185 141.205 ;
        RECT 128.885 139.965 129.185 140.295 ;
        RECT 129.365 140.275 129.595 140.915 ;
        RECT 129.775 140.655 130.085 141.025 ;
        RECT 130.265 140.835 130.935 141.205 ;
        RECT 129.775 140.455 131.005 140.655 ;
        RECT 129.365 139.965 129.890 140.275 ;
        RECT 130.070 139.965 130.535 140.275 ;
        RECT 130.715 139.785 131.005 140.455 ;
        RECT 128.475 139.495 128.685 139.505 ;
        RECT 125.625 138.995 125.955 139.495 ;
        RECT 126.125 139.255 127.760 139.495 ;
        RECT 126.125 139.165 126.355 139.255 ;
        RECT 126.465 138.995 126.795 139.035 ;
        RECT 125.625 138.825 126.795 138.995 ;
        RECT 126.985 138.655 127.340 139.075 ;
        RECT 127.510 138.825 127.760 139.255 ;
        RECT 127.930 138.655 128.260 139.415 ;
        RECT 128.430 138.825 128.685 139.495 ;
        RECT 128.895 139.545 130.055 139.785 ;
        RECT 128.895 138.835 129.155 139.545 ;
        RECT 129.325 138.655 129.655 139.365 ;
        RECT 129.825 138.835 130.055 139.545 ;
        RECT 130.235 139.565 131.005 139.785 ;
        RECT 130.235 138.835 130.505 139.565 ;
        RECT 130.685 138.655 131.025 139.385 ;
        RECT 131.195 138.835 131.455 141.025 ;
        RECT 131.635 140.480 131.925 141.205 ;
        RECT 132.095 140.260 132.435 141.035 ;
        RECT 132.605 140.745 132.775 141.205 ;
        RECT 133.015 140.770 133.375 141.035 ;
        RECT 133.015 140.765 133.370 140.770 ;
        RECT 133.015 140.755 133.365 140.765 ;
        RECT 133.015 140.750 133.360 140.755 ;
        RECT 133.015 140.740 133.355 140.750 ;
        RECT 134.005 140.745 134.175 141.205 ;
        RECT 133.015 140.735 133.350 140.740 ;
        RECT 133.015 140.725 133.340 140.735 ;
        RECT 133.015 140.715 133.330 140.725 ;
        RECT 133.015 140.575 133.315 140.715 ;
        RECT 132.605 140.385 133.315 140.575 ;
        RECT 133.505 140.575 133.835 140.655 ;
        RECT 134.345 140.575 134.685 141.035 ;
        RECT 133.505 140.385 134.685 140.575 ;
        RECT 135.935 140.385 136.225 141.205 ;
        RECT 136.395 140.475 136.725 141.035 ;
        RECT 131.635 138.655 131.925 139.820 ;
        RECT 132.095 138.825 132.375 140.260 ;
        RECT 132.605 139.815 132.890 140.385 ;
        RECT 136.475 140.215 136.725 140.475 ;
        RECT 136.905 140.385 137.195 141.205 ;
        RECT 137.365 140.565 137.695 141.035 ;
        RECT 137.865 140.735 138.035 141.205 ;
        RECT 138.205 140.565 138.535 141.035 ;
        RECT 138.705 140.735 138.875 141.205 ;
        RECT 139.045 140.565 139.375 141.035 ;
        RECT 139.545 140.735 139.715 141.205 ;
        RECT 139.885 140.565 140.215 141.035 ;
        RECT 137.365 140.385 140.215 140.565 ;
        RECT 140.385 140.385 140.665 141.205 ;
        RECT 140.835 140.385 141.095 141.205 ;
        RECT 141.265 140.385 141.595 140.805 ;
        RECT 141.775 140.720 142.565 140.985 ;
        RECT 133.075 139.985 133.545 140.215 ;
        RECT 133.715 140.195 134.045 140.215 ;
        RECT 133.715 140.015 134.165 140.195 ;
        RECT 134.355 140.015 134.685 140.215 ;
        RECT 132.605 139.600 133.755 139.815 ;
        RECT 132.545 138.655 133.255 139.430 ;
        RECT 133.425 138.825 133.755 139.600 ;
        RECT 133.950 138.900 134.165 140.015 ;
        RECT 134.455 139.675 134.685 140.015 ;
        RECT 135.775 139.970 136.305 140.215 ;
        RECT 136.475 140.015 137.955 140.215 ;
        RECT 134.345 138.655 134.675 139.375 ;
        RECT 135.820 138.655 136.225 139.795 ;
        RECT 136.475 139.715 136.725 140.015 ;
        RECT 138.125 139.845 138.455 140.385 ;
        RECT 141.345 140.295 141.595 140.385 ;
        RECT 138.950 140.015 140.390 140.215 ;
        RECT 136.395 138.825 136.725 139.715 ;
        RECT 136.895 138.995 137.275 139.715 ;
        RECT 137.445 139.545 138.455 139.845 ;
        RECT 137.445 139.165 137.615 139.545 ;
        RECT 137.785 138.995 138.115 139.355 ;
        RECT 138.285 139.165 138.455 139.545 ;
        RECT 138.625 139.625 140.665 139.835 ;
        RECT 138.625 138.995 138.955 139.625 ;
        RECT 136.895 138.825 138.955 138.995 ;
        RECT 139.125 138.655 139.375 139.455 ;
        RECT 139.545 138.825 139.715 139.625 ;
        RECT 139.885 138.655 140.215 139.455 ;
        RECT 140.385 138.825 140.665 139.625 ;
        RECT 140.835 139.335 141.175 140.215 ;
        RECT 141.345 140.045 142.140 140.295 ;
        RECT 140.835 138.655 141.095 139.165 ;
        RECT 141.345 138.825 141.515 140.045 ;
        RECT 142.310 139.865 142.565 140.720 ;
        RECT 142.735 140.565 142.935 140.985 ;
        RECT 143.125 140.745 143.455 141.205 ;
        RECT 142.735 140.045 143.145 140.565 ;
        RECT 143.625 140.555 143.885 141.035 ;
        RECT 143.315 139.865 143.545 140.295 ;
        RECT 141.755 139.695 143.545 139.865 ;
        RECT 141.755 139.330 142.005 139.695 ;
        RECT 142.175 139.335 142.505 139.525 ;
        RECT 142.725 139.400 143.440 139.695 ;
        RECT 143.715 139.525 143.885 140.555 ;
        RECT 142.175 139.160 142.370 139.335 ;
        RECT 141.755 138.655 142.370 139.160 ;
        RECT 142.540 138.825 143.015 139.165 ;
        RECT 143.185 138.655 143.400 139.200 ;
        RECT 143.610 138.825 143.885 139.525 ;
        RECT 144.055 140.555 144.315 141.035 ;
        RECT 144.485 140.745 144.815 141.205 ;
        RECT 145.005 140.565 145.205 140.985 ;
        RECT 144.055 139.525 144.225 140.555 ;
        RECT 144.395 139.865 144.625 140.295 ;
        RECT 144.795 140.045 145.205 140.565 ;
        RECT 145.375 140.720 146.165 140.985 ;
        RECT 145.375 139.865 145.630 140.720 ;
        RECT 146.345 140.385 146.675 140.805 ;
        RECT 146.845 140.385 147.105 141.205 ;
        RECT 147.275 140.405 147.970 141.035 ;
        RECT 148.175 140.405 148.485 141.205 ;
        RECT 148.655 140.660 154.000 141.205 ;
        RECT 146.345 140.295 146.595 140.385 ;
        RECT 145.800 140.045 146.595 140.295 ;
        RECT 144.395 139.695 146.185 139.865 ;
        RECT 144.055 138.825 144.330 139.525 ;
        RECT 144.500 139.400 145.215 139.695 ;
        RECT 145.435 139.335 145.765 139.525 ;
        RECT 144.540 138.655 144.755 139.200 ;
        RECT 144.925 138.825 145.400 139.165 ;
        RECT 145.570 139.160 145.765 139.335 ;
        RECT 145.935 139.330 146.185 139.695 ;
        RECT 145.570 138.655 146.185 139.160 ;
        RECT 146.425 138.825 146.595 140.045 ;
        RECT 146.765 139.335 147.105 140.215 ;
        RECT 147.295 139.965 147.630 140.215 ;
        RECT 147.800 139.805 147.970 140.405 ;
        RECT 148.140 139.965 148.475 140.235 ;
        RECT 150.240 139.830 150.580 140.660 ;
        RECT 154.175 140.435 156.765 141.205 ;
        RECT 156.935 140.455 158.145 141.205 ;
        RECT 146.845 138.655 147.105 139.165 ;
        RECT 147.275 138.655 147.535 139.795 ;
        RECT 147.705 138.825 148.035 139.805 ;
        RECT 148.205 138.655 148.485 139.795 ;
        RECT 152.060 139.090 152.410 140.340 ;
        RECT 154.175 139.915 155.385 140.435 ;
        RECT 155.555 139.745 156.765 140.265 ;
        RECT 148.655 138.655 154.000 139.090 ;
        RECT 154.175 138.655 156.765 139.745 ;
        RECT 156.935 139.745 157.455 140.285 ;
        RECT 157.625 139.915 158.145 140.455 ;
        RECT 156.935 138.655 158.145 139.745 ;
        RECT 2.750 138.485 158.230 138.655 ;
        RECT 2.835 137.395 4.045 138.485 ;
        RECT 4.220 137.815 4.475 138.315 ;
        RECT 4.645 137.985 4.975 138.485 ;
        RECT 4.220 137.645 4.970 137.815 ;
        RECT 2.835 136.685 3.355 137.225 ;
        RECT 3.525 136.855 4.045 137.395 ;
        RECT 4.220 136.825 4.570 137.475 ;
        RECT 2.835 135.935 4.045 136.685 ;
        RECT 4.740 136.655 4.970 137.645 ;
        RECT 4.220 136.485 4.970 136.655 ;
        RECT 4.220 136.195 4.475 136.485 ;
        RECT 4.645 135.935 4.975 136.315 ;
        RECT 5.145 136.195 5.315 138.315 ;
        RECT 5.485 137.515 5.810 138.300 ;
        RECT 5.980 138.025 6.230 138.485 ;
        RECT 6.400 137.985 6.650 138.315 ;
        RECT 6.865 137.985 7.545 138.315 ;
        RECT 6.400 137.855 6.570 137.985 ;
        RECT 6.175 137.685 6.570 137.855 ;
        RECT 5.545 136.465 6.005 137.515 ;
        RECT 6.175 136.325 6.345 137.685 ;
        RECT 6.740 137.425 7.205 137.815 ;
        RECT 6.515 136.615 6.865 137.235 ;
        RECT 7.035 136.835 7.205 137.425 ;
        RECT 7.375 137.205 7.545 137.985 ;
        RECT 7.715 137.885 7.885 138.225 ;
        RECT 8.120 138.055 8.450 138.485 ;
        RECT 8.620 137.885 8.790 138.225 ;
        RECT 9.085 138.025 9.455 138.485 ;
        RECT 7.715 137.715 8.790 137.885 ;
        RECT 9.625 137.855 9.795 138.315 ;
        RECT 10.030 137.975 10.900 138.315 ;
        RECT 11.070 138.025 11.320 138.485 ;
        RECT 9.235 137.685 9.795 137.855 ;
        RECT 9.235 137.545 9.405 137.685 ;
        RECT 7.905 137.375 9.405 137.545 ;
        RECT 10.100 137.515 10.560 137.805 ;
        RECT 7.375 137.035 9.065 137.205 ;
        RECT 7.035 136.615 7.390 136.835 ;
        RECT 7.560 136.325 7.730 137.035 ;
        RECT 7.935 136.615 8.725 136.865 ;
        RECT 8.895 136.855 9.065 137.035 ;
        RECT 9.235 136.685 9.405 137.375 ;
        RECT 5.675 135.935 6.005 136.295 ;
        RECT 6.175 136.155 6.670 136.325 ;
        RECT 6.875 136.155 7.730 136.325 ;
        RECT 8.605 135.935 8.935 136.395 ;
        RECT 9.145 136.295 9.405 136.685 ;
        RECT 9.595 137.505 10.560 137.515 ;
        RECT 10.730 137.595 10.900 137.975 ;
        RECT 11.490 137.935 11.660 138.225 ;
        RECT 11.840 138.105 12.170 138.485 ;
        RECT 11.490 137.765 12.290 137.935 ;
        RECT 9.595 137.345 10.270 137.505 ;
        RECT 10.730 137.425 11.950 137.595 ;
        RECT 9.595 136.555 9.805 137.345 ;
        RECT 10.730 137.335 10.900 137.425 ;
        RECT 9.975 136.555 10.325 137.175 ;
        RECT 10.495 137.165 10.900 137.335 ;
        RECT 10.495 136.385 10.665 137.165 ;
        RECT 10.835 136.715 11.055 136.995 ;
        RECT 11.235 136.885 11.775 137.255 ;
        RECT 12.120 137.175 12.290 137.765 ;
        RECT 12.510 137.345 12.815 138.485 ;
        RECT 12.985 137.295 13.240 138.175 ;
        RECT 12.120 137.145 12.860 137.175 ;
        RECT 10.835 136.545 11.365 136.715 ;
        RECT 9.145 136.125 9.495 136.295 ;
        RECT 9.715 136.105 10.665 136.385 ;
        RECT 10.835 135.935 11.025 136.375 ;
        RECT 11.195 136.315 11.365 136.545 ;
        RECT 11.535 136.485 11.775 136.885 ;
        RECT 11.945 136.845 12.860 137.145 ;
        RECT 11.945 136.670 12.270 136.845 ;
        RECT 11.945 136.315 12.265 136.670 ;
        RECT 13.030 136.645 13.240 137.295 ;
        RECT 11.195 136.145 12.265 136.315 ;
        RECT 12.510 135.935 12.815 136.395 ;
        RECT 12.985 136.115 13.240 136.645 ;
        RECT 14.335 137.410 14.605 138.315 ;
        RECT 14.775 137.725 15.105 138.485 ;
        RECT 15.285 137.555 15.455 138.315 ;
        RECT 14.335 136.610 14.505 137.410 ;
        RECT 14.790 137.385 15.455 137.555 ;
        RECT 14.790 137.240 14.960 137.385 ;
        RECT 15.715 137.320 16.005 138.485 ;
        RECT 16.180 137.345 16.515 138.315 ;
        RECT 16.685 137.345 16.855 138.485 ;
        RECT 17.025 138.145 19.055 138.315 ;
        RECT 14.675 136.910 14.960 137.240 ;
        RECT 14.790 136.655 14.960 136.910 ;
        RECT 15.195 136.835 15.525 137.205 ;
        RECT 16.180 136.675 16.350 137.345 ;
        RECT 17.025 137.175 17.195 138.145 ;
        RECT 16.520 136.845 16.775 137.175 ;
        RECT 17.000 136.845 17.195 137.175 ;
        RECT 17.365 137.805 18.490 137.975 ;
        RECT 16.605 136.675 16.775 136.845 ;
        RECT 17.365 136.675 17.535 137.805 ;
        RECT 14.335 136.105 14.595 136.610 ;
        RECT 14.790 136.485 15.455 136.655 ;
        RECT 14.775 135.935 15.105 136.315 ;
        RECT 15.285 136.105 15.455 136.485 ;
        RECT 15.715 135.935 16.005 136.660 ;
        RECT 16.180 136.105 16.435 136.675 ;
        RECT 16.605 136.505 17.535 136.675 ;
        RECT 17.705 137.465 18.715 137.635 ;
        RECT 17.705 136.665 17.875 137.465 ;
        RECT 17.360 136.470 17.535 136.505 ;
        RECT 16.605 135.935 16.935 136.335 ;
        RECT 17.360 136.105 17.890 136.470 ;
        RECT 18.080 136.445 18.355 137.265 ;
        RECT 18.075 136.275 18.355 136.445 ;
        RECT 18.080 136.105 18.355 136.275 ;
        RECT 18.525 136.105 18.715 137.465 ;
        RECT 18.885 137.480 19.055 138.145 ;
        RECT 19.225 137.725 19.395 138.485 ;
        RECT 19.630 137.725 20.145 138.135 ;
        RECT 18.885 137.290 19.635 137.480 ;
        RECT 19.805 136.915 20.145 137.725 ;
        RECT 20.315 137.395 21.985 138.485 ;
        RECT 22.160 137.815 22.415 138.315 ;
        RECT 22.585 137.985 22.915 138.485 ;
        RECT 22.160 137.645 22.910 137.815 ;
        RECT 18.915 136.745 20.145 136.915 ;
        RECT 18.895 135.935 19.405 136.470 ;
        RECT 19.625 136.140 19.870 136.745 ;
        RECT 20.315 136.705 21.065 137.225 ;
        RECT 21.235 136.875 21.985 137.395 ;
        RECT 22.160 136.825 22.510 137.475 ;
        RECT 20.315 135.935 21.985 136.705 ;
        RECT 22.680 136.655 22.910 137.645 ;
        RECT 22.160 136.485 22.910 136.655 ;
        RECT 22.160 136.195 22.415 136.485 ;
        RECT 22.585 135.935 22.915 136.315 ;
        RECT 23.085 136.195 23.255 138.315 ;
        RECT 23.425 137.515 23.750 138.300 ;
        RECT 23.920 138.025 24.170 138.485 ;
        RECT 24.340 137.985 24.590 138.315 ;
        RECT 24.805 137.985 25.485 138.315 ;
        RECT 24.340 137.855 24.510 137.985 ;
        RECT 24.115 137.685 24.510 137.855 ;
        RECT 23.485 136.465 23.945 137.515 ;
        RECT 24.115 136.325 24.285 137.685 ;
        RECT 24.680 137.425 25.145 137.815 ;
        RECT 24.455 136.615 24.805 137.235 ;
        RECT 24.975 136.835 25.145 137.425 ;
        RECT 25.315 137.205 25.485 137.985 ;
        RECT 25.655 137.885 25.825 138.225 ;
        RECT 26.060 138.055 26.390 138.485 ;
        RECT 26.560 137.885 26.730 138.225 ;
        RECT 27.025 138.025 27.395 138.485 ;
        RECT 25.655 137.715 26.730 137.885 ;
        RECT 27.565 137.855 27.735 138.315 ;
        RECT 27.970 137.975 28.840 138.315 ;
        RECT 29.010 138.025 29.260 138.485 ;
        RECT 27.175 137.685 27.735 137.855 ;
        RECT 27.175 137.545 27.345 137.685 ;
        RECT 25.845 137.375 27.345 137.545 ;
        RECT 28.040 137.515 28.500 137.805 ;
        RECT 25.315 137.035 27.005 137.205 ;
        RECT 24.975 136.615 25.330 136.835 ;
        RECT 25.500 136.325 25.670 137.035 ;
        RECT 25.875 136.615 26.665 136.865 ;
        RECT 26.835 136.855 27.005 137.035 ;
        RECT 27.175 136.685 27.345 137.375 ;
        RECT 23.615 135.935 23.945 136.295 ;
        RECT 24.115 136.155 24.610 136.325 ;
        RECT 24.815 136.155 25.670 136.325 ;
        RECT 26.545 135.935 26.875 136.395 ;
        RECT 27.085 136.295 27.345 136.685 ;
        RECT 27.535 137.505 28.500 137.515 ;
        RECT 28.670 137.595 28.840 137.975 ;
        RECT 29.430 137.935 29.600 138.225 ;
        RECT 29.780 138.105 30.110 138.485 ;
        RECT 29.430 137.765 30.230 137.935 ;
        RECT 27.535 137.345 28.210 137.505 ;
        RECT 28.670 137.425 29.890 137.595 ;
        RECT 27.535 136.555 27.745 137.345 ;
        RECT 28.670 137.335 28.840 137.425 ;
        RECT 27.915 136.555 28.265 137.175 ;
        RECT 28.435 137.165 28.840 137.335 ;
        RECT 28.435 136.385 28.605 137.165 ;
        RECT 28.775 136.715 28.995 136.995 ;
        RECT 29.175 136.885 29.715 137.255 ;
        RECT 30.060 137.175 30.230 137.765 ;
        RECT 30.450 137.345 30.755 138.485 ;
        RECT 30.925 137.295 31.180 138.175 ;
        RECT 30.060 137.145 30.800 137.175 ;
        RECT 28.775 136.545 29.305 136.715 ;
        RECT 27.085 136.125 27.435 136.295 ;
        RECT 27.655 136.105 28.605 136.385 ;
        RECT 28.775 135.935 28.965 136.375 ;
        RECT 29.135 136.315 29.305 136.545 ;
        RECT 29.475 136.485 29.715 136.885 ;
        RECT 29.885 136.845 30.800 137.145 ;
        RECT 29.885 136.670 30.210 136.845 ;
        RECT 29.885 136.315 30.205 136.670 ;
        RECT 30.970 136.645 31.180 137.295 ;
        RECT 29.135 136.145 30.205 136.315 ;
        RECT 30.450 135.935 30.755 136.395 ;
        RECT 30.925 136.115 31.180 136.645 ;
        RECT 32.280 137.295 32.535 138.175 ;
        RECT 32.705 137.345 33.010 138.485 ;
        RECT 33.350 138.105 33.680 138.485 ;
        RECT 33.860 137.935 34.030 138.225 ;
        RECT 34.200 138.025 34.450 138.485 ;
        RECT 33.230 137.765 34.030 137.935 ;
        RECT 34.620 137.975 35.490 138.315 ;
        RECT 32.280 136.645 32.490 137.295 ;
        RECT 33.230 137.175 33.400 137.765 ;
        RECT 34.620 137.595 34.790 137.975 ;
        RECT 35.725 137.855 35.895 138.315 ;
        RECT 36.065 138.025 36.435 138.485 ;
        RECT 36.730 137.885 36.900 138.225 ;
        RECT 37.070 138.055 37.400 138.485 ;
        RECT 37.635 137.885 37.805 138.225 ;
        RECT 33.570 137.425 34.790 137.595 ;
        RECT 34.960 137.515 35.420 137.805 ;
        RECT 35.725 137.685 36.285 137.855 ;
        RECT 36.730 137.715 37.805 137.885 ;
        RECT 37.975 137.985 38.655 138.315 ;
        RECT 38.870 137.985 39.120 138.315 ;
        RECT 39.290 138.025 39.540 138.485 ;
        RECT 36.115 137.545 36.285 137.685 ;
        RECT 34.960 137.505 35.925 137.515 ;
        RECT 34.620 137.335 34.790 137.425 ;
        RECT 35.250 137.345 35.925 137.505 ;
        RECT 32.660 137.145 33.400 137.175 ;
        RECT 32.660 136.845 33.575 137.145 ;
        RECT 33.250 136.670 33.575 136.845 ;
        RECT 32.280 136.115 32.535 136.645 ;
        RECT 32.705 135.935 33.010 136.395 ;
        RECT 33.255 136.315 33.575 136.670 ;
        RECT 33.745 136.885 34.285 137.255 ;
        RECT 34.620 137.165 35.025 137.335 ;
        RECT 33.745 136.485 33.985 136.885 ;
        RECT 34.465 136.715 34.685 136.995 ;
        RECT 34.155 136.545 34.685 136.715 ;
        RECT 34.155 136.315 34.325 136.545 ;
        RECT 34.855 136.385 35.025 137.165 ;
        RECT 35.195 136.555 35.545 137.175 ;
        RECT 35.715 136.555 35.925 137.345 ;
        RECT 36.115 137.375 37.615 137.545 ;
        RECT 36.115 136.685 36.285 137.375 ;
        RECT 37.975 137.205 38.145 137.985 ;
        RECT 38.950 137.855 39.120 137.985 ;
        RECT 36.455 137.035 38.145 137.205 ;
        RECT 38.315 137.425 38.780 137.815 ;
        RECT 38.950 137.685 39.345 137.855 ;
        RECT 36.455 136.855 36.625 137.035 ;
        RECT 33.255 136.145 34.325 136.315 ;
        RECT 34.495 135.935 34.685 136.375 ;
        RECT 34.855 136.105 35.805 136.385 ;
        RECT 36.115 136.295 36.375 136.685 ;
        RECT 36.795 136.615 37.585 136.865 ;
        RECT 36.025 136.125 36.375 136.295 ;
        RECT 36.585 135.935 36.915 136.395 ;
        RECT 37.790 136.325 37.960 137.035 ;
        RECT 38.315 136.835 38.485 137.425 ;
        RECT 38.130 136.615 38.485 136.835 ;
        RECT 38.655 136.615 39.005 137.235 ;
        RECT 39.175 136.325 39.345 137.685 ;
        RECT 39.710 137.515 40.035 138.300 ;
        RECT 39.515 136.465 39.975 137.515 ;
        RECT 37.790 136.155 38.645 136.325 ;
        RECT 38.850 136.155 39.345 136.325 ;
        RECT 39.515 135.935 39.845 136.295 ;
        RECT 40.205 136.195 40.375 138.315 ;
        RECT 40.545 137.985 40.875 138.485 ;
        RECT 41.045 137.815 41.300 138.315 ;
        RECT 40.550 137.645 41.300 137.815 ;
        RECT 40.550 136.655 40.780 137.645 ;
        RECT 40.950 136.825 41.300 137.475 ;
        RECT 41.475 137.320 41.765 138.485 ;
        RECT 42.860 137.815 43.115 138.315 ;
        RECT 43.285 137.985 43.615 138.485 ;
        RECT 42.860 137.645 43.610 137.815 ;
        RECT 42.860 136.825 43.210 137.475 ;
        RECT 40.550 136.485 41.300 136.655 ;
        RECT 40.545 135.935 40.875 136.315 ;
        RECT 41.045 136.195 41.300 136.485 ;
        RECT 41.475 135.935 41.765 136.660 ;
        RECT 43.380 136.655 43.610 137.645 ;
        RECT 42.860 136.485 43.610 136.655 ;
        RECT 42.860 136.195 43.115 136.485 ;
        RECT 43.285 135.935 43.615 136.315 ;
        RECT 43.785 136.195 43.955 138.315 ;
        RECT 44.125 137.515 44.450 138.300 ;
        RECT 44.620 138.025 44.870 138.485 ;
        RECT 45.040 137.985 45.290 138.315 ;
        RECT 45.505 137.985 46.185 138.315 ;
        RECT 45.040 137.855 45.210 137.985 ;
        RECT 44.815 137.685 45.210 137.855 ;
        RECT 44.185 136.465 44.645 137.515 ;
        RECT 44.815 136.325 44.985 137.685 ;
        RECT 45.380 137.425 45.845 137.815 ;
        RECT 45.155 136.615 45.505 137.235 ;
        RECT 45.675 136.835 45.845 137.425 ;
        RECT 46.015 137.205 46.185 137.985 ;
        RECT 46.355 137.885 46.525 138.225 ;
        RECT 46.760 138.055 47.090 138.485 ;
        RECT 47.260 137.885 47.430 138.225 ;
        RECT 47.725 138.025 48.095 138.485 ;
        RECT 46.355 137.715 47.430 137.885 ;
        RECT 48.265 137.855 48.435 138.315 ;
        RECT 48.670 137.975 49.540 138.315 ;
        RECT 49.710 138.025 49.960 138.485 ;
        RECT 47.875 137.685 48.435 137.855 ;
        RECT 47.875 137.545 48.045 137.685 ;
        RECT 46.545 137.375 48.045 137.545 ;
        RECT 48.740 137.515 49.200 137.805 ;
        RECT 46.015 137.035 47.705 137.205 ;
        RECT 45.675 136.615 46.030 136.835 ;
        RECT 46.200 136.325 46.370 137.035 ;
        RECT 46.575 136.615 47.365 136.865 ;
        RECT 47.535 136.855 47.705 137.035 ;
        RECT 47.875 136.685 48.045 137.375 ;
        RECT 44.315 135.935 44.645 136.295 ;
        RECT 44.815 136.155 45.310 136.325 ;
        RECT 45.515 136.155 46.370 136.325 ;
        RECT 47.245 135.935 47.575 136.395 ;
        RECT 47.785 136.295 48.045 136.685 ;
        RECT 48.235 137.505 49.200 137.515 ;
        RECT 49.370 137.595 49.540 137.975 ;
        RECT 50.130 137.935 50.300 138.225 ;
        RECT 50.480 138.105 50.810 138.485 ;
        RECT 50.130 137.765 50.930 137.935 ;
        RECT 48.235 137.345 48.910 137.505 ;
        RECT 49.370 137.425 50.590 137.595 ;
        RECT 48.235 136.555 48.445 137.345 ;
        RECT 49.370 137.335 49.540 137.425 ;
        RECT 48.615 136.555 48.965 137.175 ;
        RECT 49.135 137.165 49.540 137.335 ;
        RECT 49.135 136.385 49.305 137.165 ;
        RECT 49.475 136.715 49.695 136.995 ;
        RECT 49.875 136.885 50.415 137.255 ;
        RECT 50.760 137.175 50.930 137.765 ;
        RECT 51.150 137.345 51.455 138.485 ;
        RECT 51.625 137.295 51.880 138.175 ;
        RECT 52.605 137.555 52.775 138.315 ;
        RECT 52.955 137.725 53.285 138.485 ;
        RECT 52.605 137.385 53.270 137.555 ;
        RECT 53.455 137.410 53.725 138.315 ;
        RECT 50.760 137.145 51.500 137.175 ;
        RECT 49.475 136.545 50.005 136.715 ;
        RECT 47.785 136.125 48.135 136.295 ;
        RECT 48.355 136.105 49.305 136.385 ;
        RECT 49.475 135.935 49.665 136.375 ;
        RECT 49.835 136.315 50.005 136.545 ;
        RECT 50.175 136.485 50.415 136.885 ;
        RECT 50.585 136.845 51.500 137.145 ;
        RECT 50.585 136.670 50.910 136.845 ;
        RECT 50.585 136.315 50.905 136.670 ;
        RECT 51.670 136.645 51.880 137.295 ;
        RECT 53.100 137.240 53.270 137.385 ;
        RECT 52.535 136.835 52.865 137.205 ;
        RECT 53.100 136.910 53.385 137.240 ;
        RECT 53.100 136.655 53.270 136.910 ;
        RECT 49.835 136.145 50.905 136.315 ;
        RECT 51.150 135.935 51.455 136.395 ;
        RECT 51.625 136.115 51.880 136.645 ;
        RECT 52.605 136.485 53.270 136.655 ;
        RECT 53.555 136.610 53.725 137.410 ;
        RECT 52.605 136.105 52.775 136.485 ;
        RECT 52.955 135.935 53.285 136.315 ;
        RECT 53.465 136.105 53.725 136.610 ;
        RECT 53.900 137.345 54.235 138.315 ;
        RECT 54.405 137.345 54.575 138.485 ;
        RECT 54.745 138.145 56.775 138.315 ;
        RECT 53.900 136.675 54.070 137.345 ;
        RECT 54.745 137.175 54.915 138.145 ;
        RECT 54.240 136.845 54.495 137.175 ;
        RECT 54.720 136.845 54.915 137.175 ;
        RECT 55.085 137.805 56.210 137.975 ;
        RECT 54.325 136.675 54.495 136.845 ;
        RECT 55.085 136.675 55.255 137.805 ;
        RECT 53.900 136.105 54.155 136.675 ;
        RECT 54.325 136.505 55.255 136.675 ;
        RECT 55.425 137.465 56.435 137.635 ;
        RECT 55.425 136.665 55.595 137.465 ;
        RECT 55.800 137.125 56.075 137.265 ;
        RECT 55.795 136.955 56.075 137.125 ;
        RECT 55.080 136.470 55.255 136.505 ;
        RECT 54.325 135.935 54.655 136.335 ;
        RECT 55.080 136.105 55.610 136.470 ;
        RECT 55.800 136.105 56.075 136.955 ;
        RECT 56.245 136.105 56.435 137.465 ;
        RECT 56.605 137.480 56.775 138.145 ;
        RECT 56.945 137.725 57.115 138.485 ;
        RECT 57.350 137.725 57.865 138.135 ;
        RECT 56.605 137.290 57.355 137.480 ;
        RECT 57.525 136.915 57.865 137.725 ;
        RECT 58.040 137.815 58.295 138.315 ;
        RECT 58.465 137.985 58.795 138.485 ;
        RECT 58.040 137.645 58.790 137.815 ;
        RECT 56.635 136.745 57.865 136.915 ;
        RECT 58.040 136.825 58.390 137.475 ;
        RECT 56.615 135.935 57.125 136.470 ;
        RECT 57.345 136.140 57.590 136.745 ;
        RECT 58.560 136.655 58.790 137.645 ;
        RECT 58.040 136.485 58.790 136.655 ;
        RECT 58.040 136.195 58.295 136.485 ;
        RECT 58.465 135.935 58.795 136.315 ;
        RECT 58.965 136.195 59.135 138.315 ;
        RECT 59.305 137.515 59.630 138.300 ;
        RECT 59.800 138.025 60.050 138.485 ;
        RECT 60.220 137.985 60.470 138.315 ;
        RECT 60.685 137.985 61.365 138.315 ;
        RECT 60.220 137.855 60.390 137.985 ;
        RECT 59.995 137.685 60.390 137.855 ;
        RECT 59.365 136.465 59.825 137.515 ;
        RECT 59.995 136.325 60.165 137.685 ;
        RECT 60.560 137.425 61.025 137.815 ;
        RECT 60.335 136.615 60.685 137.235 ;
        RECT 60.855 136.835 61.025 137.425 ;
        RECT 61.195 137.205 61.365 137.985 ;
        RECT 61.535 137.885 61.705 138.225 ;
        RECT 61.940 138.055 62.270 138.485 ;
        RECT 62.440 137.885 62.610 138.225 ;
        RECT 62.905 138.025 63.275 138.485 ;
        RECT 61.535 137.715 62.610 137.885 ;
        RECT 63.445 137.855 63.615 138.315 ;
        RECT 63.850 137.975 64.720 138.315 ;
        RECT 64.890 138.025 65.140 138.485 ;
        RECT 63.055 137.685 63.615 137.855 ;
        RECT 63.055 137.545 63.225 137.685 ;
        RECT 61.725 137.375 63.225 137.545 ;
        RECT 63.920 137.515 64.380 137.805 ;
        RECT 61.195 137.035 62.885 137.205 ;
        RECT 60.855 136.615 61.210 136.835 ;
        RECT 61.380 136.325 61.550 137.035 ;
        RECT 61.755 136.615 62.545 136.865 ;
        RECT 62.715 136.855 62.885 137.035 ;
        RECT 63.055 136.685 63.225 137.375 ;
        RECT 59.495 135.935 59.825 136.295 ;
        RECT 59.995 136.155 60.490 136.325 ;
        RECT 60.695 136.155 61.550 136.325 ;
        RECT 62.425 135.935 62.755 136.395 ;
        RECT 62.965 136.295 63.225 136.685 ;
        RECT 63.415 137.505 64.380 137.515 ;
        RECT 64.550 137.595 64.720 137.975 ;
        RECT 65.310 137.935 65.480 138.225 ;
        RECT 65.660 138.105 65.990 138.485 ;
        RECT 65.310 137.765 66.110 137.935 ;
        RECT 63.415 137.345 64.090 137.505 ;
        RECT 64.550 137.425 65.770 137.595 ;
        RECT 63.415 136.555 63.625 137.345 ;
        RECT 64.550 137.335 64.720 137.425 ;
        RECT 63.795 136.555 64.145 137.175 ;
        RECT 64.315 137.165 64.720 137.335 ;
        RECT 64.315 136.385 64.485 137.165 ;
        RECT 64.655 136.715 64.875 136.995 ;
        RECT 65.055 136.885 65.595 137.255 ;
        RECT 65.940 137.175 66.110 137.765 ;
        RECT 66.330 137.345 66.635 138.485 ;
        RECT 66.805 137.295 67.060 138.175 ;
        RECT 67.235 137.320 67.525 138.485 ;
        RECT 67.755 137.345 67.965 138.485 ;
        RECT 68.135 137.335 68.465 138.315 ;
        RECT 68.635 137.345 68.865 138.485 ;
        RECT 69.080 137.345 69.430 138.485 ;
        RECT 65.940 137.145 66.680 137.175 ;
        RECT 64.655 136.545 65.185 136.715 ;
        RECT 62.965 136.125 63.315 136.295 ;
        RECT 63.535 136.105 64.485 136.385 ;
        RECT 64.655 135.935 64.845 136.375 ;
        RECT 65.015 136.315 65.185 136.545 ;
        RECT 65.355 136.485 65.595 136.885 ;
        RECT 65.765 136.845 66.680 137.145 ;
        RECT 65.765 136.670 66.090 136.845 ;
        RECT 65.765 136.315 66.085 136.670 ;
        RECT 66.850 136.645 67.060 137.295 ;
        RECT 65.015 136.145 66.085 136.315 ;
        RECT 66.330 135.935 66.635 136.395 ;
        RECT 66.805 136.115 67.060 136.645 ;
        RECT 67.235 135.935 67.525 136.660 ;
        RECT 67.755 135.935 67.965 136.755 ;
        RECT 68.135 136.735 68.385 137.335 ;
        RECT 68.555 136.925 68.885 137.175 ;
        RECT 69.080 136.925 69.430 137.175 ;
        RECT 69.600 136.925 70.045 138.315 ;
        RECT 70.450 137.175 70.690 138.255 ;
        RECT 70.215 136.925 70.690 137.175 ;
        RECT 68.135 136.105 68.465 136.735 ;
        RECT 68.635 135.935 68.865 136.755 ;
        RECT 69.165 135.935 69.335 136.755 ;
        RECT 69.505 136.585 70.690 136.755 ;
        RECT 69.505 136.105 69.835 136.585 ;
        RECT 70.005 135.935 70.175 136.415 ;
        RECT 70.360 136.105 70.690 136.585 ;
        RECT 70.935 136.675 71.150 138.315 ;
        RECT 71.320 137.345 71.665 138.485 ;
        RECT 71.835 137.975 72.135 138.485 ;
        RECT 72.305 137.805 72.635 138.315 ;
        RECT 72.805 137.975 73.435 138.485 ;
        RECT 74.015 137.975 74.395 138.145 ;
        RECT 74.565 137.975 74.865 138.485 ;
        RECT 74.225 137.805 74.395 137.975 ;
        RECT 71.835 137.635 74.055 137.805 ;
        RECT 71.320 136.845 71.665 137.175 ;
        RECT 71.835 136.675 72.005 137.635 ;
        RECT 72.175 137.295 73.715 137.465 ;
        RECT 72.175 136.845 72.420 137.295 ;
        RECT 72.680 136.925 73.375 137.125 ;
        RECT 73.545 137.095 73.715 137.295 ;
        RECT 73.885 137.435 74.055 137.635 ;
        RECT 74.225 137.605 74.885 137.805 ;
        RECT 73.885 137.265 74.545 137.435 ;
        RECT 73.545 136.925 74.145 137.095 ;
        RECT 74.375 136.845 74.545 137.265 ;
        RECT 70.935 136.110 71.665 136.675 ;
        RECT 71.835 136.130 72.300 136.675 ;
        RECT 72.805 135.935 72.975 136.755 ;
        RECT 73.145 136.675 74.055 136.755 ;
        RECT 74.715 136.675 74.885 137.605 ;
        RECT 75.055 137.395 76.725 138.485 ;
        RECT 77.445 137.865 77.615 138.295 ;
        RECT 77.785 138.035 78.115 138.485 ;
        RECT 77.445 137.635 78.120 137.865 ;
        RECT 73.145 136.585 74.395 136.675 ;
        RECT 73.145 136.105 73.475 136.585 ;
        RECT 73.885 136.505 74.395 136.585 ;
        RECT 73.645 135.935 73.995 136.325 ;
        RECT 74.165 136.105 74.395 136.505 ;
        RECT 74.565 136.195 74.885 136.675 ;
        RECT 75.055 136.705 75.805 137.225 ;
        RECT 75.975 136.875 76.725 137.395 ;
        RECT 75.055 135.935 76.725 136.705 ;
        RECT 77.415 136.615 77.715 137.465 ;
        RECT 77.885 136.985 78.120 137.635 ;
        RECT 78.290 137.325 78.575 138.270 ;
        RECT 78.755 138.015 79.440 138.485 ;
        RECT 78.750 137.495 79.445 137.805 ;
        RECT 79.620 137.430 79.925 138.215 ;
        RECT 78.290 137.175 79.150 137.325 ;
        RECT 78.290 137.155 79.575 137.175 ;
        RECT 77.885 136.655 78.420 136.985 ;
        RECT 78.590 136.795 79.575 137.155 ;
        RECT 77.885 136.505 78.105 136.655 ;
        RECT 77.360 135.935 77.695 136.440 ;
        RECT 77.865 136.130 78.105 136.505 ;
        RECT 78.590 136.460 78.760 136.795 ;
        RECT 79.750 136.625 79.925 137.430 ;
        RECT 80.125 137.875 80.455 138.305 ;
        RECT 80.635 138.045 80.830 138.485 ;
        RECT 81.000 137.875 81.330 138.305 ;
        RECT 80.125 137.705 81.330 137.875 ;
        RECT 80.125 137.375 81.020 137.705 ;
        RECT 81.500 137.535 81.775 138.305 ;
        RECT 81.190 137.345 81.775 137.535 ;
        RECT 81.955 137.395 83.165 138.485 ;
        RECT 83.335 137.975 83.635 138.485 ;
        RECT 83.805 137.805 84.135 138.315 ;
        RECT 84.305 137.975 84.935 138.485 ;
        RECT 85.515 137.975 85.895 138.145 ;
        RECT 86.065 137.975 86.365 138.485 ;
        RECT 85.725 137.805 85.895 137.975 ;
        RECT 80.130 136.845 80.425 137.175 ;
        RECT 80.605 136.845 81.020 137.175 ;
        RECT 78.385 136.265 78.760 136.460 ;
        RECT 78.385 136.120 78.555 136.265 ;
        RECT 79.120 135.935 79.515 136.430 ;
        RECT 79.685 136.105 79.925 136.625 ;
        RECT 80.125 135.935 80.425 136.665 ;
        RECT 80.605 136.225 80.835 136.845 ;
        RECT 81.190 136.675 81.365 137.345 ;
        RECT 81.035 136.495 81.365 136.675 ;
        RECT 81.535 136.525 81.775 137.175 ;
        RECT 81.955 136.685 82.475 137.225 ;
        RECT 82.645 136.855 83.165 137.395 ;
        RECT 83.335 137.635 85.555 137.805 ;
        RECT 81.035 136.115 81.260 136.495 ;
        RECT 81.430 135.935 81.760 136.325 ;
        RECT 81.955 135.935 83.165 136.685 ;
        RECT 83.335 136.675 83.505 137.635 ;
        RECT 83.675 137.295 85.215 137.465 ;
        RECT 83.675 136.845 83.920 137.295 ;
        RECT 84.180 136.925 84.875 137.125 ;
        RECT 85.045 137.095 85.215 137.295 ;
        RECT 85.385 137.435 85.555 137.635 ;
        RECT 85.725 137.605 86.385 137.805 ;
        RECT 85.385 137.265 86.045 137.435 ;
        RECT 85.045 136.925 85.645 137.095 ;
        RECT 85.875 136.845 86.045 137.265 ;
        RECT 83.335 136.130 83.800 136.675 ;
        RECT 84.305 135.935 84.475 136.755 ;
        RECT 84.645 136.675 85.555 136.755 ;
        RECT 86.215 136.675 86.385 137.605 ;
        RECT 84.645 136.585 85.895 136.675 ;
        RECT 84.645 136.105 84.975 136.585 ;
        RECT 85.385 136.505 85.895 136.585 ;
        RECT 85.145 135.935 85.495 136.325 ;
        RECT 85.665 136.105 85.895 136.505 ;
        RECT 86.065 136.195 86.385 136.675 ;
        RECT 86.555 137.345 86.825 138.315 ;
        RECT 87.035 137.685 87.315 138.485 ;
        RECT 87.495 137.935 88.690 138.265 ;
        RECT 87.820 137.515 88.240 137.765 ;
        RECT 86.995 137.345 88.240 137.515 ;
        RECT 86.555 137.295 86.785 137.345 ;
        RECT 86.555 136.610 86.725 137.295 ;
        RECT 86.995 137.175 87.165 137.345 ;
        RECT 88.465 137.175 88.635 137.735 ;
        RECT 88.885 137.345 89.140 138.485 ;
        RECT 89.325 137.425 89.655 138.275 ;
        RECT 86.935 136.845 87.165 137.175 ;
        RECT 87.895 136.845 88.635 137.175 ;
        RECT 88.805 136.925 89.140 137.175 ;
        RECT 86.995 136.675 87.165 136.845 ;
        RECT 88.385 136.755 88.635 136.845 ;
        RECT 86.555 136.265 86.825 136.610 ;
        RECT 86.995 136.505 87.735 136.675 ;
        RECT 88.385 136.585 89.120 136.755 ;
        RECT 87.015 135.935 87.395 136.335 ;
        RECT 87.565 136.155 87.735 136.505 ;
        RECT 87.905 135.935 88.640 136.415 ;
        RECT 88.810 136.115 89.120 136.585 ;
        RECT 89.325 136.660 89.515 137.425 ;
        RECT 89.825 137.345 90.075 138.485 ;
        RECT 90.265 137.845 90.515 138.265 ;
        RECT 90.745 138.015 91.075 138.485 ;
        RECT 91.305 137.845 91.555 138.265 ;
        RECT 90.265 137.675 91.555 137.845 ;
        RECT 91.735 137.845 92.065 138.275 ;
        RECT 91.735 137.675 92.190 137.845 ;
        RECT 90.255 137.175 90.470 137.505 ;
        RECT 89.685 136.845 89.995 137.175 ;
        RECT 90.165 136.845 90.470 137.175 ;
        RECT 90.645 136.845 90.930 137.505 ;
        RECT 91.125 136.845 91.390 137.505 ;
        RECT 91.605 136.845 91.850 137.505 ;
        RECT 89.825 136.675 89.995 136.845 ;
        RECT 92.020 136.675 92.190 137.675 ;
        RECT 92.995 137.320 93.285 138.485 ;
        RECT 93.455 137.395 96.045 138.485 ;
        RECT 89.325 136.150 89.655 136.660 ;
        RECT 89.825 136.505 92.190 136.675 ;
        RECT 93.455 136.705 94.665 137.225 ;
        RECT 94.835 136.875 96.045 137.395 ;
        RECT 96.215 137.345 96.490 138.315 ;
        RECT 96.700 137.685 96.980 138.485 ;
        RECT 97.150 137.975 98.765 138.305 ;
        RECT 97.150 137.635 98.325 137.805 ;
        RECT 97.150 137.515 97.320 137.635 ;
        RECT 96.660 137.345 97.320 137.515 ;
        RECT 89.825 135.935 90.155 136.335 ;
        RECT 91.205 136.165 91.535 136.505 ;
        RECT 91.705 135.935 92.035 136.335 ;
        RECT 92.995 135.935 93.285 136.660 ;
        RECT 93.455 135.935 96.045 136.705 ;
        RECT 96.215 136.610 96.385 137.345 ;
        RECT 96.660 137.175 96.830 137.345 ;
        RECT 97.580 137.175 97.825 137.465 ;
        RECT 97.995 137.345 98.325 137.635 ;
        RECT 98.585 137.175 98.755 137.735 ;
        RECT 99.005 137.345 99.265 138.485 ;
        RECT 99.435 137.395 102.025 138.485 ;
        RECT 96.555 136.845 96.830 137.175 ;
        RECT 97.000 136.845 97.825 137.175 ;
        RECT 98.040 136.845 98.755 137.175 ;
        RECT 98.925 136.925 99.260 137.175 ;
        RECT 96.660 136.675 96.830 136.845 ;
        RECT 98.505 136.755 98.755 136.845 ;
        RECT 96.215 136.265 96.490 136.610 ;
        RECT 96.660 136.505 98.325 136.675 ;
        RECT 96.680 135.935 97.055 136.335 ;
        RECT 97.225 136.155 97.395 136.505 ;
        RECT 97.565 135.935 97.895 136.335 ;
        RECT 98.065 136.105 98.325 136.505 ;
        RECT 98.505 136.335 98.835 136.755 ;
        RECT 99.005 135.935 99.265 136.755 ;
        RECT 99.435 136.705 100.645 137.225 ;
        RECT 100.815 136.875 102.025 137.395 ;
        RECT 102.655 137.345 102.930 138.315 ;
        RECT 103.140 137.685 103.420 138.485 ;
        RECT 103.590 137.975 105.205 138.305 ;
        RECT 103.590 137.635 104.765 137.805 ;
        RECT 103.590 137.515 103.760 137.635 ;
        RECT 103.100 137.345 103.760 137.515 ;
        RECT 99.435 135.935 102.025 136.705 ;
        RECT 102.655 136.610 102.825 137.345 ;
        RECT 103.100 137.175 103.270 137.345 ;
        RECT 104.020 137.175 104.265 137.465 ;
        RECT 104.435 137.345 104.765 137.635 ;
        RECT 105.025 137.175 105.195 137.735 ;
        RECT 105.445 137.345 105.705 138.485 ;
        RECT 106.010 137.675 106.260 138.485 ;
        RECT 106.430 137.465 106.680 138.315 ;
        RECT 106.850 137.645 107.100 138.485 ;
        RECT 107.270 137.465 107.520 138.315 ;
        RECT 107.690 137.975 108.460 138.485 ;
        RECT 108.630 138.145 109.720 138.315 ;
        RECT 108.630 137.975 108.880 138.145 ;
        RECT 109.470 137.975 109.720 138.145 ;
        RECT 109.890 137.975 110.220 138.485 ;
        RECT 110.390 138.145 111.480 138.315 ;
        RECT 110.390 137.975 110.640 138.145 ;
        RECT 109.050 137.805 109.300 137.975 ;
        RECT 110.810 137.805 111.060 137.975 ;
        RECT 105.875 137.295 107.520 137.465 ;
        RECT 107.690 137.635 111.060 137.805 ;
        RECT 111.230 137.635 111.480 138.145 ;
        RECT 102.995 136.845 103.270 137.175 ;
        RECT 103.440 136.845 104.265 137.175 ;
        RECT 104.480 136.845 105.195 137.175 ;
        RECT 105.365 136.925 105.700 137.175 ;
        RECT 103.100 136.675 103.270 136.845 ;
        RECT 104.945 136.755 105.195 136.845 ;
        RECT 105.875 136.755 106.160 137.295 ;
        RECT 107.690 137.125 108.020 137.635 ;
        RECT 106.330 136.925 108.020 137.125 ;
        RECT 108.210 137.295 109.970 137.465 ;
        RECT 108.210 136.925 108.745 137.295 ;
        RECT 108.915 136.925 109.470 137.125 ;
        RECT 109.640 136.925 109.970 137.295 ;
        RECT 110.140 137.295 111.525 137.465 ;
        RECT 111.695 137.305 111.900 138.485 ;
        RECT 112.315 137.345 112.590 138.315 ;
        RECT 112.800 137.685 113.080 138.485 ;
        RECT 113.250 138.145 113.890 138.305 ;
        RECT 113.250 137.975 113.925 138.145 ;
        RECT 114.115 138.055 114.860 138.225 ;
        RECT 115.525 138.055 115.855 138.485 ;
        RECT 114.115 137.805 114.285 138.055 ;
        RECT 116.025 137.885 116.285 138.305 ;
        RECT 113.250 137.635 114.285 137.805 ;
        RECT 114.455 137.715 116.285 137.885 ;
        RECT 113.250 137.515 113.420 137.635 ;
        RECT 112.760 137.345 113.420 137.515 ;
        RECT 114.455 137.435 114.625 137.715 ;
        RECT 110.140 136.925 110.470 137.295 ;
        RECT 111.355 137.125 111.525 137.295 ;
        RECT 110.690 136.925 111.185 137.125 ;
        RECT 111.355 136.925 112.145 137.125 ;
        RECT 107.730 136.755 108.020 136.925 ;
        RECT 102.655 136.265 102.930 136.610 ;
        RECT 103.100 136.505 104.765 136.675 ;
        RECT 103.120 135.935 103.495 136.335 ;
        RECT 103.665 136.155 103.835 136.505 ;
        RECT 104.005 135.935 104.335 136.335 ;
        RECT 104.505 136.105 104.765 136.505 ;
        RECT 104.945 136.335 105.275 136.755 ;
        RECT 105.445 135.935 105.705 136.755 ;
        RECT 105.875 136.575 107.560 136.755 ;
        RECT 107.730 136.585 109.760 136.755 ;
        RECT 106.050 135.935 106.220 136.405 ;
        RECT 106.390 136.115 106.720 136.575 ;
        RECT 106.890 135.935 107.060 136.405 ;
        RECT 107.230 136.105 107.560 136.575 ;
        RECT 108.205 136.495 109.760 136.585 ;
        RECT 109.930 136.585 111.940 136.755 ;
        RECT 107.730 135.935 107.900 136.405 ;
        RECT 109.930 136.325 110.260 136.585 ;
        RECT 110.770 136.575 111.940 136.585 ;
        RECT 108.170 136.105 110.260 136.325 ;
        RECT 110.430 135.935 110.600 136.405 ;
        RECT 110.770 136.105 111.100 136.575 ;
        RECT 111.270 135.935 111.440 136.405 ;
        RECT 111.610 136.105 111.940 136.575 ;
        RECT 112.315 136.610 112.485 137.345 ;
        RECT 112.760 137.175 112.930 137.345 ;
        RECT 113.975 137.265 114.625 137.435 ;
        RECT 114.795 137.375 115.380 137.545 ;
        RECT 112.655 136.845 112.930 137.175 ;
        RECT 113.100 136.845 113.755 137.175 ;
        RECT 113.975 136.845 114.145 137.265 ;
        RECT 114.795 137.095 114.965 137.375 ;
        RECT 114.540 136.925 114.965 137.095 ;
        RECT 112.760 136.675 112.930 136.845 ;
        RECT 114.795 136.675 114.965 136.925 ;
        RECT 115.135 136.845 115.425 137.175 ;
        RECT 115.595 136.845 115.945 137.545 ;
        RECT 116.115 136.675 116.285 137.715 ;
        RECT 116.525 137.515 116.885 137.690 ;
        RECT 117.470 137.685 117.640 138.485 ;
        RECT 117.810 137.855 118.140 138.315 ;
        RECT 118.310 138.025 118.480 138.485 ;
        RECT 117.810 137.685 118.585 137.855 ;
        RECT 116.525 137.345 117.985 137.515 ;
        RECT 116.520 136.785 116.715 137.175 ;
        RECT 112.315 136.265 112.590 136.610 ;
        RECT 112.760 136.505 114.355 136.675 ;
        RECT 114.795 136.505 115.295 136.675 ;
        RECT 112.780 135.935 113.160 136.335 ;
        RECT 113.330 136.155 113.500 136.505 ;
        RECT 113.670 135.935 114.000 136.335 ;
        RECT 114.185 136.155 114.355 136.505 ;
        RECT 114.525 135.935 114.900 136.335 ;
        RECT 115.125 136.300 115.295 136.505 ;
        RECT 115.545 135.935 115.715 136.675 ;
        RECT 115.970 136.300 116.285 136.675 ;
        RECT 116.515 136.615 116.715 136.785 ;
        RECT 116.885 136.445 117.065 137.345 ;
        RECT 117.235 136.615 117.645 137.175 ;
        RECT 117.815 136.845 117.985 137.345 ;
        RECT 118.155 136.675 118.585 137.685 ;
        RECT 118.755 137.320 119.045 138.485 ;
        RECT 119.225 137.535 119.500 138.305 ;
        RECT 119.670 137.875 120.000 138.305 ;
        RECT 120.170 138.045 120.365 138.485 ;
        RECT 120.545 137.875 120.875 138.305 ;
        RECT 119.670 137.705 120.875 137.875 ;
        RECT 119.225 137.345 119.810 137.535 ;
        RECT 119.980 137.375 120.875 137.705 ;
        RECT 122.065 137.865 122.235 138.295 ;
        RECT 122.405 138.035 122.735 138.485 ;
        RECT 122.065 137.635 122.740 137.865 ;
        RECT 117.890 136.505 118.585 136.675 ;
        RECT 116.475 135.935 116.715 136.445 ;
        RECT 116.885 136.105 117.175 136.445 ;
        RECT 117.405 135.935 117.720 136.445 ;
        RECT 117.890 136.235 118.060 136.505 ;
        RECT 118.230 135.935 118.560 136.335 ;
        RECT 118.755 135.935 119.045 136.660 ;
        RECT 119.225 136.525 119.465 137.175 ;
        RECT 119.635 136.675 119.810 137.345 ;
        RECT 119.980 136.845 120.395 137.175 ;
        RECT 120.575 136.845 120.870 137.175 ;
        RECT 119.635 136.495 119.965 136.675 ;
        RECT 119.240 135.935 119.570 136.325 ;
        RECT 119.740 136.115 119.965 136.495 ;
        RECT 120.165 136.225 120.395 136.845 ;
        RECT 120.575 135.935 120.875 136.665 ;
        RECT 122.035 136.615 122.335 137.465 ;
        RECT 122.505 136.985 122.740 137.635 ;
        RECT 122.910 137.325 123.195 138.270 ;
        RECT 123.375 138.015 124.060 138.485 ;
        RECT 123.370 137.495 124.065 137.805 ;
        RECT 124.240 137.430 124.545 138.215 ;
        RECT 122.910 137.175 123.770 137.325 ;
        RECT 124.335 137.295 124.545 137.430 ;
        RECT 122.910 137.155 124.195 137.175 ;
        RECT 122.505 136.655 123.040 136.985 ;
        RECT 123.210 136.795 124.195 137.155 ;
        RECT 122.505 136.505 122.725 136.655 ;
        RECT 121.980 135.935 122.315 136.440 ;
        RECT 122.485 136.130 122.725 136.505 ;
        RECT 123.210 136.460 123.380 136.795 ;
        RECT 124.370 136.625 124.545 137.295 ;
        RECT 123.005 136.265 123.380 136.460 ;
        RECT 123.005 136.120 123.175 136.265 ;
        RECT 123.740 135.935 124.135 136.430 ;
        RECT 124.305 136.105 124.545 136.625 ;
        RECT 124.735 137.345 125.005 138.315 ;
        RECT 125.215 137.685 125.495 138.485 ;
        RECT 125.675 137.935 126.870 138.265 ;
        RECT 126.000 137.515 126.420 137.765 ;
        RECT 125.175 137.345 126.420 137.515 ;
        RECT 124.735 136.610 124.905 137.345 ;
        RECT 125.175 137.175 125.345 137.345 ;
        RECT 126.645 137.175 126.815 137.735 ;
        RECT 127.065 137.345 127.320 138.485 ;
        RECT 127.510 137.635 128.235 138.305 ;
        RECT 125.115 136.845 125.345 137.175 ;
        RECT 126.075 136.845 126.815 137.175 ;
        RECT 126.985 136.925 127.320 137.175 ;
        RECT 125.175 136.675 125.345 136.845 ;
        RECT 126.565 136.755 126.815 136.845 ;
        RECT 124.735 136.265 125.005 136.610 ;
        RECT 125.175 136.505 125.915 136.675 ;
        RECT 126.565 136.585 127.300 136.755 ;
        RECT 125.195 135.935 125.575 136.335 ;
        RECT 125.745 136.155 125.915 136.505 ;
        RECT 126.085 135.935 126.820 136.415 ;
        RECT 126.990 136.115 127.300 136.585 ;
        RECT 127.510 136.665 127.725 137.635 ;
        RECT 127.935 136.845 128.235 137.465 ;
        RECT 128.415 137.175 128.645 138.305 ;
        RECT 128.815 137.575 129.000 138.305 ;
        RECT 129.170 137.755 129.500 138.485 ;
        RECT 129.670 137.575 129.920 138.305 ;
        RECT 128.815 137.375 129.920 137.575 ;
        RECT 130.255 137.395 131.925 138.485 ;
        RECT 128.415 136.845 128.745 137.175 ;
        RECT 128.925 136.845 129.565 137.175 ;
        RECT 127.510 136.475 128.990 136.665 ;
        RECT 127.890 136.115 128.115 136.475 ;
        RECT 128.295 135.935 128.625 136.305 ;
        RECT 128.805 136.115 128.990 136.475 ;
        RECT 129.315 136.115 129.565 136.845 ;
        RECT 129.735 136.615 130.075 137.175 ;
        RECT 130.255 136.705 131.005 137.225 ;
        RECT 131.175 136.875 131.925 137.395 ;
        RECT 129.745 135.935 130.085 136.445 ;
        RECT 130.255 135.935 131.925 136.705 ;
        RECT 132.105 136.115 132.365 138.305 ;
        RECT 132.535 137.755 132.875 138.485 ;
        RECT 133.055 137.575 133.325 138.305 ;
        RECT 132.555 137.355 133.325 137.575 ;
        RECT 133.505 137.595 133.735 138.305 ;
        RECT 133.905 137.775 134.235 138.485 ;
        RECT 134.405 137.595 134.665 138.305 ;
        RECT 133.505 137.355 134.665 137.595 ;
        RECT 134.855 137.475 135.115 138.485 ;
        RECT 135.285 137.645 135.560 138.315 ;
        RECT 132.555 136.685 132.845 137.355 ;
        RECT 135.285 137.295 135.455 137.645 ;
        RECT 135.760 137.640 135.975 138.485 ;
        RECT 136.160 137.975 136.635 138.315 ;
        RECT 136.815 137.980 137.445 138.485 ;
        RECT 136.815 137.805 137.005 137.980 ;
        RECT 136.200 137.445 136.450 137.740 ;
        RECT 136.675 137.615 137.005 137.805 ;
        RECT 137.175 137.445 137.430 137.810 ;
        RECT 133.025 136.865 133.490 137.175 ;
        RECT 133.670 136.865 134.195 137.175 ;
        RECT 132.555 136.485 133.785 136.685 ;
        RECT 132.625 135.935 133.295 136.305 ;
        RECT 133.475 136.115 133.785 136.485 ;
        RECT 133.965 136.225 134.195 136.865 ;
        RECT 134.375 136.845 134.675 137.175 ;
        RECT 134.855 136.775 135.470 137.295 ;
        RECT 135.640 137.275 137.430 137.445 ;
        RECT 137.615 137.345 137.905 138.485 ;
        RECT 138.075 137.765 138.525 138.315 ;
        RECT 138.715 137.765 139.045 138.485 ;
        RECT 135.640 136.845 135.870 137.275 ;
        RECT 134.375 135.935 134.665 136.665 ;
        RECT 134.855 135.935 135.130 136.595 ;
        RECT 135.300 136.565 135.470 136.775 ;
        RECT 136.055 136.600 136.465 137.095 ;
        RECT 135.300 136.105 135.550 136.565 ;
        RECT 135.725 135.935 136.055 136.430 ;
        RECT 136.235 136.155 136.465 136.600 ;
        RECT 136.635 136.420 136.890 137.275 ;
        RECT 137.060 136.615 137.445 137.095 ;
        RECT 136.635 136.155 137.425 136.420 ;
        RECT 137.615 135.935 137.905 136.735 ;
        RECT 138.075 136.395 138.325 137.765 ;
        RECT 139.255 137.595 139.555 138.145 ;
        RECT 139.725 137.815 140.005 138.485 ;
        RECT 140.415 138.145 141.555 138.315 ;
        RECT 140.415 137.685 140.715 138.145 ;
        RECT 138.615 137.425 139.555 137.595 ;
        RECT 138.615 137.175 138.785 137.425 ;
        RECT 139.890 137.175 140.205 137.615 ;
        RECT 140.885 137.515 141.215 137.975 ;
        RECT 138.495 136.845 138.785 137.175 ;
        RECT 138.955 136.925 139.285 137.175 ;
        RECT 139.515 136.925 140.205 137.175 ;
        RECT 140.455 137.295 141.215 137.515 ;
        RECT 141.385 137.515 141.555 138.145 ;
        RECT 141.725 137.685 142.055 138.485 ;
        RECT 142.225 137.515 142.500 138.315 ;
        RECT 141.385 137.305 142.500 137.515 ;
        RECT 142.675 137.395 144.345 138.485 ;
        RECT 138.615 136.755 138.785 136.845 ;
        RECT 140.455 136.785 140.670 137.295 ;
        RECT 140.840 136.925 141.610 137.125 ;
        RECT 141.780 136.925 142.500 137.125 ;
        RECT 140.435 136.755 140.670 136.785 ;
        RECT 138.615 136.565 140.005 136.755 ;
        RECT 140.435 136.615 142.055 136.755 ;
        RECT 140.455 136.585 142.055 136.615 ;
        RECT 138.075 136.105 138.625 136.395 ;
        RECT 138.795 135.935 139.045 136.395 ;
        RECT 139.675 136.205 140.005 136.565 ;
        RECT 140.885 136.575 142.055 136.585 ;
        RECT 140.425 135.935 140.715 136.405 ;
        RECT 140.885 136.105 141.215 136.575 ;
        RECT 141.385 135.935 141.555 136.405 ;
        RECT 141.725 136.105 142.055 136.575 ;
        RECT 142.225 135.935 142.500 136.755 ;
        RECT 142.675 136.705 143.425 137.225 ;
        RECT 143.595 136.875 144.345 137.395 ;
        RECT 144.515 137.320 144.805 138.485 ;
        RECT 145.010 137.695 145.545 138.315 ;
        RECT 142.675 135.935 144.345 136.705 ;
        RECT 145.010 136.675 145.325 137.695 ;
        RECT 145.715 137.685 146.045 138.485 ;
        RECT 146.530 137.515 146.920 137.690 ;
        RECT 145.495 137.345 146.920 137.515 ;
        RECT 147.365 137.555 147.535 138.315 ;
        RECT 147.750 137.725 148.080 138.485 ;
        RECT 147.365 137.385 148.080 137.555 ;
        RECT 148.250 137.410 148.505 138.315 ;
        RECT 145.495 136.845 145.665 137.345 ;
        RECT 144.515 135.935 144.805 136.660 ;
        RECT 145.010 136.105 145.625 136.675 ;
        RECT 145.915 136.615 146.180 137.175 ;
        RECT 146.350 136.445 146.520 137.345 ;
        RECT 146.690 136.615 147.045 137.175 ;
        RECT 147.275 136.835 147.630 137.205 ;
        RECT 147.910 137.175 148.080 137.385 ;
        RECT 147.910 136.845 148.165 137.175 ;
        RECT 147.910 136.655 148.080 136.845 ;
        RECT 148.335 136.680 148.505 137.410 ;
        RECT 148.680 137.335 148.940 138.485 ;
        RECT 149.115 138.050 154.460 138.485 ;
        RECT 147.365 136.485 148.080 136.655 ;
        RECT 145.795 135.935 146.010 136.445 ;
        RECT 146.240 136.115 146.520 136.445 ;
        RECT 146.700 135.935 146.940 136.445 ;
        RECT 147.365 136.105 147.535 136.485 ;
        RECT 147.750 135.935 148.080 136.315 ;
        RECT 148.250 136.105 148.505 136.680 ;
        RECT 148.680 135.935 148.940 136.775 ;
        RECT 150.700 136.480 151.040 137.310 ;
        RECT 152.520 136.800 152.870 138.050 ;
        RECT 154.635 137.395 156.305 138.485 ;
        RECT 154.635 136.705 155.385 137.225 ;
        RECT 155.555 136.875 156.305 137.395 ;
        RECT 156.935 137.395 158.145 138.485 ;
        RECT 156.935 136.855 157.455 137.395 ;
        RECT 149.115 135.935 154.460 136.480 ;
        RECT 154.635 135.935 156.305 136.705 ;
        RECT 157.625 136.685 158.145 137.225 ;
        RECT 156.935 135.935 158.145 136.685 ;
        RECT 2.750 135.765 158.230 135.935 ;
        RECT 2.835 135.015 4.045 135.765 ;
        RECT 4.765 135.215 4.935 135.595 ;
        RECT 5.115 135.385 5.445 135.765 ;
        RECT 4.765 135.045 5.430 135.215 ;
        RECT 5.625 135.090 5.885 135.595 ;
        RECT 2.835 134.475 3.355 135.015 ;
        RECT 3.525 134.305 4.045 134.845 ;
        RECT 4.695 134.495 5.025 134.865 ;
        RECT 5.260 134.790 5.430 135.045 ;
        RECT 5.260 134.460 5.545 134.790 ;
        RECT 5.260 134.315 5.430 134.460 ;
        RECT 2.835 133.215 4.045 134.305 ;
        RECT 4.765 134.145 5.430 134.315 ;
        RECT 5.715 134.290 5.885 135.090 ;
        RECT 4.765 133.385 4.935 134.145 ;
        RECT 5.115 133.215 5.445 133.975 ;
        RECT 5.615 133.385 5.885 134.290 ;
        RECT 6.055 135.090 6.315 135.595 ;
        RECT 6.495 135.385 6.825 135.765 ;
        RECT 7.005 135.215 7.175 135.595 ;
        RECT 6.055 134.290 6.225 135.090 ;
        RECT 6.510 135.045 7.175 135.215 ;
        RECT 6.510 134.790 6.680 135.045 ;
        RECT 8.360 135.025 8.615 135.595 ;
        RECT 8.785 135.365 9.115 135.765 ;
        RECT 9.540 135.230 10.070 135.595 ;
        RECT 10.260 135.425 10.535 135.595 ;
        RECT 10.255 135.255 10.535 135.425 ;
        RECT 9.540 135.195 9.715 135.230 ;
        RECT 8.785 135.025 9.715 135.195 ;
        RECT 6.395 134.460 6.680 134.790 ;
        RECT 6.915 134.495 7.245 134.865 ;
        RECT 6.510 134.315 6.680 134.460 ;
        RECT 8.360 134.355 8.530 135.025 ;
        RECT 8.785 134.855 8.955 135.025 ;
        RECT 8.700 134.525 8.955 134.855 ;
        RECT 9.180 134.525 9.375 134.855 ;
        RECT 6.055 133.385 6.325 134.290 ;
        RECT 6.510 134.145 7.175 134.315 ;
        RECT 6.495 133.215 6.825 133.975 ;
        RECT 7.005 133.385 7.175 134.145 ;
        RECT 8.360 133.385 8.695 134.355 ;
        RECT 8.865 133.215 9.035 134.355 ;
        RECT 9.205 133.555 9.375 134.525 ;
        RECT 9.545 133.895 9.715 135.025 ;
        RECT 9.885 134.235 10.055 135.035 ;
        RECT 10.260 134.435 10.535 135.255 ;
        RECT 10.705 134.235 10.895 135.595 ;
        RECT 11.075 135.230 11.585 135.765 ;
        RECT 11.805 134.955 12.050 135.560 ;
        RECT 12.500 135.215 12.755 135.505 ;
        RECT 12.925 135.385 13.255 135.765 ;
        RECT 12.500 135.045 13.250 135.215 ;
        RECT 11.095 134.785 12.325 134.955 ;
        RECT 9.885 134.065 10.895 134.235 ;
        RECT 11.065 134.220 11.815 134.410 ;
        RECT 9.545 133.725 10.670 133.895 ;
        RECT 11.065 133.555 11.235 134.220 ;
        RECT 11.985 133.975 12.325 134.785 ;
        RECT 12.500 134.225 12.850 134.875 ;
        RECT 13.020 134.055 13.250 135.045 ;
        RECT 9.205 133.385 11.235 133.555 ;
        RECT 11.405 133.215 11.575 133.975 ;
        RECT 11.810 133.565 12.325 133.975 ;
        RECT 12.500 133.885 13.250 134.055 ;
        RECT 12.500 133.385 12.755 133.885 ;
        RECT 12.925 133.215 13.255 133.715 ;
        RECT 13.425 133.385 13.595 135.505 ;
        RECT 13.955 135.405 14.285 135.765 ;
        RECT 14.455 135.375 14.950 135.545 ;
        RECT 15.155 135.375 16.010 135.545 ;
        RECT 13.825 134.185 14.285 135.235 ;
        RECT 13.765 133.400 14.090 134.185 ;
        RECT 14.455 134.015 14.625 135.375 ;
        RECT 14.795 134.465 15.145 135.085 ;
        RECT 15.315 134.865 15.670 135.085 ;
        RECT 15.315 134.275 15.485 134.865 ;
        RECT 15.840 134.665 16.010 135.375 ;
        RECT 16.885 135.305 17.215 135.765 ;
        RECT 17.425 135.405 17.775 135.575 ;
        RECT 16.215 134.835 17.005 135.085 ;
        RECT 17.425 135.015 17.685 135.405 ;
        RECT 17.995 135.315 18.945 135.595 ;
        RECT 19.115 135.325 19.305 135.765 ;
        RECT 19.475 135.385 20.545 135.555 ;
        RECT 17.175 134.665 17.345 134.845 ;
        RECT 14.455 133.845 14.850 134.015 ;
        RECT 15.020 133.885 15.485 134.275 ;
        RECT 15.655 134.495 17.345 134.665 ;
        RECT 14.680 133.715 14.850 133.845 ;
        RECT 15.655 133.715 15.825 134.495 ;
        RECT 17.515 134.325 17.685 135.015 ;
        RECT 16.185 134.155 17.685 134.325 ;
        RECT 17.875 134.355 18.085 135.145 ;
        RECT 18.255 134.525 18.605 135.145 ;
        RECT 18.775 134.535 18.945 135.315 ;
        RECT 19.475 135.155 19.645 135.385 ;
        RECT 19.115 134.985 19.645 135.155 ;
        RECT 19.115 134.705 19.335 134.985 ;
        RECT 19.815 134.815 20.055 135.215 ;
        RECT 18.775 134.365 19.180 134.535 ;
        RECT 19.515 134.445 20.055 134.815 ;
        RECT 20.225 135.030 20.545 135.385 ;
        RECT 20.790 135.305 21.095 135.765 ;
        RECT 21.265 135.055 21.520 135.585 ;
        RECT 20.225 134.855 20.550 135.030 ;
        RECT 20.225 134.555 21.140 134.855 ;
        RECT 20.400 134.525 21.140 134.555 ;
        RECT 17.875 134.195 18.550 134.355 ;
        RECT 19.010 134.275 19.180 134.365 ;
        RECT 17.875 134.185 18.840 134.195 ;
        RECT 17.515 134.015 17.685 134.155 ;
        RECT 14.260 133.215 14.510 133.675 ;
        RECT 14.680 133.385 14.930 133.715 ;
        RECT 15.145 133.385 15.825 133.715 ;
        RECT 15.995 133.815 17.070 133.985 ;
        RECT 17.515 133.845 18.075 134.015 ;
        RECT 18.380 133.895 18.840 134.185 ;
        RECT 19.010 134.105 20.230 134.275 ;
        RECT 15.995 133.475 16.165 133.815 ;
        RECT 16.400 133.215 16.730 133.645 ;
        RECT 16.900 133.475 17.070 133.815 ;
        RECT 17.365 133.215 17.735 133.675 ;
        RECT 17.905 133.385 18.075 133.845 ;
        RECT 19.010 133.725 19.180 134.105 ;
        RECT 20.400 133.935 20.570 134.525 ;
        RECT 21.310 134.405 21.520 135.055 ;
        RECT 21.695 135.015 22.905 135.765 ;
        RECT 23.165 135.215 23.335 135.595 ;
        RECT 23.515 135.385 23.845 135.765 ;
        RECT 23.165 135.045 23.830 135.215 ;
        RECT 24.025 135.090 24.285 135.595 ;
        RECT 21.695 134.475 22.215 135.015 ;
        RECT 18.310 133.385 19.180 133.725 ;
        RECT 19.770 133.765 20.570 133.935 ;
        RECT 19.350 133.215 19.600 133.675 ;
        RECT 19.770 133.475 19.940 133.765 ;
        RECT 20.120 133.215 20.450 133.595 ;
        RECT 20.790 133.215 21.095 134.355 ;
        RECT 21.265 133.525 21.520 134.405 ;
        RECT 22.385 134.305 22.905 134.845 ;
        RECT 23.095 134.495 23.425 134.865 ;
        RECT 23.660 134.790 23.830 135.045 ;
        RECT 23.660 134.460 23.945 134.790 ;
        RECT 23.660 134.315 23.830 134.460 ;
        RECT 21.695 133.215 22.905 134.305 ;
        RECT 23.165 134.145 23.830 134.315 ;
        RECT 24.115 134.290 24.285 135.090 ;
        RECT 23.165 133.385 23.335 134.145 ;
        RECT 23.515 133.215 23.845 133.975 ;
        RECT 24.015 133.385 24.285 134.290 ;
        RECT 24.460 135.025 24.715 135.595 ;
        RECT 24.885 135.365 25.215 135.765 ;
        RECT 25.640 135.230 26.170 135.595 ;
        RECT 26.360 135.425 26.635 135.595 ;
        RECT 26.355 135.255 26.635 135.425 ;
        RECT 25.640 135.195 25.815 135.230 ;
        RECT 24.885 135.025 25.815 135.195 ;
        RECT 24.460 134.355 24.630 135.025 ;
        RECT 24.885 134.855 25.055 135.025 ;
        RECT 24.800 134.525 25.055 134.855 ;
        RECT 25.280 134.525 25.475 134.855 ;
        RECT 24.460 133.385 24.795 134.355 ;
        RECT 24.965 133.215 25.135 134.355 ;
        RECT 25.305 133.555 25.475 134.525 ;
        RECT 25.645 133.895 25.815 135.025 ;
        RECT 25.985 134.235 26.155 135.035 ;
        RECT 26.360 134.435 26.635 135.255 ;
        RECT 26.805 134.235 26.995 135.595 ;
        RECT 27.175 135.230 27.685 135.765 ;
        RECT 27.905 134.955 28.150 135.560 ;
        RECT 28.595 135.040 28.885 135.765 ;
        RECT 29.115 135.285 29.395 135.765 ;
        RECT 29.565 135.115 29.825 135.505 ;
        RECT 30.000 135.285 30.255 135.765 ;
        RECT 30.425 135.115 30.720 135.505 ;
        RECT 30.900 135.285 31.175 135.765 ;
        RECT 31.345 135.265 31.645 135.595 ;
        RECT 27.195 134.785 28.425 134.955 ;
        RECT 25.985 134.065 26.995 134.235 ;
        RECT 27.165 134.220 27.915 134.410 ;
        RECT 25.645 133.725 26.770 133.895 ;
        RECT 27.165 133.555 27.335 134.220 ;
        RECT 28.085 133.975 28.425 134.785 ;
        RECT 29.070 134.945 30.720 135.115 ;
        RECT 29.070 134.435 29.475 134.945 ;
        RECT 29.645 134.605 30.785 134.775 ;
        RECT 25.305 133.385 27.335 133.555 ;
        RECT 27.505 133.215 27.675 133.975 ;
        RECT 27.910 133.565 28.425 133.975 ;
        RECT 28.595 133.215 28.885 134.380 ;
        RECT 29.070 134.265 29.825 134.435 ;
        RECT 29.110 133.215 29.395 134.085 ;
        RECT 29.565 134.015 29.825 134.265 ;
        RECT 30.615 134.355 30.785 134.605 ;
        RECT 30.955 134.525 31.305 135.095 ;
        RECT 31.475 134.355 31.645 135.265 ;
        RECT 31.820 135.215 32.075 135.505 ;
        RECT 32.245 135.385 32.575 135.765 ;
        RECT 31.820 135.045 32.570 135.215 ;
        RECT 30.615 134.185 31.645 134.355 ;
        RECT 31.820 134.225 32.170 134.875 ;
        RECT 29.565 133.845 30.685 134.015 ;
        RECT 29.565 133.385 29.825 133.845 ;
        RECT 30.000 133.215 30.255 133.675 ;
        RECT 30.425 133.385 30.685 133.845 ;
        RECT 30.855 133.215 31.165 134.015 ;
        RECT 31.335 133.385 31.645 134.185 ;
        RECT 32.340 134.055 32.570 135.045 ;
        RECT 31.820 133.885 32.570 134.055 ;
        RECT 31.820 133.385 32.075 133.885 ;
        RECT 32.245 133.215 32.575 133.715 ;
        RECT 32.745 133.385 32.915 135.505 ;
        RECT 33.275 135.405 33.605 135.765 ;
        RECT 33.775 135.375 34.270 135.545 ;
        RECT 34.475 135.375 35.330 135.545 ;
        RECT 33.145 134.185 33.605 135.235 ;
        RECT 33.085 133.400 33.410 134.185 ;
        RECT 33.775 134.015 33.945 135.375 ;
        RECT 34.115 134.465 34.465 135.085 ;
        RECT 34.635 134.865 34.990 135.085 ;
        RECT 34.635 134.275 34.805 134.865 ;
        RECT 35.160 134.665 35.330 135.375 ;
        RECT 36.205 135.305 36.535 135.765 ;
        RECT 36.745 135.405 37.095 135.575 ;
        RECT 35.535 134.835 36.325 135.085 ;
        RECT 36.745 135.015 37.005 135.405 ;
        RECT 37.315 135.315 38.265 135.595 ;
        RECT 38.435 135.325 38.625 135.765 ;
        RECT 38.795 135.385 39.865 135.555 ;
        RECT 36.495 134.665 36.665 134.845 ;
        RECT 33.775 133.845 34.170 134.015 ;
        RECT 34.340 133.885 34.805 134.275 ;
        RECT 34.975 134.495 36.665 134.665 ;
        RECT 34.000 133.715 34.170 133.845 ;
        RECT 34.975 133.715 35.145 134.495 ;
        RECT 36.835 134.325 37.005 135.015 ;
        RECT 35.505 134.155 37.005 134.325 ;
        RECT 37.195 134.355 37.405 135.145 ;
        RECT 37.575 134.525 37.925 135.145 ;
        RECT 38.095 134.535 38.265 135.315 ;
        RECT 38.795 135.155 38.965 135.385 ;
        RECT 38.435 134.985 38.965 135.155 ;
        RECT 38.435 134.705 38.655 134.985 ;
        RECT 39.135 134.815 39.375 135.215 ;
        RECT 38.095 134.365 38.500 134.535 ;
        RECT 38.835 134.445 39.375 134.815 ;
        RECT 39.545 135.030 39.865 135.385 ;
        RECT 40.110 135.305 40.415 135.765 ;
        RECT 40.585 135.055 40.840 135.585 ;
        RECT 39.545 134.855 39.870 135.030 ;
        RECT 39.545 134.555 40.460 134.855 ;
        RECT 39.720 134.525 40.460 134.555 ;
        RECT 37.195 134.195 37.870 134.355 ;
        RECT 38.330 134.275 38.500 134.365 ;
        RECT 37.195 134.185 38.160 134.195 ;
        RECT 36.835 134.015 37.005 134.155 ;
        RECT 33.580 133.215 33.830 133.675 ;
        RECT 34.000 133.385 34.250 133.715 ;
        RECT 34.465 133.385 35.145 133.715 ;
        RECT 35.315 133.815 36.390 133.985 ;
        RECT 36.835 133.845 37.395 134.015 ;
        RECT 37.700 133.895 38.160 134.185 ;
        RECT 38.330 134.105 39.550 134.275 ;
        RECT 35.315 133.475 35.485 133.815 ;
        RECT 35.720 133.215 36.050 133.645 ;
        RECT 36.220 133.475 36.390 133.815 ;
        RECT 36.685 133.215 37.055 133.675 ;
        RECT 37.225 133.385 37.395 133.845 ;
        RECT 38.330 133.725 38.500 134.105 ;
        RECT 39.720 133.935 39.890 134.525 ;
        RECT 40.630 134.405 40.840 135.055 ;
        RECT 37.630 133.385 38.500 133.725 ;
        RECT 39.090 133.765 39.890 133.935 ;
        RECT 38.670 133.215 38.920 133.675 ;
        RECT 39.090 133.475 39.260 133.765 ;
        RECT 39.440 133.215 39.770 133.595 ;
        RECT 40.110 133.215 40.415 134.355 ;
        RECT 40.585 133.525 40.840 134.405 ;
        RECT 41.940 135.055 42.195 135.585 ;
        RECT 42.365 135.305 42.670 135.765 ;
        RECT 42.915 135.385 43.985 135.555 ;
        RECT 41.940 134.405 42.150 135.055 ;
        RECT 42.915 135.030 43.235 135.385 ;
        RECT 42.910 134.855 43.235 135.030 ;
        RECT 42.320 134.555 43.235 134.855 ;
        RECT 43.405 134.815 43.645 135.215 ;
        RECT 43.815 135.155 43.985 135.385 ;
        RECT 44.155 135.325 44.345 135.765 ;
        RECT 44.515 135.315 45.465 135.595 ;
        RECT 45.685 135.405 46.035 135.575 ;
        RECT 43.815 134.985 44.345 135.155 ;
        RECT 42.320 134.525 43.060 134.555 ;
        RECT 41.940 133.525 42.195 134.405 ;
        RECT 42.365 133.215 42.670 134.355 ;
        RECT 42.890 133.935 43.060 134.525 ;
        RECT 43.405 134.445 43.945 134.815 ;
        RECT 44.125 134.705 44.345 134.985 ;
        RECT 44.515 134.535 44.685 135.315 ;
        RECT 44.280 134.365 44.685 134.535 ;
        RECT 44.855 134.525 45.205 135.145 ;
        RECT 44.280 134.275 44.450 134.365 ;
        RECT 45.375 134.355 45.585 135.145 ;
        RECT 43.230 134.105 44.450 134.275 ;
        RECT 44.910 134.195 45.585 134.355 ;
        RECT 42.890 133.765 43.690 133.935 ;
        RECT 43.010 133.215 43.340 133.595 ;
        RECT 43.520 133.475 43.690 133.765 ;
        RECT 44.280 133.725 44.450 134.105 ;
        RECT 44.620 134.185 45.585 134.195 ;
        RECT 45.775 135.015 46.035 135.405 ;
        RECT 46.245 135.305 46.575 135.765 ;
        RECT 47.450 135.375 48.305 135.545 ;
        RECT 48.510 135.375 49.005 135.545 ;
        RECT 49.175 135.405 49.505 135.765 ;
        RECT 45.775 134.325 45.945 135.015 ;
        RECT 46.115 134.665 46.285 134.845 ;
        RECT 46.455 134.835 47.245 135.085 ;
        RECT 47.450 134.665 47.620 135.375 ;
        RECT 47.790 134.865 48.145 135.085 ;
        RECT 46.115 134.495 47.805 134.665 ;
        RECT 44.620 133.895 45.080 134.185 ;
        RECT 45.775 134.155 47.275 134.325 ;
        RECT 45.775 134.015 45.945 134.155 ;
        RECT 45.385 133.845 45.945 134.015 ;
        RECT 43.860 133.215 44.110 133.675 ;
        RECT 44.280 133.385 45.150 133.725 ;
        RECT 45.385 133.385 45.555 133.845 ;
        RECT 46.390 133.815 47.465 133.985 ;
        RECT 45.725 133.215 46.095 133.675 ;
        RECT 46.390 133.475 46.560 133.815 ;
        RECT 46.730 133.215 47.060 133.645 ;
        RECT 47.295 133.475 47.465 133.815 ;
        RECT 47.635 133.715 47.805 134.495 ;
        RECT 47.975 134.275 48.145 134.865 ;
        RECT 48.315 134.465 48.665 135.085 ;
        RECT 47.975 133.885 48.440 134.275 ;
        RECT 48.835 134.015 49.005 135.375 ;
        RECT 49.175 134.185 49.635 135.235 ;
        RECT 48.610 133.845 49.005 134.015 ;
        RECT 48.610 133.715 48.780 133.845 ;
        RECT 47.635 133.385 48.315 133.715 ;
        RECT 48.530 133.385 48.780 133.715 ;
        RECT 48.950 133.215 49.200 133.675 ;
        RECT 49.370 133.400 49.695 134.185 ;
        RECT 49.865 133.385 50.035 135.505 ;
        RECT 50.205 135.385 50.535 135.765 ;
        RECT 50.705 135.215 50.960 135.505 ;
        RECT 50.210 135.045 50.960 135.215 ;
        RECT 51.135 135.090 51.395 135.595 ;
        RECT 51.575 135.385 51.905 135.765 ;
        RECT 52.085 135.215 52.255 135.595 ;
        RECT 50.210 134.055 50.440 135.045 ;
        RECT 50.610 134.225 50.960 134.875 ;
        RECT 51.135 134.290 51.305 135.090 ;
        RECT 51.590 135.045 52.255 135.215 ;
        RECT 52.605 135.215 52.775 135.595 ;
        RECT 52.955 135.385 53.285 135.765 ;
        RECT 52.605 135.045 53.270 135.215 ;
        RECT 53.465 135.090 53.725 135.595 ;
        RECT 51.590 134.790 51.760 135.045 ;
        RECT 51.475 134.460 51.760 134.790 ;
        RECT 51.995 134.495 52.325 134.865 ;
        RECT 52.535 134.495 52.865 134.865 ;
        RECT 53.100 134.790 53.270 135.045 ;
        RECT 51.590 134.315 51.760 134.460 ;
        RECT 53.100 134.460 53.385 134.790 ;
        RECT 53.100 134.315 53.270 134.460 ;
        RECT 50.210 133.885 50.960 134.055 ;
        RECT 50.205 133.215 50.535 133.715 ;
        RECT 50.705 133.385 50.960 133.885 ;
        RECT 51.135 133.385 51.405 134.290 ;
        RECT 51.590 134.145 52.255 134.315 ;
        RECT 51.575 133.215 51.905 133.975 ;
        RECT 52.085 133.385 52.255 134.145 ;
        RECT 52.605 134.145 53.270 134.315 ;
        RECT 53.555 134.290 53.725 135.090 ;
        RECT 54.355 135.040 54.645 135.765 ;
        RECT 54.905 135.215 55.075 135.595 ;
        RECT 55.255 135.385 55.585 135.765 ;
        RECT 54.905 135.045 55.570 135.215 ;
        RECT 55.765 135.090 56.025 135.595 ;
        RECT 54.835 134.495 55.165 134.865 ;
        RECT 55.400 134.790 55.570 135.045 ;
        RECT 55.400 134.460 55.685 134.790 ;
        RECT 52.605 133.385 52.775 134.145 ;
        RECT 52.955 133.215 53.285 133.975 ;
        RECT 53.455 133.385 53.725 134.290 ;
        RECT 54.355 133.215 54.645 134.380 ;
        RECT 55.400 134.315 55.570 134.460 ;
        RECT 54.905 134.145 55.570 134.315 ;
        RECT 55.855 134.290 56.025 135.090 ;
        RECT 56.200 135.215 56.455 135.505 ;
        RECT 56.625 135.385 56.955 135.765 ;
        RECT 56.200 135.045 56.950 135.215 ;
        RECT 54.905 133.385 55.075 134.145 ;
        RECT 55.255 133.215 55.585 133.975 ;
        RECT 55.755 133.385 56.025 134.290 ;
        RECT 56.200 134.225 56.550 134.875 ;
        RECT 56.720 134.055 56.950 135.045 ;
        RECT 56.200 133.885 56.950 134.055 ;
        RECT 56.200 133.385 56.455 133.885 ;
        RECT 56.625 133.215 56.955 133.715 ;
        RECT 57.125 133.385 57.295 135.505 ;
        RECT 57.655 135.405 57.985 135.765 ;
        RECT 58.155 135.375 58.650 135.545 ;
        RECT 58.855 135.375 59.710 135.545 ;
        RECT 57.525 134.185 57.985 135.235 ;
        RECT 57.465 133.400 57.790 134.185 ;
        RECT 58.155 134.015 58.325 135.375 ;
        RECT 58.495 134.465 58.845 135.085 ;
        RECT 59.015 134.865 59.370 135.085 ;
        RECT 59.015 134.275 59.185 134.865 ;
        RECT 59.540 134.665 59.710 135.375 ;
        RECT 60.585 135.305 60.915 135.765 ;
        RECT 61.125 135.405 61.475 135.575 ;
        RECT 59.915 134.835 60.705 135.085 ;
        RECT 61.125 135.015 61.385 135.405 ;
        RECT 61.695 135.315 62.645 135.595 ;
        RECT 62.815 135.325 63.005 135.765 ;
        RECT 63.175 135.385 64.245 135.555 ;
        RECT 60.875 134.665 61.045 134.845 ;
        RECT 58.155 133.845 58.550 134.015 ;
        RECT 58.720 133.885 59.185 134.275 ;
        RECT 59.355 134.495 61.045 134.665 ;
        RECT 58.380 133.715 58.550 133.845 ;
        RECT 59.355 133.715 59.525 134.495 ;
        RECT 61.215 134.325 61.385 135.015 ;
        RECT 59.885 134.155 61.385 134.325 ;
        RECT 61.575 134.355 61.785 135.145 ;
        RECT 61.955 134.525 62.305 135.145 ;
        RECT 62.475 134.535 62.645 135.315 ;
        RECT 63.175 135.155 63.345 135.385 ;
        RECT 62.815 134.985 63.345 135.155 ;
        RECT 62.815 134.705 63.035 134.985 ;
        RECT 63.515 134.815 63.755 135.215 ;
        RECT 62.475 134.365 62.880 134.535 ;
        RECT 63.215 134.445 63.755 134.815 ;
        RECT 63.925 135.030 64.245 135.385 ;
        RECT 64.490 135.305 64.795 135.765 ;
        RECT 64.965 135.055 65.220 135.585 ;
        RECT 63.925 134.855 64.250 135.030 ;
        RECT 63.925 134.555 64.840 134.855 ;
        RECT 64.100 134.525 64.840 134.555 ;
        RECT 61.575 134.195 62.250 134.355 ;
        RECT 62.710 134.275 62.880 134.365 ;
        RECT 61.575 134.185 62.540 134.195 ;
        RECT 61.215 134.015 61.385 134.155 ;
        RECT 57.960 133.215 58.210 133.675 ;
        RECT 58.380 133.385 58.630 133.715 ;
        RECT 58.845 133.385 59.525 133.715 ;
        RECT 59.695 133.815 60.770 133.985 ;
        RECT 61.215 133.845 61.775 134.015 ;
        RECT 62.080 133.895 62.540 134.185 ;
        RECT 62.710 134.105 63.930 134.275 ;
        RECT 59.695 133.475 59.865 133.815 ;
        RECT 60.100 133.215 60.430 133.645 ;
        RECT 60.600 133.475 60.770 133.815 ;
        RECT 61.065 133.215 61.435 133.675 ;
        RECT 61.605 133.385 61.775 133.845 ;
        RECT 62.710 133.725 62.880 134.105 ;
        RECT 64.100 133.935 64.270 134.525 ;
        RECT 65.010 134.405 65.220 135.055 ;
        RECT 62.010 133.385 62.880 133.725 ;
        RECT 63.470 133.765 64.270 133.935 ;
        RECT 63.050 133.215 63.300 133.675 ;
        RECT 63.470 133.475 63.640 133.765 ;
        RECT 63.820 133.215 64.150 133.595 ;
        RECT 64.490 133.215 64.795 134.355 ;
        RECT 64.965 133.525 65.220 134.405 ;
        RECT 65.395 135.090 65.655 135.595 ;
        RECT 65.835 135.385 66.165 135.765 ;
        RECT 66.345 135.215 66.515 135.595 ;
        RECT 65.395 134.290 65.565 135.090 ;
        RECT 65.850 135.045 66.515 135.215 ;
        RECT 65.850 134.790 66.020 135.045 ;
        RECT 66.780 134.965 67.035 135.765 ;
        RECT 67.205 135.100 67.455 135.595 ;
        RECT 67.625 135.385 67.955 135.765 ;
        RECT 68.125 135.385 69.420 135.555 ;
        RECT 68.125 135.215 68.295 135.385 ;
        RECT 65.735 134.460 66.020 134.790 ;
        RECT 66.255 134.495 66.585 134.865 ;
        RECT 65.850 134.315 66.020 134.460 ;
        RECT 65.395 133.385 65.665 134.290 ;
        RECT 65.850 134.145 66.515 134.315 ;
        RECT 65.835 133.215 66.165 133.975 ;
        RECT 66.345 133.385 66.515 134.145 ;
        RECT 66.780 133.215 67.035 134.355 ;
        RECT 67.205 134.255 67.375 135.100 ;
        RECT 67.685 135.045 68.295 135.215 ;
        RECT 69.590 135.115 69.780 135.430 ;
        RECT 70.040 135.265 70.240 135.765 ;
        RECT 67.685 134.855 67.855 135.045 ;
        RECT 67.545 134.525 67.855 134.855 ;
        RECT 67.205 133.385 67.515 134.255 ;
        RECT 67.685 134.015 67.855 134.525 ;
        RECT 68.025 134.355 68.195 134.855 ;
        RECT 68.505 134.570 69.135 135.085 ;
        RECT 69.315 134.825 69.780 135.115 ;
        RECT 68.965 134.535 69.135 134.570 ;
        RECT 68.025 134.185 68.685 134.355 ;
        RECT 68.965 134.225 69.780 134.535 ;
        RECT 70.050 134.225 70.240 135.095 ;
        RECT 68.515 134.015 68.685 134.185 ;
        RECT 70.410 134.015 70.740 135.595 ;
        RECT 70.915 135.015 72.125 135.765 ;
        RECT 70.915 134.475 71.435 135.015 ;
        RECT 72.305 134.955 72.575 135.765 ;
        RECT 72.745 134.955 73.075 135.595 ;
        RECT 73.245 134.955 73.485 135.765 ;
        RECT 73.685 134.955 73.955 135.765 ;
        RECT 74.125 134.955 74.455 135.595 ;
        RECT 74.625 134.955 74.865 135.765 ;
        RECT 71.605 134.305 72.125 134.845 ;
        RECT 72.295 134.525 72.645 134.775 ;
        RECT 72.815 134.355 72.985 134.955 ;
        RECT 73.155 134.525 73.505 134.775 ;
        RECT 73.675 134.525 74.025 134.775 ;
        RECT 74.195 134.355 74.365 134.955 ;
        RECT 74.535 134.525 74.885 134.775 ;
        RECT 67.685 133.845 68.345 134.015 ;
        RECT 68.515 133.845 70.740 134.015 ;
        RECT 67.715 133.215 68.005 133.675 ;
        RECT 68.175 133.595 68.345 133.845 ;
        RECT 68.175 133.425 69.485 133.595 ;
        RECT 70.015 133.215 70.235 133.675 ;
        RECT 70.405 133.385 70.740 133.845 ;
        RECT 70.915 133.215 72.125 134.305 ;
        RECT 72.305 133.215 72.635 134.355 ;
        RECT 72.815 134.185 73.495 134.355 ;
        RECT 73.165 133.400 73.495 134.185 ;
        RECT 73.685 133.215 74.015 134.355 ;
        RECT 74.195 134.185 74.875 134.355 ;
        RECT 74.545 133.400 74.875 134.185 ;
        RECT 75.065 133.395 75.325 135.585 ;
        RECT 75.585 135.395 76.255 135.765 ;
        RECT 76.435 135.215 76.745 135.585 ;
        RECT 75.515 135.015 76.745 135.215 ;
        RECT 75.515 134.345 75.805 135.015 ;
        RECT 76.925 134.835 77.155 135.475 ;
        RECT 77.335 135.035 77.625 135.765 ;
        RECT 77.905 135.215 78.075 135.595 ;
        RECT 78.290 135.385 78.620 135.765 ;
        RECT 77.905 135.045 78.620 135.215 ;
        RECT 75.985 134.525 76.450 134.835 ;
        RECT 76.630 134.525 77.155 134.835 ;
        RECT 77.335 134.525 77.635 134.855 ;
        RECT 77.815 134.495 78.170 134.865 ;
        RECT 78.450 134.855 78.620 135.045 ;
        RECT 78.790 135.020 79.045 135.595 ;
        RECT 78.450 134.525 78.705 134.855 ;
        RECT 75.515 134.125 76.285 134.345 ;
        RECT 75.495 133.215 75.835 133.945 ;
        RECT 76.015 133.395 76.285 134.125 ;
        RECT 76.465 134.105 77.625 134.345 ;
        RECT 78.450 134.315 78.620 134.525 ;
        RECT 76.465 133.395 76.695 134.105 ;
        RECT 76.865 133.215 77.195 133.925 ;
        RECT 77.365 133.395 77.625 134.105 ;
        RECT 77.905 134.145 78.620 134.315 ;
        RECT 78.875 134.290 79.045 135.020 ;
        RECT 79.220 134.925 79.480 135.765 ;
        RECT 80.115 135.040 80.405 135.765 ;
        RECT 80.595 134.955 80.835 135.765 ;
        RECT 81.005 134.955 81.335 135.595 ;
        RECT 81.505 134.955 81.775 135.765 ;
        RECT 81.955 135.015 83.165 135.765 ;
        RECT 83.370 135.025 83.985 135.595 ;
        RECT 84.155 135.255 84.370 135.765 ;
        RECT 84.600 135.255 84.880 135.585 ;
        RECT 85.060 135.255 85.300 135.765 ;
        RECT 80.575 134.525 80.925 134.775 ;
        RECT 77.905 133.385 78.075 134.145 ;
        RECT 78.290 133.215 78.620 133.975 ;
        RECT 78.790 133.385 79.045 134.290 ;
        RECT 79.220 133.215 79.480 134.365 ;
        RECT 80.115 133.215 80.405 134.380 ;
        RECT 81.095 134.355 81.265 134.955 ;
        RECT 81.435 134.525 81.785 134.775 ;
        RECT 81.955 134.475 82.475 135.015 ;
        RECT 80.585 134.185 81.265 134.355 ;
        RECT 80.585 133.400 80.915 134.185 ;
        RECT 81.445 133.215 81.775 134.355 ;
        RECT 82.645 134.305 83.165 134.845 ;
        RECT 81.955 133.215 83.165 134.305 ;
        RECT 83.370 134.005 83.685 135.025 ;
        RECT 83.855 134.355 84.025 134.855 ;
        RECT 84.275 134.525 84.540 135.085 ;
        RECT 84.710 134.355 84.880 135.255 ;
        RECT 85.660 135.115 85.970 135.585 ;
        RECT 86.140 135.285 86.875 135.765 ;
        RECT 87.045 135.195 87.215 135.545 ;
        RECT 87.385 135.365 87.765 135.765 ;
        RECT 85.050 134.525 85.405 135.085 ;
        RECT 85.660 134.945 86.395 135.115 ;
        RECT 87.045 135.025 87.785 135.195 ;
        RECT 87.955 135.090 88.225 135.435 ;
        RECT 86.145 134.855 86.395 134.945 ;
        RECT 87.615 134.855 87.785 135.025 ;
        RECT 85.640 134.525 85.975 134.775 ;
        RECT 86.145 134.525 86.885 134.855 ;
        RECT 87.615 134.525 87.845 134.855 ;
        RECT 83.855 134.185 85.280 134.355 ;
        RECT 83.370 133.385 83.905 134.005 ;
        RECT 84.075 133.215 84.405 134.015 ;
        RECT 84.890 134.010 85.280 134.185 ;
        RECT 85.640 133.215 85.895 134.355 ;
        RECT 86.145 133.965 86.315 134.525 ;
        RECT 87.615 134.355 87.785 134.525 ;
        RECT 88.055 134.355 88.225 135.090 ;
        RECT 88.870 135.195 89.125 135.545 ;
        RECT 89.295 135.365 89.625 135.765 ;
        RECT 89.795 135.195 89.965 135.545 ;
        RECT 90.135 135.365 90.515 135.765 ;
        RECT 88.870 135.025 90.535 135.195 ;
        RECT 90.705 135.090 90.980 135.435 ;
        RECT 90.365 134.855 90.535 135.025 ;
        RECT 88.855 134.525 89.200 134.855 ;
        RECT 89.370 134.525 90.195 134.855 ;
        RECT 90.365 134.525 90.640 134.855 ;
        RECT 86.540 134.185 87.785 134.355 ;
        RECT 86.540 133.935 86.960 134.185 ;
        RECT 86.090 133.435 87.285 133.765 ;
        RECT 87.465 133.215 87.745 134.015 ;
        RECT 87.955 133.385 88.225 134.355 ;
        RECT 88.875 134.065 89.200 134.355 ;
        RECT 89.370 134.235 89.565 134.525 ;
        RECT 90.365 134.355 90.535 134.525 ;
        RECT 90.810 134.355 90.980 135.090 ;
        RECT 91.245 135.085 91.415 135.460 ;
        RECT 91.215 134.915 91.415 135.085 ;
        RECT 91.605 135.235 91.835 135.540 ;
        RECT 92.005 135.405 92.335 135.765 ;
        RECT 92.530 135.235 92.820 135.585 ;
        RECT 91.605 135.065 92.820 135.235 ;
        RECT 91.245 134.895 91.415 134.915 ;
        RECT 92.995 134.995 95.585 135.765 ;
        RECT 91.245 134.725 91.765 134.895 ;
        RECT 89.875 134.185 90.535 134.355 ;
        RECT 89.875 134.065 90.045 134.185 ;
        RECT 88.875 133.895 90.045 134.065 ;
        RECT 88.855 133.435 90.045 133.725 ;
        RECT 90.215 133.215 90.495 134.015 ;
        RECT 90.705 133.385 90.980 134.355 ;
        RECT 91.160 134.195 91.405 134.555 ;
        RECT 91.595 134.345 91.765 134.725 ;
        RECT 91.935 134.525 92.320 134.855 ;
        RECT 92.500 134.745 92.760 134.855 ;
        RECT 92.500 134.575 92.765 134.745 ;
        RECT 92.500 134.525 92.760 134.575 ;
        RECT 91.595 134.065 91.945 134.345 ;
        RECT 91.160 133.215 91.415 134.015 ;
        RECT 91.615 133.385 91.945 134.065 ;
        RECT 92.125 133.475 92.320 134.525 ;
        RECT 92.995 134.475 94.205 134.995 ;
        RECT 96.215 134.965 96.910 135.595 ;
        RECT 97.115 134.965 97.425 135.765 ;
        RECT 97.635 135.255 98.035 135.765 ;
        RECT 98.610 135.150 98.780 135.595 ;
        RECT 98.950 135.365 99.670 135.765 ;
        RECT 99.840 135.195 100.010 135.595 ;
        RECT 100.245 135.320 100.675 135.765 ;
        RECT 92.500 133.215 92.820 134.355 ;
        RECT 94.375 134.305 95.585 134.825 ;
        RECT 96.235 134.525 96.570 134.775 ;
        RECT 96.740 134.365 96.910 134.965 ;
        RECT 97.080 134.525 97.415 134.795 ;
        RECT 92.995 133.215 95.585 134.305 ;
        RECT 96.215 133.215 96.475 134.355 ;
        RECT 96.645 133.385 96.975 134.365 ;
        RECT 97.145 133.215 97.425 134.355 ;
        RECT 97.650 134.195 97.910 135.085 ;
        RECT 98.110 134.495 98.370 135.085 ;
        RECT 98.610 134.980 98.960 135.150 ;
        RECT 98.110 134.195 98.590 134.495 ;
        RECT 97.675 133.845 98.615 134.015 ;
        RECT 97.675 133.385 97.855 133.845 ;
        RECT 98.025 133.215 98.275 133.675 ;
        RECT 98.445 133.595 98.615 133.845 ;
        RECT 98.790 133.955 98.960 134.980 ;
        RECT 99.130 135.025 100.010 135.195 ;
        RECT 100.845 135.040 101.105 135.595 ;
        RECT 99.130 134.305 99.300 135.025 ;
        RECT 99.490 134.475 99.780 134.855 ;
        RECT 99.130 134.135 99.650 134.305 ;
        RECT 99.950 134.235 100.280 134.855 ;
        RECT 100.505 134.525 100.760 134.855 ;
        RECT 98.790 133.785 99.200 133.955 ;
        RECT 99.480 133.945 99.650 134.135 ;
        RECT 100.505 134.045 100.675 134.525 ;
        RECT 100.930 134.325 101.105 135.040 ;
        RECT 98.945 133.650 99.200 133.785 ;
        RECT 99.915 133.875 100.675 134.045 ;
        RECT 99.915 133.650 100.085 133.875 ;
        RECT 98.445 133.425 98.775 133.595 ;
        RECT 98.945 133.480 100.085 133.650 ;
        RECT 98.945 133.385 99.200 133.480 ;
        RECT 100.345 133.215 100.675 133.615 ;
        RECT 100.845 133.385 101.105 134.325 ;
        RECT 101.295 135.265 101.550 135.595 ;
        RECT 101.765 135.285 102.095 135.765 ;
        RECT 102.265 135.345 103.800 135.595 ;
        RECT 101.295 135.185 101.480 135.265 ;
        RECT 101.295 134.065 101.465 135.185 ;
        RECT 102.265 135.115 102.435 135.345 ;
        RECT 101.635 134.945 102.435 135.115 ;
        RECT 101.635 134.395 101.805 134.945 ;
        RECT 102.615 134.775 102.900 135.175 ;
        RECT 102.035 134.575 102.400 134.775 ;
        RECT 102.570 134.575 102.900 134.775 ;
        RECT 103.170 134.775 103.450 135.175 ;
        RECT 103.630 135.115 103.800 135.345 ;
        RECT 104.025 135.285 104.355 135.765 ;
        RECT 104.525 135.115 104.695 135.595 ;
        RECT 103.630 134.945 104.695 135.115 ;
        RECT 105.875 135.040 106.165 135.765 ;
        RECT 106.335 134.995 108.005 135.765 ;
        RECT 108.190 135.375 109.360 135.595 ;
        RECT 109.550 135.375 111.640 135.595 ;
        RECT 103.170 134.575 103.645 134.775 ;
        RECT 103.815 134.575 104.260 134.775 ;
        RECT 104.430 134.565 104.780 134.775 ;
        RECT 106.335 134.475 107.085 134.995 ;
        RECT 108.190 134.955 108.440 135.375 ;
        RECT 109.110 135.205 109.360 135.375 ;
        RECT 108.610 134.985 108.940 135.205 ;
        RECT 101.635 134.225 104.695 134.395 ;
        RECT 101.295 134.055 101.505 134.065 ;
        RECT 101.295 133.385 101.550 134.055 ;
        RECT 101.720 133.215 102.050 133.975 ;
        RECT 102.220 133.815 103.855 134.055 ;
        RECT 102.220 133.385 102.470 133.815 ;
        RECT 103.625 133.725 103.855 133.815 ;
        RECT 102.640 133.215 102.995 133.635 ;
        RECT 103.185 133.555 103.515 133.595 ;
        RECT 104.025 133.555 104.355 134.055 ;
        RECT 103.185 133.385 104.355 133.555 ;
        RECT 104.525 133.385 104.695 134.225 ;
        RECT 105.875 133.215 106.165 134.380 ;
        RECT 107.255 134.305 108.005 134.825 ;
        RECT 108.175 134.575 108.525 134.775 ;
        RECT 108.695 134.405 108.940 134.985 ;
        RECT 109.110 134.945 111.140 135.205 ;
        RECT 111.310 135.115 111.640 135.375 ;
        RECT 111.810 135.295 111.980 135.765 ;
        RECT 112.150 135.125 112.480 135.595 ;
        RECT 112.650 135.295 112.820 135.765 ;
        RECT 112.990 135.125 113.320 135.595 ;
        RECT 112.150 135.115 113.320 135.125 ;
        RECT 111.310 134.945 113.320 135.115 ;
        RECT 114.820 134.985 115.320 135.595 ;
        RECT 106.335 133.215 108.005 134.305 ;
        RECT 108.230 133.215 108.480 134.395 ;
        RECT 108.650 134.065 108.940 134.405 ;
        RECT 109.110 134.405 110.125 134.775 ;
        RECT 110.295 134.575 110.850 134.775 ;
        RECT 111.020 134.405 111.350 134.775 ;
        RECT 109.110 134.235 111.350 134.405 ;
        RECT 111.520 134.405 111.850 134.775 ;
        RECT 112.070 134.575 112.565 134.775 ;
        RECT 112.735 134.575 113.525 134.775 ;
        RECT 112.735 134.405 112.905 134.575 ;
        RECT 114.615 134.525 114.965 134.775 ;
        RECT 111.520 134.235 112.905 134.405 ;
        RECT 108.650 133.895 112.440 134.065 ;
        RECT 108.650 133.385 108.900 133.895 ;
        RECT 110.430 133.725 110.680 133.895 ;
        RECT 112.190 133.725 112.440 133.895 ;
        RECT 109.070 133.215 109.840 133.725 ;
        RECT 110.010 133.555 110.260 133.725 ;
        RECT 110.850 133.555 111.100 133.725 ;
        RECT 110.010 133.385 111.100 133.555 ;
        RECT 111.270 133.215 111.600 133.725 ;
        RECT 111.770 133.555 112.020 133.725 ;
        RECT 112.610 133.555 112.860 134.065 ;
        RECT 111.770 133.385 112.860 133.555 ;
        RECT 113.075 133.215 113.280 134.395 ;
        RECT 115.150 134.355 115.320 134.985 ;
        RECT 115.950 135.115 116.280 135.595 ;
        RECT 116.450 135.305 116.675 135.765 ;
        RECT 116.845 135.115 117.175 135.595 ;
        RECT 115.950 134.945 117.175 135.115 ;
        RECT 117.365 134.965 117.615 135.765 ;
        RECT 117.785 134.965 118.125 135.595 ;
        RECT 118.295 135.155 118.635 135.570 ;
        RECT 118.805 135.325 118.975 135.765 ;
        RECT 119.145 135.375 120.395 135.555 ;
        RECT 119.145 135.155 119.475 135.375 ;
        RECT 120.665 135.305 120.835 135.765 ;
        RECT 118.295 134.985 119.475 135.155 ;
        RECT 119.645 135.135 120.010 135.205 ;
        RECT 115.490 134.575 115.820 134.775 ;
        RECT 115.990 134.575 116.320 134.775 ;
        RECT 116.490 134.575 116.910 134.775 ;
        RECT 117.085 134.605 117.780 134.775 ;
        RECT 117.085 134.355 117.255 134.605 ;
        RECT 117.950 134.405 118.125 134.965 ;
        RECT 119.645 134.955 120.895 135.135 ;
        RECT 118.295 134.575 118.760 134.775 ;
        RECT 118.935 134.525 119.265 134.775 ;
        RECT 119.435 134.745 119.900 134.775 ;
        RECT 119.435 134.575 119.905 134.745 ;
        RECT 119.435 134.525 119.900 134.575 ;
        RECT 120.095 134.525 120.450 134.775 ;
        RECT 118.935 134.405 119.115 134.525 ;
        RECT 117.895 134.355 118.125 134.405 ;
        RECT 114.820 134.185 117.255 134.355 ;
        RECT 114.820 133.385 115.150 134.185 ;
        RECT 115.320 133.215 115.650 134.015 ;
        RECT 115.950 133.385 116.280 134.185 ;
        RECT 116.925 133.215 117.175 134.015 ;
        RECT 117.445 133.215 117.615 134.355 ;
        RECT 117.785 133.385 118.125 134.355 ;
        RECT 118.295 133.215 118.615 134.395 ;
        RECT 118.785 134.235 119.115 134.405 ;
        RECT 120.620 134.355 120.895 134.955 ;
        RECT 118.785 133.445 118.985 134.235 ;
        RECT 119.285 134.145 120.895 134.355 ;
        RECT 119.285 134.045 119.695 134.145 ;
        RECT 119.310 133.385 119.695 134.045 ;
        RECT 120.090 133.215 120.875 133.975 ;
        RECT 121.065 133.385 121.345 135.485 ;
        RECT 121.515 135.015 122.725 135.765 ;
        RECT 122.895 135.025 123.215 135.505 ;
        RECT 123.385 135.195 123.615 135.595 ;
        RECT 123.785 135.375 124.135 135.765 ;
        RECT 123.385 135.115 123.895 135.195 ;
        RECT 124.305 135.115 124.635 135.595 ;
        RECT 123.385 135.025 124.635 135.115 ;
        RECT 121.515 134.475 122.035 135.015 ;
        RECT 122.205 134.305 122.725 134.845 ;
        RECT 121.515 133.215 122.725 134.305 ;
        RECT 122.895 134.095 123.065 135.025 ;
        RECT 123.725 134.945 124.635 135.025 ;
        RECT 124.805 134.945 124.975 135.765 ;
        RECT 125.480 135.025 125.945 135.570 ;
        RECT 123.235 134.435 123.405 134.855 ;
        RECT 123.635 134.605 124.235 134.775 ;
        RECT 123.235 134.265 123.895 134.435 ;
        RECT 122.895 133.895 123.555 134.095 ;
        RECT 123.725 134.065 123.895 134.265 ;
        RECT 124.065 134.405 124.235 134.605 ;
        RECT 124.405 134.575 125.100 134.775 ;
        RECT 125.360 134.405 125.605 134.855 ;
        RECT 124.065 134.235 125.605 134.405 ;
        RECT 125.775 134.065 125.945 135.025 ;
        RECT 123.725 133.895 125.945 134.065 ;
        RECT 127.040 134.165 127.375 135.585 ;
        RECT 127.555 135.395 128.300 135.765 ;
        RECT 128.865 135.225 129.120 135.585 ;
        RECT 129.300 135.395 129.630 135.765 ;
        RECT 129.810 135.225 130.035 135.585 ;
        RECT 127.550 135.035 130.035 135.225 ;
        RECT 127.550 134.345 127.775 135.035 ;
        RECT 130.255 135.015 131.465 135.765 ;
        RECT 131.635 135.040 131.925 135.765 ;
        RECT 132.095 135.385 132.985 135.555 ;
        RECT 127.975 134.525 128.255 134.855 ;
        RECT 128.435 134.525 129.010 134.855 ;
        RECT 129.190 134.525 129.625 134.855 ;
        RECT 129.805 134.525 130.075 134.855 ;
        RECT 130.255 134.475 130.775 135.015 ;
        RECT 127.550 134.165 130.045 134.345 ;
        RECT 130.945 134.305 131.465 134.845 ;
        RECT 132.095 134.830 132.645 135.215 ;
        RECT 132.815 134.660 132.985 135.385 ;
        RECT 132.095 134.590 132.985 134.660 ;
        RECT 133.155 135.085 133.375 135.545 ;
        RECT 133.545 135.225 133.795 135.765 ;
        RECT 133.965 135.115 134.225 135.595 ;
        RECT 133.155 135.060 133.405 135.085 ;
        RECT 133.155 134.635 133.485 135.060 ;
        RECT 132.095 134.565 132.990 134.590 ;
        RECT 132.095 134.550 133.000 134.565 ;
        RECT 132.095 134.535 133.005 134.550 ;
        RECT 132.095 134.530 133.015 134.535 ;
        RECT 132.095 134.520 133.020 134.530 ;
        RECT 132.095 134.510 133.025 134.520 ;
        RECT 132.095 134.505 133.035 134.510 ;
        RECT 132.095 134.495 133.045 134.505 ;
        RECT 132.095 134.490 133.055 134.495 ;
        RECT 123.385 133.725 123.555 133.895 ;
        RECT 122.915 133.215 123.215 133.725 ;
        RECT 123.385 133.555 123.765 133.725 ;
        RECT 124.345 133.215 124.975 133.725 ;
        RECT 125.145 133.385 125.475 133.895 ;
        RECT 125.645 133.215 125.945 133.725 ;
        RECT 127.040 133.395 127.305 134.165 ;
        RECT 127.475 133.215 127.805 133.935 ;
        RECT 127.995 133.755 129.185 133.985 ;
        RECT 127.995 133.395 128.255 133.755 ;
        RECT 128.425 133.215 128.755 133.585 ;
        RECT 128.925 133.395 129.185 133.755 ;
        RECT 129.755 133.395 130.045 134.165 ;
        RECT 130.255 133.215 131.465 134.305 ;
        RECT 131.635 133.215 131.925 134.380 ;
        RECT 132.095 134.040 132.355 134.490 ;
        RECT 132.720 134.485 133.055 134.490 ;
        RECT 132.720 134.480 133.070 134.485 ;
        RECT 132.720 134.470 133.085 134.480 ;
        RECT 132.720 134.465 133.110 134.470 ;
        RECT 133.655 134.465 133.885 134.860 ;
        RECT 132.720 134.460 133.885 134.465 ;
        RECT 132.750 134.425 133.885 134.460 ;
        RECT 132.785 134.400 133.885 134.425 ;
        RECT 132.815 134.370 133.885 134.400 ;
        RECT 132.835 134.340 133.885 134.370 ;
        RECT 132.855 134.310 133.885 134.340 ;
        RECT 132.925 134.300 133.885 134.310 ;
        RECT 132.950 134.290 133.885 134.300 ;
        RECT 132.970 134.275 133.885 134.290 ;
        RECT 132.990 134.260 133.885 134.275 ;
        RECT 132.995 134.250 133.780 134.260 ;
        RECT 133.010 134.215 133.780 134.250 ;
        RECT 132.525 133.895 132.855 134.140 ;
        RECT 133.025 133.965 133.780 134.215 ;
        RECT 134.055 134.085 134.225 135.115 ;
        RECT 132.525 133.870 132.710 133.895 ;
        RECT 132.095 133.770 132.710 133.870 ;
        RECT 132.095 133.215 132.700 133.770 ;
        RECT 132.875 133.385 133.355 133.725 ;
        RECT 133.525 133.215 133.780 133.760 ;
        RECT 133.950 133.385 134.225 134.085 ;
        RECT 134.395 135.025 134.860 135.570 ;
        RECT 134.395 134.065 134.565 135.025 ;
        RECT 135.365 134.945 135.535 135.765 ;
        RECT 135.705 135.115 136.035 135.595 ;
        RECT 136.205 135.375 136.555 135.765 ;
        RECT 136.725 135.195 136.955 135.595 ;
        RECT 136.445 135.115 136.955 135.195 ;
        RECT 135.705 135.025 136.955 135.115 ;
        RECT 137.125 135.025 137.445 135.505 ;
        RECT 137.780 135.255 138.020 135.765 ;
        RECT 138.200 135.255 138.480 135.585 ;
        RECT 138.710 135.255 138.925 135.765 ;
        RECT 135.705 134.945 136.615 135.025 ;
        RECT 134.735 134.405 134.980 134.855 ;
        RECT 135.240 134.575 135.935 134.775 ;
        RECT 136.105 134.605 136.705 134.775 ;
        RECT 136.105 134.405 136.275 134.605 ;
        RECT 136.935 134.435 137.105 134.855 ;
        RECT 134.735 134.235 136.275 134.405 ;
        RECT 136.445 134.265 137.105 134.435 ;
        RECT 136.445 134.065 136.615 134.265 ;
        RECT 137.275 134.095 137.445 135.025 ;
        RECT 137.675 134.525 138.030 135.085 ;
        RECT 138.200 134.355 138.370 135.255 ;
        RECT 138.540 134.525 138.805 135.085 ;
        RECT 139.095 135.025 139.710 135.595 ;
        RECT 139.915 135.220 145.260 135.765 ;
        RECT 145.435 135.220 150.780 135.765 ;
        RECT 150.955 135.220 156.300 135.765 ;
        RECT 139.055 134.355 139.225 134.855 ;
        RECT 134.395 133.895 136.615 134.065 ;
        RECT 136.785 133.895 137.445 134.095 ;
        RECT 137.800 134.185 139.225 134.355 ;
        RECT 137.800 134.010 138.190 134.185 ;
        RECT 134.395 133.215 134.695 133.725 ;
        RECT 134.865 133.385 135.195 133.895 ;
        RECT 136.785 133.725 136.955 133.895 ;
        RECT 135.365 133.215 135.995 133.725 ;
        RECT 136.575 133.555 136.955 133.725 ;
        RECT 137.125 133.215 137.425 133.725 ;
        RECT 138.675 133.215 139.005 134.015 ;
        RECT 139.395 134.005 139.710 135.025 ;
        RECT 141.500 134.390 141.840 135.220 ;
        RECT 139.175 133.385 139.710 134.005 ;
        RECT 143.320 133.650 143.670 134.900 ;
        RECT 147.020 134.390 147.360 135.220 ;
        RECT 148.840 133.650 149.190 134.900 ;
        RECT 152.540 134.390 152.880 135.220 ;
        RECT 156.935 135.015 158.145 135.765 ;
        RECT 154.360 133.650 154.710 134.900 ;
        RECT 156.935 134.305 157.455 134.845 ;
        RECT 157.625 134.475 158.145 135.015 ;
        RECT 139.915 133.215 145.260 133.650 ;
        RECT 145.435 133.215 150.780 133.650 ;
        RECT 150.955 133.215 156.300 133.650 ;
        RECT 156.935 133.215 158.145 134.305 ;
        RECT 2.750 133.045 158.230 133.215 ;
        RECT 2.835 131.955 4.045 133.045 ;
        RECT 2.835 131.245 3.355 131.785 ;
        RECT 3.525 131.415 4.045 131.955 ;
        RECT 4.305 132.115 4.475 132.875 ;
        RECT 4.655 132.285 4.985 133.045 ;
        RECT 4.305 131.945 4.970 132.115 ;
        RECT 5.155 131.970 5.425 132.875 ;
        RECT 5.600 132.375 5.855 132.875 ;
        RECT 6.025 132.545 6.355 133.045 ;
        RECT 5.600 132.205 6.350 132.375 ;
        RECT 4.800 131.800 4.970 131.945 ;
        RECT 4.235 131.395 4.565 131.765 ;
        RECT 4.800 131.470 5.085 131.800 ;
        RECT 2.835 130.495 4.045 131.245 ;
        RECT 4.800 131.215 4.970 131.470 ;
        RECT 4.305 131.045 4.970 131.215 ;
        RECT 5.255 131.170 5.425 131.970 ;
        RECT 5.600 131.385 5.950 132.035 ;
        RECT 6.120 131.215 6.350 132.205 ;
        RECT 4.305 130.665 4.475 131.045 ;
        RECT 4.655 130.495 4.985 130.875 ;
        RECT 5.165 130.665 5.425 131.170 ;
        RECT 5.600 131.045 6.350 131.215 ;
        RECT 5.600 130.755 5.855 131.045 ;
        RECT 6.025 130.495 6.355 130.875 ;
        RECT 6.525 130.755 6.695 132.875 ;
        RECT 6.865 132.075 7.190 132.860 ;
        RECT 7.360 132.585 7.610 133.045 ;
        RECT 7.780 132.545 8.030 132.875 ;
        RECT 8.245 132.545 8.925 132.875 ;
        RECT 7.780 132.415 7.950 132.545 ;
        RECT 7.555 132.245 7.950 132.415 ;
        RECT 6.925 131.025 7.385 132.075 ;
        RECT 7.555 130.885 7.725 132.245 ;
        RECT 8.120 131.985 8.585 132.375 ;
        RECT 7.895 131.175 8.245 131.795 ;
        RECT 8.415 131.395 8.585 131.985 ;
        RECT 8.755 131.765 8.925 132.545 ;
        RECT 9.095 132.445 9.265 132.785 ;
        RECT 9.500 132.615 9.830 133.045 ;
        RECT 10.000 132.445 10.170 132.785 ;
        RECT 10.465 132.585 10.835 133.045 ;
        RECT 9.095 132.275 10.170 132.445 ;
        RECT 11.005 132.415 11.175 132.875 ;
        RECT 11.410 132.535 12.280 132.875 ;
        RECT 12.450 132.585 12.700 133.045 ;
        RECT 10.615 132.245 11.175 132.415 ;
        RECT 10.615 132.105 10.785 132.245 ;
        RECT 9.285 131.935 10.785 132.105 ;
        RECT 11.480 132.075 11.940 132.365 ;
        RECT 8.755 131.595 10.445 131.765 ;
        RECT 8.415 131.175 8.770 131.395 ;
        RECT 8.940 130.885 9.110 131.595 ;
        RECT 9.315 131.175 10.105 131.425 ;
        RECT 10.275 131.415 10.445 131.595 ;
        RECT 10.615 131.245 10.785 131.935 ;
        RECT 7.055 130.495 7.385 130.855 ;
        RECT 7.555 130.715 8.050 130.885 ;
        RECT 8.255 130.715 9.110 130.885 ;
        RECT 9.985 130.495 10.315 130.955 ;
        RECT 10.525 130.855 10.785 131.245 ;
        RECT 10.975 132.065 11.940 132.075 ;
        RECT 12.110 132.155 12.280 132.535 ;
        RECT 12.870 132.495 13.040 132.785 ;
        RECT 13.220 132.665 13.550 133.045 ;
        RECT 12.870 132.325 13.670 132.495 ;
        RECT 10.975 131.905 11.650 132.065 ;
        RECT 12.110 131.985 13.330 132.155 ;
        RECT 10.975 131.115 11.185 131.905 ;
        RECT 12.110 131.895 12.280 131.985 ;
        RECT 11.355 131.115 11.705 131.735 ;
        RECT 11.875 131.725 12.280 131.895 ;
        RECT 11.875 130.945 12.045 131.725 ;
        RECT 12.215 131.275 12.435 131.555 ;
        RECT 12.615 131.445 13.155 131.815 ;
        RECT 13.500 131.735 13.670 132.325 ;
        RECT 13.890 131.905 14.195 133.045 ;
        RECT 14.365 131.855 14.620 132.735 ;
        RECT 15.715 131.880 16.005 133.045 ;
        RECT 16.180 131.905 16.515 132.875 ;
        RECT 16.685 131.905 16.855 133.045 ;
        RECT 17.025 132.705 19.055 132.875 ;
        RECT 13.500 131.705 14.240 131.735 ;
        RECT 12.215 131.105 12.745 131.275 ;
        RECT 10.525 130.685 10.875 130.855 ;
        RECT 11.095 130.665 12.045 130.945 ;
        RECT 12.215 130.495 12.405 130.935 ;
        RECT 12.575 130.875 12.745 131.105 ;
        RECT 12.915 131.045 13.155 131.445 ;
        RECT 13.325 131.405 14.240 131.705 ;
        RECT 13.325 131.230 13.650 131.405 ;
        RECT 13.325 130.875 13.645 131.230 ;
        RECT 14.410 131.205 14.620 131.855 ;
        RECT 16.180 131.235 16.350 131.905 ;
        RECT 17.025 131.735 17.195 132.705 ;
        RECT 16.520 131.405 16.775 131.735 ;
        RECT 17.000 131.405 17.195 131.735 ;
        RECT 17.365 132.365 18.490 132.535 ;
        RECT 16.605 131.235 16.775 131.405 ;
        RECT 17.365 131.235 17.535 132.365 ;
        RECT 12.575 130.705 13.645 130.875 ;
        RECT 13.890 130.495 14.195 130.955 ;
        RECT 14.365 130.675 14.620 131.205 ;
        RECT 15.715 130.495 16.005 131.220 ;
        RECT 16.180 130.665 16.435 131.235 ;
        RECT 16.605 131.065 17.535 131.235 ;
        RECT 17.705 132.025 18.715 132.195 ;
        RECT 17.705 131.225 17.875 132.025 ;
        RECT 17.360 131.030 17.535 131.065 ;
        RECT 16.605 130.495 16.935 130.895 ;
        RECT 17.360 130.665 17.890 131.030 ;
        RECT 18.080 131.005 18.355 131.825 ;
        RECT 18.075 130.835 18.355 131.005 ;
        RECT 18.080 130.665 18.355 130.835 ;
        RECT 18.525 130.665 18.715 132.025 ;
        RECT 18.885 132.040 19.055 132.705 ;
        RECT 19.225 132.285 19.395 133.045 ;
        RECT 19.630 132.285 20.145 132.695 ;
        RECT 18.885 131.850 19.635 132.040 ;
        RECT 19.805 131.475 20.145 132.285 ;
        RECT 18.915 131.305 20.145 131.475 ;
        RECT 21.235 131.970 21.505 132.875 ;
        RECT 21.675 132.285 22.005 133.045 ;
        RECT 22.185 132.115 22.355 132.875 ;
        RECT 22.620 132.375 22.875 132.875 ;
        RECT 23.045 132.545 23.375 133.045 ;
        RECT 22.620 132.205 23.370 132.375 ;
        RECT 18.895 130.495 19.405 131.030 ;
        RECT 19.625 130.700 19.870 131.305 ;
        RECT 21.235 131.170 21.405 131.970 ;
        RECT 21.690 131.945 22.355 132.115 ;
        RECT 21.690 131.800 21.860 131.945 ;
        RECT 21.575 131.470 21.860 131.800 ;
        RECT 21.690 131.215 21.860 131.470 ;
        RECT 22.095 131.395 22.425 131.765 ;
        RECT 22.620 131.385 22.970 132.035 ;
        RECT 23.140 131.215 23.370 132.205 ;
        RECT 21.235 130.665 21.495 131.170 ;
        RECT 21.690 131.045 22.355 131.215 ;
        RECT 21.675 130.495 22.005 130.875 ;
        RECT 22.185 130.665 22.355 131.045 ;
        RECT 22.620 131.045 23.370 131.215 ;
        RECT 22.620 130.755 22.875 131.045 ;
        RECT 23.045 130.495 23.375 130.875 ;
        RECT 23.545 130.755 23.715 132.875 ;
        RECT 23.885 132.075 24.210 132.860 ;
        RECT 24.380 132.585 24.630 133.045 ;
        RECT 24.800 132.545 25.050 132.875 ;
        RECT 25.265 132.545 25.945 132.875 ;
        RECT 24.800 132.415 24.970 132.545 ;
        RECT 24.575 132.245 24.970 132.415 ;
        RECT 23.945 131.025 24.405 132.075 ;
        RECT 24.575 130.885 24.745 132.245 ;
        RECT 25.140 131.985 25.605 132.375 ;
        RECT 24.915 131.175 25.265 131.795 ;
        RECT 25.435 131.395 25.605 131.985 ;
        RECT 25.775 131.765 25.945 132.545 ;
        RECT 26.115 132.445 26.285 132.785 ;
        RECT 26.520 132.615 26.850 133.045 ;
        RECT 27.020 132.445 27.190 132.785 ;
        RECT 27.485 132.585 27.855 133.045 ;
        RECT 26.115 132.275 27.190 132.445 ;
        RECT 28.025 132.415 28.195 132.875 ;
        RECT 28.430 132.535 29.300 132.875 ;
        RECT 29.470 132.585 29.720 133.045 ;
        RECT 27.635 132.245 28.195 132.415 ;
        RECT 27.635 132.105 27.805 132.245 ;
        RECT 26.305 131.935 27.805 132.105 ;
        RECT 28.500 132.075 28.960 132.365 ;
        RECT 25.775 131.595 27.465 131.765 ;
        RECT 25.435 131.175 25.790 131.395 ;
        RECT 25.960 130.885 26.130 131.595 ;
        RECT 26.335 131.175 27.125 131.425 ;
        RECT 27.295 131.415 27.465 131.595 ;
        RECT 27.635 131.245 27.805 131.935 ;
        RECT 24.075 130.495 24.405 130.855 ;
        RECT 24.575 130.715 25.070 130.885 ;
        RECT 25.275 130.715 26.130 130.885 ;
        RECT 27.005 130.495 27.335 130.955 ;
        RECT 27.545 130.855 27.805 131.245 ;
        RECT 27.995 132.065 28.960 132.075 ;
        RECT 29.130 132.155 29.300 132.535 ;
        RECT 29.890 132.495 30.060 132.785 ;
        RECT 30.240 132.665 30.570 133.045 ;
        RECT 29.890 132.325 30.690 132.495 ;
        RECT 27.995 131.905 28.670 132.065 ;
        RECT 29.130 131.985 30.350 132.155 ;
        RECT 27.995 131.115 28.205 131.905 ;
        RECT 29.130 131.895 29.300 131.985 ;
        RECT 28.375 131.115 28.725 131.735 ;
        RECT 28.895 131.725 29.300 131.895 ;
        RECT 28.895 130.945 29.065 131.725 ;
        RECT 29.235 131.275 29.455 131.555 ;
        RECT 29.635 131.445 30.175 131.815 ;
        RECT 30.520 131.735 30.690 132.325 ;
        RECT 30.910 131.905 31.215 133.045 ;
        RECT 31.385 131.855 31.640 132.735 ;
        RECT 31.930 132.415 32.215 132.875 ;
        RECT 32.385 132.585 32.655 133.045 ;
        RECT 31.930 132.195 32.885 132.415 ;
        RECT 30.520 131.705 31.260 131.735 ;
        RECT 29.235 131.105 29.765 131.275 ;
        RECT 27.545 130.685 27.895 130.855 ;
        RECT 28.115 130.665 29.065 130.945 ;
        RECT 29.235 130.495 29.425 130.935 ;
        RECT 29.595 130.875 29.765 131.105 ;
        RECT 29.935 131.045 30.175 131.445 ;
        RECT 30.345 131.405 31.260 131.705 ;
        RECT 30.345 131.230 30.670 131.405 ;
        RECT 30.345 130.875 30.665 131.230 ;
        RECT 31.430 131.205 31.640 131.855 ;
        RECT 31.815 131.465 32.505 132.025 ;
        RECT 32.675 131.295 32.885 132.195 ;
        RECT 29.595 130.705 30.665 130.875 ;
        RECT 30.910 130.495 31.215 130.955 ;
        RECT 31.385 130.675 31.640 131.205 ;
        RECT 31.930 131.125 32.885 131.295 ;
        RECT 33.055 132.025 33.455 132.875 ;
        RECT 33.645 132.415 33.925 132.875 ;
        RECT 34.445 132.585 34.770 133.045 ;
        RECT 33.645 132.195 34.770 132.415 ;
        RECT 33.055 131.465 34.150 132.025 ;
        RECT 34.320 131.735 34.770 132.195 ;
        RECT 34.940 131.905 35.325 132.875 ;
        RECT 31.930 130.665 32.215 131.125 ;
        RECT 32.385 130.495 32.655 130.955 ;
        RECT 33.055 130.665 33.455 131.465 ;
        RECT 34.320 131.405 34.875 131.735 ;
        RECT 34.320 131.295 34.770 131.405 ;
        RECT 33.645 131.125 34.770 131.295 ;
        RECT 35.045 131.235 35.325 131.905 ;
        RECT 33.645 130.665 33.925 131.125 ;
        RECT 34.445 130.495 34.770 130.955 ;
        RECT 34.940 130.665 35.325 131.235 ;
        RECT 35.500 131.905 35.835 132.875 ;
        RECT 36.005 131.905 36.175 133.045 ;
        RECT 36.345 132.705 38.375 132.875 ;
        RECT 35.500 131.235 35.670 131.905 ;
        RECT 36.345 131.735 36.515 132.705 ;
        RECT 35.840 131.405 36.095 131.735 ;
        RECT 36.320 131.405 36.515 131.735 ;
        RECT 36.685 132.365 37.810 132.535 ;
        RECT 35.925 131.235 36.095 131.405 ;
        RECT 36.685 131.235 36.855 132.365 ;
        RECT 35.500 130.665 35.755 131.235 ;
        RECT 35.925 131.065 36.855 131.235 ;
        RECT 37.025 132.025 38.035 132.195 ;
        RECT 37.025 131.225 37.195 132.025 ;
        RECT 37.400 131.685 37.675 131.825 ;
        RECT 37.395 131.515 37.675 131.685 ;
        RECT 36.680 131.030 36.855 131.065 ;
        RECT 35.925 130.495 36.255 130.895 ;
        RECT 36.680 130.665 37.210 131.030 ;
        RECT 37.400 130.665 37.675 131.515 ;
        RECT 37.845 130.665 38.035 132.025 ;
        RECT 38.205 132.040 38.375 132.705 ;
        RECT 38.545 132.285 38.715 133.045 ;
        RECT 38.950 132.285 39.465 132.695 ;
        RECT 38.205 131.850 38.955 132.040 ;
        RECT 39.125 131.475 39.465 132.285 ;
        RECT 40.185 132.115 40.355 132.875 ;
        RECT 40.535 132.285 40.865 133.045 ;
        RECT 40.185 131.945 40.850 132.115 ;
        RECT 41.035 131.970 41.305 132.875 ;
        RECT 40.680 131.800 40.850 131.945 ;
        RECT 38.235 131.305 39.465 131.475 ;
        RECT 40.115 131.395 40.445 131.765 ;
        RECT 40.680 131.470 40.965 131.800 ;
        RECT 38.215 130.495 38.725 131.030 ;
        RECT 38.945 130.700 39.190 131.305 ;
        RECT 40.680 131.215 40.850 131.470 ;
        RECT 40.185 131.045 40.850 131.215 ;
        RECT 41.135 131.170 41.305 131.970 ;
        RECT 41.475 131.880 41.765 133.045 ;
        RECT 42.025 132.115 42.195 132.875 ;
        RECT 42.375 132.285 42.705 133.045 ;
        RECT 42.025 131.945 42.690 132.115 ;
        RECT 42.875 131.970 43.145 132.875 ;
        RECT 42.520 131.800 42.690 131.945 ;
        RECT 41.955 131.395 42.285 131.765 ;
        RECT 42.520 131.470 42.805 131.800 ;
        RECT 40.185 130.665 40.355 131.045 ;
        RECT 40.535 130.495 40.865 130.875 ;
        RECT 41.045 130.665 41.305 131.170 ;
        RECT 41.475 130.495 41.765 131.220 ;
        RECT 42.520 131.215 42.690 131.470 ;
        RECT 42.025 131.045 42.690 131.215 ;
        RECT 42.975 131.170 43.145 131.970 ;
        RECT 43.315 132.285 43.830 132.695 ;
        RECT 44.065 132.285 44.235 133.045 ;
        RECT 44.405 132.705 46.435 132.875 ;
        RECT 43.315 131.475 43.655 132.285 ;
        RECT 44.405 132.040 44.575 132.705 ;
        RECT 44.970 132.365 46.095 132.535 ;
        RECT 43.825 131.850 44.575 132.040 ;
        RECT 44.745 132.025 45.755 132.195 ;
        RECT 43.315 131.305 44.545 131.475 ;
        RECT 42.025 130.665 42.195 131.045 ;
        RECT 42.375 130.495 42.705 130.875 ;
        RECT 42.885 130.665 43.145 131.170 ;
        RECT 43.590 130.700 43.835 131.305 ;
        RECT 44.055 130.495 44.565 131.030 ;
        RECT 44.745 130.665 44.935 132.025 ;
        RECT 45.105 131.345 45.380 131.825 ;
        RECT 45.105 131.175 45.385 131.345 ;
        RECT 45.585 131.225 45.755 132.025 ;
        RECT 45.925 131.235 46.095 132.365 ;
        RECT 46.265 131.735 46.435 132.705 ;
        RECT 46.605 131.905 46.775 133.045 ;
        RECT 46.945 131.905 47.280 132.875 ;
        RECT 47.455 132.035 47.715 133.045 ;
        RECT 47.885 132.205 48.160 132.875 ;
        RECT 46.265 131.405 46.460 131.735 ;
        RECT 46.685 131.405 46.940 131.735 ;
        RECT 46.685 131.235 46.855 131.405 ;
        RECT 47.110 131.235 47.280 131.905 ;
        RECT 47.885 131.855 48.055 132.205 ;
        RECT 48.360 132.200 48.575 133.045 ;
        RECT 48.760 132.535 49.235 132.875 ;
        RECT 49.415 132.540 50.045 133.045 ;
        RECT 49.415 132.365 49.605 132.540 ;
        RECT 48.800 132.005 49.050 132.300 ;
        RECT 49.275 132.175 49.605 132.365 ;
        RECT 49.775 132.005 50.030 132.370 ;
        RECT 47.455 131.335 48.070 131.855 ;
        RECT 48.240 131.835 50.030 132.005 ;
        RECT 50.220 131.905 50.555 132.875 ;
        RECT 50.725 131.905 50.895 133.045 ;
        RECT 51.065 132.705 53.095 132.875 ;
        RECT 48.240 131.405 48.470 131.835 ;
        RECT 45.105 130.665 45.380 131.175 ;
        RECT 45.925 131.065 46.855 131.235 ;
        RECT 45.925 131.030 46.100 131.065 ;
        RECT 45.570 130.665 46.100 131.030 ;
        RECT 46.525 130.495 46.855 130.895 ;
        RECT 47.025 130.665 47.280 131.235 ;
        RECT 47.455 130.495 47.730 131.155 ;
        RECT 47.900 131.125 48.070 131.335 ;
        RECT 48.655 131.160 49.065 131.655 ;
        RECT 47.900 130.665 48.150 131.125 ;
        RECT 48.325 130.495 48.655 130.990 ;
        RECT 48.835 130.715 49.065 131.160 ;
        RECT 49.235 130.980 49.490 131.835 ;
        RECT 49.660 131.175 50.045 131.655 ;
        RECT 50.220 131.235 50.390 131.905 ;
        RECT 51.065 131.735 51.235 132.705 ;
        RECT 50.560 131.405 50.815 131.735 ;
        RECT 51.040 131.405 51.235 131.735 ;
        RECT 51.405 132.365 52.530 132.535 ;
        RECT 50.645 131.235 50.815 131.405 ;
        RECT 51.405 131.235 51.575 132.365 ;
        RECT 49.235 130.715 50.025 130.980 ;
        RECT 50.220 130.665 50.475 131.235 ;
        RECT 50.645 131.065 51.575 131.235 ;
        RECT 51.745 132.025 52.755 132.195 ;
        RECT 51.745 131.225 51.915 132.025 ;
        RECT 51.400 131.030 51.575 131.065 ;
        RECT 50.645 130.495 50.975 130.895 ;
        RECT 51.400 130.665 51.930 131.030 ;
        RECT 52.120 131.005 52.395 131.825 ;
        RECT 52.115 130.835 52.395 131.005 ;
        RECT 52.120 130.665 52.395 130.835 ;
        RECT 52.565 130.665 52.755 132.025 ;
        RECT 52.925 132.040 53.095 132.705 ;
        RECT 53.265 132.285 53.435 133.045 ;
        RECT 53.670 132.285 54.185 132.695 ;
        RECT 52.925 131.850 53.675 132.040 ;
        RECT 53.845 131.475 54.185 132.285 ;
        RECT 52.955 131.305 54.185 131.475 ;
        RECT 54.360 131.905 54.695 132.875 ;
        RECT 54.865 131.905 55.035 133.045 ;
        RECT 55.205 132.705 57.235 132.875 ;
        RECT 52.935 130.495 53.445 131.030 ;
        RECT 53.665 130.700 53.910 131.305 ;
        RECT 54.360 131.235 54.530 131.905 ;
        RECT 55.205 131.735 55.375 132.705 ;
        RECT 54.700 131.405 54.955 131.735 ;
        RECT 55.180 131.405 55.375 131.735 ;
        RECT 55.545 132.365 56.670 132.535 ;
        RECT 54.785 131.235 54.955 131.405 ;
        RECT 55.545 131.235 55.715 132.365 ;
        RECT 54.360 130.665 54.615 131.235 ;
        RECT 54.785 131.065 55.715 131.235 ;
        RECT 55.885 132.025 56.895 132.195 ;
        RECT 55.885 131.225 56.055 132.025 ;
        RECT 56.260 131.685 56.535 131.825 ;
        RECT 56.255 131.515 56.535 131.685 ;
        RECT 55.540 131.030 55.715 131.065 ;
        RECT 54.785 130.495 55.115 130.895 ;
        RECT 55.540 130.665 56.070 131.030 ;
        RECT 56.260 130.665 56.535 131.515 ;
        RECT 56.705 130.665 56.895 132.025 ;
        RECT 57.065 132.040 57.235 132.705 ;
        RECT 57.405 132.285 57.575 133.045 ;
        RECT 57.810 132.285 58.325 132.695 ;
        RECT 58.495 132.610 63.840 133.045 ;
        RECT 57.065 131.850 57.815 132.040 ;
        RECT 57.985 131.475 58.325 132.285 ;
        RECT 57.095 131.305 58.325 131.475 ;
        RECT 57.075 130.495 57.585 131.030 ;
        RECT 57.805 130.700 58.050 131.305 ;
        RECT 60.080 131.040 60.420 131.870 ;
        RECT 61.900 131.360 62.250 132.610 ;
        RECT 64.015 131.955 66.605 133.045 ;
        RECT 64.015 131.265 65.225 131.785 ;
        RECT 65.395 131.435 66.605 131.955 ;
        RECT 67.235 131.880 67.525 133.045 ;
        RECT 68.165 132.325 68.495 133.045 ;
        RECT 68.665 132.155 68.835 132.875 ;
        RECT 69.005 132.325 69.335 133.045 ;
        RECT 69.505 132.155 69.675 132.875 ;
        RECT 69.845 132.665 70.175 133.045 ;
        RECT 70.345 132.515 70.515 132.875 ;
        RECT 70.820 132.685 72.600 132.855 ;
        RECT 70.345 132.345 72.060 132.515 ;
        RECT 72.250 132.345 72.600 132.685 ;
        RECT 72.770 132.245 73.075 133.045 ;
        RECT 68.160 131.985 69.675 132.155 ;
        RECT 69.855 132.175 70.025 132.195 ;
        RECT 69.855 132.005 71.610 132.175 ;
        RECT 73.245 132.075 73.500 132.875 ;
        RECT 58.495 130.495 63.840 131.040 ;
        RECT 64.015 130.495 66.605 131.265 ;
        RECT 67.235 130.495 67.525 131.220 ;
        RECT 68.160 131.215 68.390 131.985 ;
        RECT 69.855 131.655 70.025 132.005 ;
        RECT 68.560 131.485 70.025 131.655 ;
        RECT 69.855 131.235 70.025 131.485 ;
        RECT 70.195 131.405 70.910 131.735 ;
        RECT 71.155 131.405 71.625 131.735 ;
        RECT 71.840 131.405 72.110 132.025 ;
        RECT 72.510 131.905 73.500 132.075 ;
        RECT 72.510 131.405 72.680 131.905 ;
        RECT 72.850 131.405 73.160 131.735 ;
        RECT 68.160 131.045 69.675 131.215 ;
        RECT 69.855 131.065 70.530 131.235 ;
        RECT 68.165 130.495 68.495 130.875 ;
        RECT 68.665 130.665 68.835 131.045 ;
        RECT 69.005 130.495 69.335 130.875 ;
        RECT 69.505 130.665 69.675 131.045 ;
        RECT 70.360 130.875 70.530 131.065 ;
        RECT 70.740 131.215 70.910 131.405 ;
        RECT 72.850 131.215 73.020 131.405 ;
        RECT 70.740 131.045 73.020 131.215 ;
        RECT 73.330 131.035 73.500 131.905 ;
        RECT 69.845 130.495 70.175 130.875 ;
        RECT 70.360 130.705 71.615 130.875 ;
        RECT 72.745 130.495 73.075 130.875 ;
        RECT 73.245 130.705 73.500 131.035 ;
        RECT 73.680 131.905 73.955 132.875 ;
        RECT 74.165 132.245 74.445 133.045 ;
        RECT 74.615 132.535 75.805 132.825 ;
        RECT 74.615 132.195 75.785 132.365 ;
        RECT 74.615 132.075 74.785 132.195 ;
        RECT 74.125 131.905 74.785 132.075 ;
        RECT 73.680 131.170 73.850 131.905 ;
        RECT 74.125 131.735 74.295 131.905 ;
        RECT 75.095 131.735 75.290 132.025 ;
        RECT 75.460 131.905 75.785 132.195 ;
        RECT 76.140 132.135 76.390 132.865 ;
        RECT 76.560 132.315 76.890 133.045 ;
        RECT 77.060 132.135 77.245 132.865 ;
        RECT 76.140 131.935 77.245 132.135 ;
        RECT 77.415 131.735 77.645 132.865 ;
        RECT 77.825 132.195 78.550 132.865 ;
        RECT 74.020 131.405 74.295 131.735 ;
        RECT 74.465 131.405 75.290 131.735 ;
        RECT 75.460 131.405 75.805 131.735 ;
        RECT 74.125 131.235 74.295 131.405 ;
        RECT 73.680 130.825 73.955 131.170 ;
        RECT 74.125 131.065 75.790 131.235 ;
        RECT 75.985 131.175 76.325 131.735 ;
        RECT 76.495 131.405 77.135 131.735 ;
        RECT 77.315 131.405 77.645 131.735 ;
        RECT 77.825 131.405 78.125 132.025 ;
        RECT 74.145 130.495 74.525 130.895 ;
        RECT 74.695 130.715 74.865 131.065 ;
        RECT 75.035 130.495 75.365 130.895 ;
        RECT 75.535 130.715 75.790 131.065 ;
        RECT 75.975 130.495 76.315 131.005 ;
        RECT 76.495 130.675 76.745 131.405 ;
        RECT 78.335 131.225 78.550 132.195 ;
        RECT 78.735 131.955 80.405 133.045 ;
        RECT 77.070 131.035 78.550 131.225 ;
        RECT 78.735 131.265 79.485 131.785 ;
        RECT 79.655 131.435 80.405 131.955 ;
        RECT 77.070 130.675 77.255 131.035 ;
        RECT 77.435 130.495 77.765 130.865 ;
        RECT 77.945 130.675 78.170 131.035 ;
        RECT 78.735 130.495 80.405 131.265 ;
        RECT 81.050 130.675 81.330 132.865 ;
        RECT 81.520 131.905 81.805 133.045 ;
        RECT 82.070 132.395 82.240 132.865 ;
        RECT 82.415 132.565 82.745 133.045 ;
        RECT 82.915 132.395 83.095 132.865 ;
        RECT 82.070 132.195 83.095 132.395 ;
        RECT 81.530 131.225 81.790 131.735 ;
        RECT 82.000 131.405 82.260 132.025 ;
        RECT 82.455 131.405 82.880 132.025 ;
        RECT 83.265 131.755 83.595 132.865 ;
        RECT 83.765 132.635 84.115 133.045 ;
        RECT 84.285 132.455 84.525 132.845 ;
        RECT 83.050 131.455 83.595 131.755 ;
        RECT 83.775 132.255 84.525 132.455 ;
        RECT 83.775 131.575 84.115 132.255 ;
        RECT 83.050 131.225 83.270 131.455 ;
        RECT 81.530 131.035 83.270 131.225 ;
        RECT 81.530 130.495 82.260 130.865 ;
        RECT 82.840 130.675 83.270 131.035 ;
        RECT 83.440 130.495 83.685 131.275 ;
        RECT 83.885 130.675 84.115 131.575 ;
        RECT 84.295 130.735 84.525 132.075 ;
        RECT 84.715 131.905 84.975 133.045 ;
        RECT 85.145 131.895 85.475 132.875 ;
        RECT 85.645 131.905 85.925 133.045 ;
        RECT 86.095 131.955 88.685 133.045 ;
        RECT 84.735 131.485 85.070 131.735 ;
        RECT 85.240 131.295 85.410 131.895 ;
        RECT 85.580 131.465 85.915 131.735 ;
        RECT 84.715 130.665 85.410 131.295 ;
        RECT 85.615 130.495 85.925 131.295 ;
        RECT 86.095 131.265 87.305 131.785 ;
        RECT 87.475 131.435 88.685 131.955 ;
        RECT 88.860 132.690 89.940 132.860 ;
        RECT 88.860 131.905 89.195 132.690 ;
        RECT 89.365 131.735 89.600 132.415 ;
        RECT 89.770 132.075 89.940 132.690 ;
        RECT 90.205 132.245 90.520 133.045 ;
        RECT 89.770 131.905 90.085 132.075 ;
        RECT 88.860 131.405 89.195 131.735 ;
        RECT 89.365 131.405 89.745 131.735 ;
        RECT 86.095 130.495 88.685 131.265 ;
        RECT 89.915 131.235 90.085 131.905 ;
        RECT 88.860 131.065 90.085 131.235 ;
        RECT 90.255 131.065 90.525 132.075 ;
        RECT 90.695 131.955 92.365 133.045 ;
        RECT 90.695 131.265 91.445 131.785 ;
        RECT 91.615 131.435 92.365 131.955 ;
        RECT 92.995 131.880 93.285 133.045 ;
        RECT 93.455 131.955 94.665 133.045 ;
        RECT 88.860 130.795 89.115 131.065 ;
        RECT 89.285 130.495 89.615 130.895 ;
        RECT 89.785 130.795 89.955 131.065 ;
        RECT 90.125 130.495 90.455 130.895 ;
        RECT 90.695 130.495 92.365 131.265 ;
        RECT 93.455 131.245 93.975 131.785 ;
        RECT 94.145 131.415 94.665 131.955 ;
        RECT 94.840 132.095 95.105 132.865 ;
        RECT 95.275 132.325 95.605 133.045 ;
        RECT 95.795 132.505 96.055 132.865 ;
        RECT 96.225 132.675 96.555 133.045 ;
        RECT 96.725 132.505 96.985 132.865 ;
        RECT 95.795 132.275 96.985 132.505 ;
        RECT 97.555 132.095 97.845 132.865 ;
        RECT 92.995 130.495 93.285 131.220 ;
        RECT 93.455 130.495 94.665 131.245 ;
        RECT 94.840 130.675 95.175 132.095 ;
        RECT 95.350 131.915 97.845 132.095 ;
        RECT 98.055 131.955 99.265 133.045 ;
        RECT 95.350 131.225 95.575 131.915 ;
        RECT 95.775 131.405 96.055 131.735 ;
        RECT 96.235 131.405 96.810 131.735 ;
        RECT 96.990 131.405 97.425 131.735 ;
        RECT 97.605 131.405 97.875 131.735 ;
        RECT 98.055 131.245 98.575 131.785 ;
        RECT 98.745 131.415 99.265 131.955 ;
        RECT 99.440 132.095 99.705 132.865 ;
        RECT 99.875 132.325 100.205 133.045 ;
        RECT 100.395 132.505 100.655 132.865 ;
        RECT 100.825 132.675 101.155 133.045 ;
        RECT 101.325 132.505 101.585 132.865 ;
        RECT 100.395 132.275 101.585 132.505 ;
        RECT 102.155 132.095 102.445 132.865 ;
        RECT 95.350 131.035 97.835 131.225 ;
        RECT 95.355 130.495 96.100 130.865 ;
        RECT 96.665 130.675 96.920 131.035 ;
        RECT 97.100 130.495 97.430 130.865 ;
        RECT 97.610 130.675 97.835 131.035 ;
        RECT 98.055 130.495 99.265 131.245 ;
        RECT 99.440 130.675 99.775 132.095 ;
        RECT 99.950 131.915 102.445 132.095 ;
        RECT 102.655 131.955 103.865 133.045 ;
        RECT 99.950 131.225 100.175 131.915 ;
        RECT 100.375 131.405 100.655 131.735 ;
        RECT 100.835 131.405 101.410 131.735 ;
        RECT 101.590 131.405 102.025 131.735 ;
        RECT 102.205 131.405 102.475 131.735 ;
        RECT 102.655 131.245 103.175 131.785 ;
        RECT 103.345 131.415 103.865 131.955 ;
        RECT 104.125 132.035 104.295 132.875 ;
        RECT 104.465 132.705 105.635 132.875 ;
        RECT 104.465 132.205 104.795 132.705 ;
        RECT 105.305 132.665 105.635 132.705 ;
        RECT 105.825 132.625 106.180 133.045 ;
        RECT 104.965 132.445 105.195 132.535 ;
        RECT 106.350 132.445 106.600 132.875 ;
        RECT 104.965 132.205 106.600 132.445 ;
        RECT 106.770 132.285 107.100 133.045 ;
        RECT 107.270 132.205 107.525 132.875 ;
        RECT 104.125 131.865 107.185 132.035 ;
        RECT 104.040 131.485 104.390 131.695 ;
        RECT 104.560 131.485 105.005 131.685 ;
        RECT 105.175 131.485 105.650 131.685 ;
        RECT 99.950 131.035 102.435 131.225 ;
        RECT 99.955 130.495 100.700 130.865 ;
        RECT 101.265 130.675 101.520 131.035 ;
        RECT 101.700 130.495 102.030 130.865 ;
        RECT 102.210 130.675 102.435 131.035 ;
        RECT 102.655 130.495 103.865 131.245 ;
        RECT 104.125 131.145 105.190 131.315 ;
        RECT 104.125 130.665 104.295 131.145 ;
        RECT 104.465 130.495 104.795 130.975 ;
        RECT 105.020 130.915 105.190 131.145 ;
        RECT 105.370 131.085 105.650 131.485 ;
        RECT 105.920 131.485 106.250 131.685 ;
        RECT 106.420 131.485 106.785 131.685 ;
        RECT 105.920 131.085 106.205 131.485 ;
        RECT 107.015 131.315 107.185 131.865 ;
        RECT 106.385 131.145 107.185 131.315 ;
        RECT 106.385 130.915 106.555 131.145 ;
        RECT 107.355 131.075 107.525 132.205 ;
        RECT 107.340 131.005 107.525 131.075 ;
        RECT 107.315 130.995 107.525 131.005 ;
        RECT 105.020 130.665 106.555 130.915 ;
        RECT 106.725 130.495 107.055 130.975 ;
        RECT 107.270 130.665 107.525 130.995 ;
        RECT 107.715 131.440 107.995 132.875 ;
        RECT 108.165 132.270 108.875 133.045 ;
        RECT 109.045 132.100 109.375 132.875 ;
        RECT 108.225 131.885 109.375 132.100 ;
        RECT 107.715 130.665 108.055 131.440 ;
        RECT 108.225 131.315 108.510 131.885 ;
        RECT 108.695 131.485 109.165 131.715 ;
        RECT 109.570 131.685 109.785 132.800 ;
        RECT 109.965 132.325 110.295 133.045 ;
        RECT 110.075 131.685 110.305 132.025 ;
        RECT 110.475 131.955 111.685 133.045 ;
        RECT 112.055 132.375 112.335 133.045 ;
        RECT 112.505 132.155 112.805 132.705 ;
        RECT 113.005 132.325 113.335 133.045 ;
        RECT 113.525 132.325 113.985 132.875 ;
        RECT 109.335 131.505 109.785 131.685 ;
        RECT 109.335 131.485 109.665 131.505 ;
        RECT 109.975 131.485 110.305 131.685 ;
        RECT 108.225 131.125 108.935 131.315 ;
        RECT 108.635 130.985 108.935 131.125 ;
        RECT 109.125 131.125 110.305 131.315 ;
        RECT 109.125 131.045 109.455 131.125 ;
        RECT 108.635 130.975 108.950 130.985 ;
        RECT 108.635 130.965 108.960 130.975 ;
        RECT 108.635 130.960 108.970 130.965 ;
        RECT 108.225 130.495 108.395 130.955 ;
        RECT 108.635 130.950 108.975 130.960 ;
        RECT 108.635 130.945 108.980 130.950 ;
        RECT 108.635 130.935 108.985 130.945 ;
        RECT 108.635 130.930 108.990 130.935 ;
        RECT 108.635 130.665 108.995 130.930 ;
        RECT 109.625 130.495 109.795 130.955 ;
        RECT 109.965 130.665 110.305 131.125 ;
        RECT 110.475 131.245 110.995 131.785 ;
        RECT 111.165 131.415 111.685 131.955 ;
        RECT 111.870 131.735 112.135 132.095 ;
        RECT 112.505 131.985 113.445 132.155 ;
        RECT 113.275 131.735 113.445 131.985 ;
        RECT 111.870 131.485 112.545 131.735 ;
        RECT 112.765 131.485 113.105 131.735 ;
        RECT 113.275 131.405 113.565 131.735 ;
        RECT 113.275 131.315 113.445 131.405 ;
        RECT 110.475 130.495 111.685 131.245 ;
        RECT 112.055 131.125 113.445 131.315 ;
        RECT 112.055 130.765 112.385 131.125 ;
        RECT 113.735 130.955 113.985 132.325 ;
        RECT 114.365 132.065 114.695 132.875 ;
        RECT 114.865 132.235 115.035 133.045 ;
        RECT 115.205 132.065 115.535 132.875 ;
        RECT 115.705 132.235 115.875 133.045 ;
        RECT 116.045 132.705 118.155 132.875 ;
        RECT 116.045 132.065 116.295 132.705 ;
        RECT 114.365 131.895 116.295 132.065 ;
        RECT 116.510 132.065 116.895 132.535 ;
        RECT 117.065 132.235 117.235 132.705 ;
        RECT 117.405 132.065 117.735 132.535 ;
        RECT 117.905 132.235 118.155 132.705 ;
        RECT 118.325 132.065 118.575 132.875 ;
        RECT 116.510 131.895 118.575 132.065 ;
        RECT 114.170 131.515 115.305 131.685 ;
        RECT 114.170 131.485 115.280 131.515 ;
        RECT 115.570 131.485 116.225 131.685 ;
        RECT 113.005 130.495 113.255 130.955 ;
        RECT 113.425 130.665 113.985 130.955 ;
        RECT 114.295 131.090 115.455 131.260 ;
        RECT 116.510 131.255 116.800 131.895 ;
        RECT 118.755 131.880 119.045 133.045 ;
        RECT 119.215 131.905 119.490 132.875 ;
        RECT 119.700 132.245 119.980 133.045 ;
        RECT 120.150 132.535 121.765 132.865 ;
        RECT 120.150 132.195 121.325 132.365 ;
        RECT 120.150 132.075 120.320 132.195 ;
        RECT 119.660 131.905 120.320 132.075 ;
        RECT 116.970 131.515 117.605 131.685 ;
        RECT 117.890 131.515 118.525 131.685 ;
        RECT 116.970 131.485 117.600 131.515 ;
        RECT 117.890 131.485 118.520 131.515 ;
        RECT 114.295 130.665 114.615 131.090 ;
        RECT 114.785 130.495 115.115 130.920 ;
        RECT 115.285 130.915 115.455 131.090 ;
        RECT 115.625 131.085 117.315 131.255 ;
        RECT 117.485 131.090 118.575 131.260 ;
        RECT 117.485 130.915 117.655 131.090 ;
        RECT 115.285 130.665 116.375 130.915 ;
        RECT 116.565 130.665 117.655 130.915 ;
        RECT 117.825 130.495 118.155 130.920 ;
        RECT 118.325 130.665 118.575 131.090 ;
        RECT 118.755 130.495 119.045 131.220 ;
        RECT 119.215 131.170 119.385 131.905 ;
        RECT 119.660 131.735 119.830 131.905 ;
        RECT 120.580 131.735 120.825 132.025 ;
        RECT 120.995 131.905 121.325 132.195 ;
        RECT 121.585 131.735 121.755 132.295 ;
        RECT 122.005 131.905 122.265 133.045 ;
        RECT 122.435 131.955 123.645 133.045 ;
        RECT 119.555 131.405 119.830 131.735 ;
        RECT 120.000 131.405 120.825 131.735 ;
        RECT 121.040 131.405 121.755 131.735 ;
        RECT 121.925 131.485 122.260 131.735 ;
        RECT 119.660 131.235 119.830 131.405 ;
        RECT 121.505 131.315 121.755 131.405 ;
        RECT 119.215 130.825 119.490 131.170 ;
        RECT 119.660 131.065 121.325 131.235 ;
        RECT 119.680 130.495 120.055 130.895 ;
        RECT 120.225 130.715 120.395 131.065 ;
        RECT 120.565 130.495 120.895 130.895 ;
        RECT 121.065 130.665 121.325 131.065 ;
        RECT 121.505 130.895 121.835 131.315 ;
        RECT 122.005 130.495 122.265 131.315 ;
        RECT 122.435 131.245 122.955 131.785 ;
        RECT 123.125 131.415 123.645 131.955 ;
        RECT 122.435 130.495 123.645 131.245 ;
        RECT 123.830 130.675 124.110 132.865 ;
        RECT 124.300 131.905 124.585 133.045 ;
        RECT 124.850 132.395 125.020 132.865 ;
        RECT 125.195 132.565 125.525 133.045 ;
        RECT 125.695 132.395 125.875 132.865 ;
        RECT 124.850 132.195 125.875 132.395 ;
        RECT 124.310 131.225 124.570 131.735 ;
        RECT 124.780 131.405 125.040 132.025 ;
        RECT 125.235 131.405 125.660 132.025 ;
        RECT 126.045 131.755 126.375 132.865 ;
        RECT 126.545 132.635 126.895 133.045 ;
        RECT 127.065 132.455 127.305 132.845 ;
        RECT 125.830 131.455 126.375 131.755 ;
        RECT 126.555 132.255 127.305 132.455 ;
        RECT 126.555 131.575 126.895 132.255 ;
        RECT 125.830 131.225 126.050 131.455 ;
        RECT 124.310 131.035 126.050 131.225 ;
        RECT 124.310 130.495 125.040 130.865 ;
        RECT 125.620 130.675 126.050 131.035 ;
        RECT 126.220 130.495 126.465 131.275 ;
        RECT 126.665 130.675 126.895 131.575 ;
        RECT 127.075 130.735 127.305 132.075 ;
        RECT 127.505 131.905 127.835 133.045 ;
        RECT 128.365 132.075 128.695 132.860 ;
        RECT 128.885 132.325 129.215 133.045 ;
        RECT 128.015 131.905 128.695 132.075 ;
        RECT 127.495 131.485 127.845 131.735 ;
        RECT 128.015 131.305 128.185 131.905 ;
        RECT 128.355 131.485 128.705 131.735 ;
        RECT 128.875 131.685 129.105 132.025 ;
        RECT 129.395 131.685 129.610 132.800 ;
        RECT 129.805 132.100 130.135 132.875 ;
        RECT 130.305 132.270 131.015 133.045 ;
        RECT 129.805 131.885 130.955 132.100 ;
        RECT 128.875 131.485 129.205 131.685 ;
        RECT 129.395 131.505 129.845 131.685 ;
        RECT 129.515 131.485 129.845 131.505 ;
        RECT 130.015 131.485 130.485 131.715 ;
        RECT 130.670 131.315 130.955 131.885 ;
        RECT 131.185 131.440 131.465 132.875 ;
        RECT 127.505 130.495 127.775 131.305 ;
        RECT 127.945 130.665 128.275 131.305 ;
        RECT 128.445 130.495 128.685 131.305 ;
        RECT 128.875 131.125 130.055 131.315 ;
        RECT 128.875 130.665 129.215 131.125 ;
        RECT 129.725 131.045 130.055 131.125 ;
        RECT 130.245 131.125 130.955 131.315 ;
        RECT 130.245 130.985 130.545 131.125 ;
        RECT 130.230 130.975 130.545 130.985 ;
        RECT 130.220 130.965 130.545 130.975 ;
        RECT 130.210 130.960 130.545 130.965 ;
        RECT 129.385 130.495 129.555 130.955 ;
        RECT 130.205 130.950 130.545 130.960 ;
        RECT 130.200 130.945 130.545 130.950 ;
        RECT 130.195 130.935 130.545 130.945 ;
        RECT 130.190 130.930 130.545 130.935 ;
        RECT 130.185 130.665 130.545 130.930 ;
        RECT 130.785 130.495 130.955 130.955 ;
        RECT 131.125 130.665 131.465 131.440 ;
        RECT 131.655 132.205 131.910 132.875 ;
        RECT 132.080 132.285 132.410 133.045 ;
        RECT 132.580 132.445 132.830 132.875 ;
        RECT 133.000 132.625 133.355 133.045 ;
        RECT 133.545 132.705 134.715 132.875 ;
        RECT 133.545 132.665 133.875 132.705 ;
        RECT 133.985 132.445 134.215 132.535 ;
        RECT 132.580 132.205 134.215 132.445 ;
        RECT 134.385 132.205 134.715 132.705 ;
        RECT 131.655 132.195 131.865 132.205 ;
        RECT 131.655 131.075 131.825 132.195 ;
        RECT 134.885 132.035 135.055 132.875 ;
        RECT 131.995 131.865 135.055 132.035 ;
        RECT 135.355 132.095 135.645 132.865 ;
        RECT 136.215 132.505 136.475 132.865 ;
        RECT 136.645 132.675 136.975 133.045 ;
        RECT 137.145 132.505 137.405 132.865 ;
        RECT 136.215 132.275 137.405 132.505 ;
        RECT 137.595 132.325 137.925 133.045 ;
        RECT 138.095 132.095 138.360 132.865 ;
        RECT 135.355 131.915 137.850 132.095 ;
        RECT 131.995 131.315 132.165 131.865 ;
        RECT 132.395 131.485 132.760 131.685 ;
        RECT 132.930 131.485 133.260 131.685 ;
        RECT 131.995 131.145 132.795 131.315 ;
        RECT 131.655 130.995 131.840 131.075 ;
        RECT 131.655 130.665 131.910 130.995 ;
        RECT 132.125 130.495 132.455 130.975 ;
        RECT 132.625 130.915 132.795 131.145 ;
        RECT 132.975 131.085 133.260 131.485 ;
        RECT 133.530 131.485 134.005 131.685 ;
        RECT 134.175 131.485 134.620 131.685 ;
        RECT 134.790 131.485 135.140 131.695 ;
        RECT 133.530 131.085 133.810 131.485 ;
        RECT 135.325 131.405 135.595 131.735 ;
        RECT 135.775 131.405 136.210 131.735 ;
        RECT 136.390 131.405 136.965 131.735 ;
        RECT 137.145 131.405 137.425 131.735 ;
        RECT 133.990 131.145 135.055 131.315 ;
        RECT 137.625 131.225 137.850 131.915 ;
        RECT 133.990 130.915 134.160 131.145 ;
        RECT 132.625 130.665 134.160 130.915 ;
        RECT 134.385 130.495 134.715 130.975 ;
        RECT 134.885 130.665 135.055 131.145 ;
        RECT 135.365 131.035 137.850 131.225 ;
        RECT 135.365 130.675 135.590 131.035 ;
        RECT 135.770 130.495 136.100 130.865 ;
        RECT 136.280 130.675 136.535 131.035 ;
        RECT 137.100 130.495 137.845 130.865 ;
        RECT 138.025 130.675 138.360 132.095 ;
        RECT 138.700 132.135 138.950 132.865 ;
        RECT 139.120 132.315 139.450 133.045 ;
        RECT 139.620 132.135 139.805 132.865 ;
        RECT 138.700 131.935 139.805 132.135 ;
        RECT 139.975 131.735 140.205 132.865 ;
        RECT 140.385 132.195 141.110 132.865 ;
        RECT 138.545 131.175 138.885 131.735 ;
        RECT 139.055 131.405 139.695 131.735 ;
        RECT 139.875 131.405 140.205 131.735 ;
        RECT 140.385 131.405 140.685 132.025 ;
        RECT 138.535 130.495 138.875 131.005 ;
        RECT 139.055 130.675 139.305 131.405 ;
        RECT 140.895 131.225 141.110 132.195 ;
        RECT 141.295 131.955 143.885 133.045 ;
        RECT 139.630 131.035 141.110 131.225 ;
        RECT 141.295 131.265 142.505 131.785 ;
        RECT 142.675 131.435 143.885 131.955 ;
        RECT 144.515 131.880 144.805 133.045 ;
        RECT 144.975 132.610 150.320 133.045 ;
        RECT 150.495 132.610 155.840 133.045 ;
        RECT 139.630 130.675 139.815 131.035 ;
        RECT 139.995 130.495 140.325 130.865 ;
        RECT 140.505 130.675 140.730 131.035 ;
        RECT 141.295 130.495 143.885 131.265 ;
        RECT 144.515 130.495 144.805 131.220 ;
        RECT 146.560 131.040 146.900 131.870 ;
        RECT 148.380 131.360 148.730 132.610 ;
        RECT 152.080 131.040 152.420 131.870 ;
        RECT 153.900 131.360 154.250 132.610 ;
        RECT 156.935 131.955 158.145 133.045 ;
        RECT 156.935 131.415 157.455 131.955 ;
        RECT 157.625 131.245 158.145 131.785 ;
        RECT 144.975 130.495 150.320 131.040 ;
        RECT 150.495 130.495 155.840 131.040 ;
        RECT 156.935 130.495 158.145 131.245 ;
        RECT 2.750 130.325 158.230 130.495 ;
        RECT 2.835 129.575 4.045 130.325 ;
        RECT 2.835 129.035 3.355 129.575 ;
        RECT 4.215 129.555 6.805 130.325 ;
        RECT 7.435 129.650 7.695 130.155 ;
        RECT 7.875 129.945 8.205 130.325 ;
        RECT 8.385 129.775 8.555 130.155 ;
        RECT 3.525 128.865 4.045 129.405 ;
        RECT 4.215 129.035 5.425 129.555 ;
        RECT 5.595 128.865 6.805 129.385 ;
        RECT 2.835 127.775 4.045 128.865 ;
        RECT 4.215 127.775 6.805 128.865 ;
        RECT 7.435 128.850 7.605 129.650 ;
        RECT 7.890 129.605 8.555 129.775 ;
        RECT 7.890 129.350 8.060 129.605 ;
        RECT 8.815 129.575 10.025 130.325 ;
        RECT 10.200 129.775 10.455 130.065 ;
        RECT 10.625 129.945 10.955 130.325 ;
        RECT 10.200 129.605 10.950 129.775 ;
        RECT 7.775 129.020 8.060 129.350 ;
        RECT 8.295 129.055 8.625 129.425 ;
        RECT 8.815 129.035 9.335 129.575 ;
        RECT 7.890 128.875 8.060 129.020 ;
        RECT 7.435 127.945 7.705 128.850 ;
        RECT 7.890 128.705 8.555 128.875 ;
        RECT 9.505 128.865 10.025 129.405 ;
        RECT 7.875 127.775 8.205 128.535 ;
        RECT 8.385 127.945 8.555 128.705 ;
        RECT 8.815 127.775 10.025 128.865 ;
        RECT 10.200 128.785 10.550 129.435 ;
        RECT 10.720 128.615 10.950 129.605 ;
        RECT 10.200 128.445 10.950 128.615 ;
        RECT 10.200 127.945 10.455 128.445 ;
        RECT 10.625 127.775 10.955 128.275 ;
        RECT 11.125 127.945 11.295 130.065 ;
        RECT 11.655 129.965 11.985 130.325 ;
        RECT 12.155 129.935 12.650 130.105 ;
        RECT 12.855 129.935 13.710 130.105 ;
        RECT 11.525 128.745 11.985 129.795 ;
        RECT 11.465 127.960 11.790 128.745 ;
        RECT 12.155 128.575 12.325 129.935 ;
        RECT 12.495 129.025 12.845 129.645 ;
        RECT 13.015 129.425 13.370 129.645 ;
        RECT 13.015 128.835 13.185 129.425 ;
        RECT 13.540 129.225 13.710 129.935 ;
        RECT 14.585 129.865 14.915 130.325 ;
        RECT 15.125 129.965 15.475 130.135 ;
        RECT 13.915 129.395 14.705 129.645 ;
        RECT 15.125 129.575 15.385 129.965 ;
        RECT 15.695 129.875 16.645 130.155 ;
        RECT 16.815 129.885 17.005 130.325 ;
        RECT 17.175 129.945 18.245 130.115 ;
        RECT 14.875 129.225 15.045 129.405 ;
        RECT 12.155 128.405 12.550 128.575 ;
        RECT 12.720 128.445 13.185 128.835 ;
        RECT 13.355 129.055 15.045 129.225 ;
        RECT 12.380 128.275 12.550 128.405 ;
        RECT 13.355 128.275 13.525 129.055 ;
        RECT 15.215 128.885 15.385 129.575 ;
        RECT 13.885 128.715 15.385 128.885 ;
        RECT 15.575 128.915 15.785 129.705 ;
        RECT 15.955 129.085 16.305 129.705 ;
        RECT 16.475 129.095 16.645 129.875 ;
        RECT 17.175 129.715 17.345 129.945 ;
        RECT 16.815 129.545 17.345 129.715 ;
        RECT 16.815 129.265 17.035 129.545 ;
        RECT 17.515 129.375 17.755 129.775 ;
        RECT 16.475 128.925 16.880 129.095 ;
        RECT 17.215 129.005 17.755 129.375 ;
        RECT 17.925 129.590 18.245 129.945 ;
        RECT 18.490 129.865 18.795 130.325 ;
        RECT 18.965 129.615 19.220 130.145 ;
        RECT 17.925 129.415 18.250 129.590 ;
        RECT 17.925 129.115 18.840 129.415 ;
        RECT 18.100 129.085 18.840 129.115 ;
        RECT 15.575 128.755 16.250 128.915 ;
        RECT 16.710 128.835 16.880 128.925 ;
        RECT 15.575 128.745 16.540 128.755 ;
        RECT 15.215 128.575 15.385 128.715 ;
        RECT 11.960 127.775 12.210 128.235 ;
        RECT 12.380 127.945 12.630 128.275 ;
        RECT 12.845 127.945 13.525 128.275 ;
        RECT 13.695 128.375 14.770 128.545 ;
        RECT 15.215 128.405 15.775 128.575 ;
        RECT 16.080 128.455 16.540 128.745 ;
        RECT 16.710 128.665 17.930 128.835 ;
        RECT 13.695 128.035 13.865 128.375 ;
        RECT 14.100 127.775 14.430 128.205 ;
        RECT 14.600 128.035 14.770 128.375 ;
        RECT 15.065 127.775 15.435 128.235 ;
        RECT 15.605 127.945 15.775 128.405 ;
        RECT 16.710 128.285 16.880 128.665 ;
        RECT 18.100 128.495 18.270 129.085 ;
        RECT 19.010 128.965 19.220 129.615 ;
        RECT 19.400 129.775 19.655 130.065 ;
        RECT 19.825 129.945 20.155 130.325 ;
        RECT 19.400 129.605 20.150 129.775 ;
        RECT 16.010 127.945 16.880 128.285 ;
        RECT 17.470 128.325 18.270 128.495 ;
        RECT 17.050 127.775 17.300 128.235 ;
        RECT 17.470 128.035 17.640 128.325 ;
        RECT 17.820 127.775 18.150 128.155 ;
        RECT 18.490 127.775 18.795 128.915 ;
        RECT 18.965 128.085 19.220 128.965 ;
        RECT 19.400 128.785 19.750 129.435 ;
        RECT 19.920 128.615 20.150 129.605 ;
        RECT 19.400 128.445 20.150 128.615 ;
        RECT 19.400 127.945 19.655 128.445 ;
        RECT 19.825 127.775 20.155 128.275 ;
        RECT 20.325 127.945 20.495 130.065 ;
        RECT 20.855 129.965 21.185 130.325 ;
        RECT 21.355 129.935 21.850 130.105 ;
        RECT 22.055 129.935 22.910 130.105 ;
        RECT 20.725 128.745 21.185 129.795 ;
        RECT 20.665 127.960 20.990 128.745 ;
        RECT 21.355 128.575 21.525 129.935 ;
        RECT 21.695 129.025 22.045 129.645 ;
        RECT 22.215 129.425 22.570 129.645 ;
        RECT 22.215 128.835 22.385 129.425 ;
        RECT 22.740 129.225 22.910 129.935 ;
        RECT 23.785 129.865 24.115 130.325 ;
        RECT 24.325 129.965 24.675 130.135 ;
        RECT 23.115 129.395 23.905 129.645 ;
        RECT 24.325 129.575 24.585 129.965 ;
        RECT 24.895 129.875 25.845 130.155 ;
        RECT 26.015 129.885 26.205 130.325 ;
        RECT 26.375 129.945 27.445 130.115 ;
        RECT 24.075 129.225 24.245 129.405 ;
        RECT 21.355 128.405 21.750 128.575 ;
        RECT 21.920 128.445 22.385 128.835 ;
        RECT 22.555 129.055 24.245 129.225 ;
        RECT 21.580 128.275 21.750 128.405 ;
        RECT 22.555 128.275 22.725 129.055 ;
        RECT 24.415 128.885 24.585 129.575 ;
        RECT 23.085 128.715 24.585 128.885 ;
        RECT 24.775 128.915 24.985 129.705 ;
        RECT 25.155 129.085 25.505 129.705 ;
        RECT 25.675 129.095 25.845 129.875 ;
        RECT 26.375 129.715 26.545 129.945 ;
        RECT 26.015 129.545 26.545 129.715 ;
        RECT 26.015 129.265 26.235 129.545 ;
        RECT 26.715 129.375 26.955 129.775 ;
        RECT 25.675 128.925 26.080 129.095 ;
        RECT 26.415 129.005 26.955 129.375 ;
        RECT 27.125 129.590 27.445 129.945 ;
        RECT 27.690 129.865 27.995 130.325 ;
        RECT 28.165 129.615 28.420 130.145 ;
        RECT 27.125 129.415 27.450 129.590 ;
        RECT 27.125 129.115 28.040 129.415 ;
        RECT 27.300 129.085 28.040 129.115 ;
        RECT 24.775 128.755 25.450 128.915 ;
        RECT 25.910 128.835 26.080 128.925 ;
        RECT 24.775 128.745 25.740 128.755 ;
        RECT 24.415 128.575 24.585 128.715 ;
        RECT 21.160 127.775 21.410 128.235 ;
        RECT 21.580 127.945 21.830 128.275 ;
        RECT 22.045 127.945 22.725 128.275 ;
        RECT 22.895 128.375 23.970 128.545 ;
        RECT 24.415 128.405 24.975 128.575 ;
        RECT 25.280 128.455 25.740 128.745 ;
        RECT 25.910 128.665 27.130 128.835 ;
        RECT 22.895 128.035 23.065 128.375 ;
        RECT 23.300 127.775 23.630 128.205 ;
        RECT 23.800 128.035 23.970 128.375 ;
        RECT 24.265 127.775 24.635 128.235 ;
        RECT 24.805 127.945 24.975 128.405 ;
        RECT 25.910 128.285 26.080 128.665 ;
        RECT 27.300 128.495 27.470 129.085 ;
        RECT 28.210 128.965 28.420 129.615 ;
        RECT 28.595 129.600 28.885 130.325 ;
        RECT 30.065 129.775 30.235 130.155 ;
        RECT 30.415 129.945 30.745 130.325 ;
        RECT 30.065 129.605 30.730 129.775 ;
        RECT 30.925 129.650 31.185 130.155 ;
        RECT 29.995 129.055 30.325 129.425 ;
        RECT 30.560 129.350 30.730 129.605 ;
        RECT 25.210 127.945 26.080 128.285 ;
        RECT 26.670 128.325 27.470 128.495 ;
        RECT 26.250 127.775 26.500 128.235 ;
        RECT 26.670 128.035 26.840 128.325 ;
        RECT 27.020 127.775 27.350 128.155 ;
        RECT 27.690 127.775 27.995 128.915 ;
        RECT 28.165 128.085 28.420 128.965 ;
        RECT 30.560 129.020 30.845 129.350 ;
        RECT 28.595 127.775 28.885 128.940 ;
        RECT 30.560 128.875 30.730 129.020 ;
        RECT 30.065 128.705 30.730 128.875 ;
        RECT 31.015 128.850 31.185 129.650 ;
        RECT 31.360 129.775 31.615 130.065 ;
        RECT 31.785 129.945 32.115 130.325 ;
        RECT 31.360 129.605 32.110 129.775 ;
        RECT 30.065 127.945 30.235 128.705 ;
        RECT 30.415 127.775 30.745 128.535 ;
        RECT 30.915 127.945 31.185 128.850 ;
        RECT 31.360 128.785 31.710 129.435 ;
        RECT 31.880 128.615 32.110 129.605 ;
        RECT 31.360 128.445 32.110 128.615 ;
        RECT 31.360 127.945 31.615 128.445 ;
        RECT 31.785 127.775 32.115 128.275 ;
        RECT 32.285 127.945 32.455 130.065 ;
        RECT 32.815 129.965 33.145 130.325 ;
        RECT 33.315 129.935 33.810 130.105 ;
        RECT 34.015 129.935 34.870 130.105 ;
        RECT 32.685 128.745 33.145 129.795 ;
        RECT 32.625 127.960 32.950 128.745 ;
        RECT 33.315 128.575 33.485 129.935 ;
        RECT 33.655 129.025 34.005 129.645 ;
        RECT 34.175 129.425 34.530 129.645 ;
        RECT 34.175 128.835 34.345 129.425 ;
        RECT 34.700 129.225 34.870 129.935 ;
        RECT 35.745 129.865 36.075 130.325 ;
        RECT 36.285 129.965 36.635 130.135 ;
        RECT 35.075 129.395 35.865 129.645 ;
        RECT 36.285 129.575 36.545 129.965 ;
        RECT 36.855 129.875 37.805 130.155 ;
        RECT 37.975 129.885 38.165 130.325 ;
        RECT 38.335 129.945 39.405 130.115 ;
        RECT 36.035 129.225 36.205 129.405 ;
        RECT 33.315 128.405 33.710 128.575 ;
        RECT 33.880 128.445 34.345 128.835 ;
        RECT 34.515 129.055 36.205 129.225 ;
        RECT 33.540 128.275 33.710 128.405 ;
        RECT 34.515 128.275 34.685 129.055 ;
        RECT 36.375 128.885 36.545 129.575 ;
        RECT 35.045 128.715 36.545 128.885 ;
        RECT 36.735 128.915 36.945 129.705 ;
        RECT 37.115 129.085 37.465 129.705 ;
        RECT 37.635 129.095 37.805 129.875 ;
        RECT 38.335 129.715 38.505 129.945 ;
        RECT 37.975 129.545 38.505 129.715 ;
        RECT 37.975 129.265 38.195 129.545 ;
        RECT 38.675 129.375 38.915 129.775 ;
        RECT 37.635 128.925 38.040 129.095 ;
        RECT 38.375 129.005 38.915 129.375 ;
        RECT 39.085 129.590 39.405 129.945 ;
        RECT 39.650 129.865 39.955 130.325 ;
        RECT 40.125 129.615 40.380 130.145 ;
        RECT 39.085 129.415 39.410 129.590 ;
        RECT 39.085 129.115 40.000 129.415 ;
        RECT 39.260 129.085 40.000 129.115 ;
        RECT 36.735 128.755 37.410 128.915 ;
        RECT 37.870 128.835 38.040 128.925 ;
        RECT 36.735 128.745 37.700 128.755 ;
        RECT 36.375 128.575 36.545 128.715 ;
        RECT 33.120 127.775 33.370 128.235 ;
        RECT 33.540 127.945 33.790 128.275 ;
        RECT 34.005 127.945 34.685 128.275 ;
        RECT 34.855 128.375 35.930 128.545 ;
        RECT 36.375 128.405 36.935 128.575 ;
        RECT 37.240 128.455 37.700 128.745 ;
        RECT 37.870 128.665 39.090 128.835 ;
        RECT 34.855 128.035 35.025 128.375 ;
        RECT 35.260 127.775 35.590 128.205 ;
        RECT 35.760 128.035 35.930 128.375 ;
        RECT 36.225 127.775 36.595 128.235 ;
        RECT 36.765 127.945 36.935 128.405 ;
        RECT 37.870 128.285 38.040 128.665 ;
        RECT 39.260 128.495 39.430 129.085 ;
        RECT 40.170 128.965 40.380 129.615 ;
        RECT 40.560 129.775 40.815 130.065 ;
        RECT 40.985 129.945 41.315 130.325 ;
        RECT 40.560 129.605 41.310 129.775 ;
        RECT 37.170 127.945 38.040 128.285 ;
        RECT 38.630 128.325 39.430 128.495 ;
        RECT 38.210 127.775 38.460 128.235 ;
        RECT 38.630 128.035 38.800 128.325 ;
        RECT 38.980 127.775 39.310 128.155 ;
        RECT 39.650 127.775 39.955 128.915 ;
        RECT 40.125 128.085 40.380 128.965 ;
        RECT 40.560 128.785 40.910 129.435 ;
        RECT 41.080 128.615 41.310 129.605 ;
        RECT 40.560 128.445 41.310 128.615 ;
        RECT 40.560 127.945 40.815 128.445 ;
        RECT 40.985 127.775 41.315 128.275 ;
        RECT 41.485 127.945 41.655 130.065 ;
        RECT 42.015 129.965 42.345 130.325 ;
        RECT 42.515 129.935 43.010 130.105 ;
        RECT 43.215 129.935 44.070 130.105 ;
        RECT 41.885 128.745 42.345 129.795 ;
        RECT 41.825 127.960 42.150 128.745 ;
        RECT 42.515 128.575 42.685 129.935 ;
        RECT 42.855 129.025 43.205 129.645 ;
        RECT 43.375 129.425 43.730 129.645 ;
        RECT 43.375 128.835 43.545 129.425 ;
        RECT 43.900 129.225 44.070 129.935 ;
        RECT 44.945 129.865 45.275 130.325 ;
        RECT 45.485 129.965 45.835 130.135 ;
        RECT 44.275 129.395 45.065 129.645 ;
        RECT 45.485 129.575 45.745 129.965 ;
        RECT 46.055 129.875 47.005 130.155 ;
        RECT 47.175 129.885 47.365 130.325 ;
        RECT 47.535 129.945 48.605 130.115 ;
        RECT 45.235 129.225 45.405 129.405 ;
        RECT 42.515 128.405 42.910 128.575 ;
        RECT 43.080 128.445 43.545 128.835 ;
        RECT 43.715 129.055 45.405 129.225 ;
        RECT 42.740 128.275 42.910 128.405 ;
        RECT 43.715 128.275 43.885 129.055 ;
        RECT 45.575 128.885 45.745 129.575 ;
        RECT 44.245 128.715 45.745 128.885 ;
        RECT 45.935 128.915 46.145 129.705 ;
        RECT 46.315 129.085 46.665 129.705 ;
        RECT 46.835 129.095 47.005 129.875 ;
        RECT 47.535 129.715 47.705 129.945 ;
        RECT 47.175 129.545 47.705 129.715 ;
        RECT 47.175 129.265 47.395 129.545 ;
        RECT 47.875 129.375 48.115 129.775 ;
        RECT 46.835 128.925 47.240 129.095 ;
        RECT 47.575 129.005 48.115 129.375 ;
        RECT 48.285 129.590 48.605 129.945 ;
        RECT 48.850 129.865 49.155 130.325 ;
        RECT 49.325 129.615 49.580 130.145 ;
        RECT 48.285 129.415 48.610 129.590 ;
        RECT 48.285 129.115 49.200 129.415 ;
        RECT 48.460 129.085 49.200 129.115 ;
        RECT 45.935 128.755 46.610 128.915 ;
        RECT 47.070 128.835 47.240 128.925 ;
        RECT 45.935 128.745 46.900 128.755 ;
        RECT 45.575 128.575 45.745 128.715 ;
        RECT 42.320 127.775 42.570 128.235 ;
        RECT 42.740 127.945 42.990 128.275 ;
        RECT 43.205 127.945 43.885 128.275 ;
        RECT 44.055 128.375 45.130 128.545 ;
        RECT 45.575 128.405 46.135 128.575 ;
        RECT 46.440 128.455 46.900 128.745 ;
        RECT 47.070 128.665 48.290 128.835 ;
        RECT 44.055 128.035 44.225 128.375 ;
        RECT 44.460 127.775 44.790 128.205 ;
        RECT 44.960 128.035 45.130 128.375 ;
        RECT 45.425 127.775 45.795 128.235 ;
        RECT 45.965 127.945 46.135 128.405 ;
        RECT 47.070 128.285 47.240 128.665 ;
        RECT 48.460 128.495 48.630 129.085 ;
        RECT 49.370 128.965 49.580 129.615 ;
        RECT 46.370 127.945 47.240 128.285 ;
        RECT 47.830 128.325 48.630 128.495 ;
        RECT 47.410 127.775 47.660 128.235 ;
        RECT 47.830 128.035 48.000 128.325 ;
        RECT 48.180 127.775 48.510 128.155 ;
        RECT 48.850 127.775 49.155 128.915 ;
        RECT 49.325 128.085 49.580 128.965 ;
        RECT 49.755 129.585 50.140 130.155 ;
        RECT 50.310 129.865 50.635 130.325 ;
        RECT 51.155 129.695 51.435 130.155 ;
        RECT 49.755 128.915 50.035 129.585 ;
        RECT 50.310 129.525 51.435 129.695 ;
        RECT 50.310 129.415 50.760 129.525 ;
        RECT 50.205 129.085 50.760 129.415 ;
        RECT 51.625 129.355 52.025 130.155 ;
        RECT 52.425 129.865 52.695 130.325 ;
        RECT 52.865 129.695 53.150 130.155 ;
        RECT 49.755 127.945 50.140 128.915 ;
        RECT 50.310 128.625 50.760 129.085 ;
        RECT 50.930 128.795 52.025 129.355 ;
        RECT 50.310 128.405 51.435 128.625 ;
        RECT 50.310 127.775 50.635 128.235 ;
        RECT 51.155 127.945 51.435 128.405 ;
        RECT 51.625 127.945 52.025 128.795 ;
        RECT 52.195 129.525 53.150 129.695 ;
        RECT 54.355 129.600 54.645 130.325 ;
        RECT 55.365 129.775 55.535 130.155 ;
        RECT 55.715 129.945 56.045 130.325 ;
        RECT 55.365 129.605 56.030 129.775 ;
        RECT 56.225 129.650 56.485 130.155 ;
        RECT 52.195 128.625 52.405 129.525 ;
        RECT 52.575 128.795 53.265 129.355 ;
        RECT 55.295 129.055 55.625 129.425 ;
        RECT 55.860 129.350 56.030 129.605 ;
        RECT 55.860 129.020 56.145 129.350 ;
        RECT 52.195 128.405 53.150 128.625 ;
        RECT 52.425 127.775 52.695 128.235 ;
        RECT 52.865 127.945 53.150 128.405 ;
        RECT 54.355 127.775 54.645 128.940 ;
        RECT 55.860 128.875 56.030 129.020 ;
        RECT 55.365 128.705 56.030 128.875 ;
        RECT 56.315 128.850 56.485 129.650 ;
        RECT 56.660 129.775 56.915 130.065 ;
        RECT 57.085 129.945 57.415 130.325 ;
        RECT 56.660 129.605 57.410 129.775 ;
        RECT 55.365 127.945 55.535 128.705 ;
        RECT 55.715 127.775 56.045 128.535 ;
        RECT 56.215 127.945 56.485 128.850 ;
        RECT 56.660 128.785 57.010 129.435 ;
        RECT 57.180 128.615 57.410 129.605 ;
        RECT 56.660 128.445 57.410 128.615 ;
        RECT 56.660 127.945 56.915 128.445 ;
        RECT 57.085 127.775 57.415 128.275 ;
        RECT 57.585 127.945 57.755 130.065 ;
        RECT 58.115 129.965 58.445 130.325 ;
        RECT 58.615 129.935 59.110 130.105 ;
        RECT 59.315 129.935 60.170 130.105 ;
        RECT 57.985 128.745 58.445 129.795 ;
        RECT 57.925 127.960 58.250 128.745 ;
        RECT 58.615 128.575 58.785 129.935 ;
        RECT 58.955 129.025 59.305 129.645 ;
        RECT 59.475 129.425 59.830 129.645 ;
        RECT 59.475 128.835 59.645 129.425 ;
        RECT 60.000 129.225 60.170 129.935 ;
        RECT 61.045 129.865 61.375 130.325 ;
        RECT 61.585 129.965 61.935 130.135 ;
        RECT 60.375 129.395 61.165 129.645 ;
        RECT 61.585 129.575 61.845 129.965 ;
        RECT 62.155 129.875 63.105 130.155 ;
        RECT 63.275 129.885 63.465 130.325 ;
        RECT 63.635 129.945 64.705 130.115 ;
        RECT 61.335 129.225 61.505 129.405 ;
        RECT 58.615 128.405 59.010 128.575 ;
        RECT 59.180 128.445 59.645 128.835 ;
        RECT 59.815 129.055 61.505 129.225 ;
        RECT 58.840 128.275 59.010 128.405 ;
        RECT 59.815 128.275 59.985 129.055 ;
        RECT 61.675 128.885 61.845 129.575 ;
        RECT 60.345 128.715 61.845 128.885 ;
        RECT 62.035 128.915 62.245 129.705 ;
        RECT 62.415 129.085 62.765 129.705 ;
        RECT 62.935 129.095 63.105 129.875 ;
        RECT 63.635 129.715 63.805 129.945 ;
        RECT 63.275 129.545 63.805 129.715 ;
        RECT 63.275 129.265 63.495 129.545 ;
        RECT 63.975 129.375 64.215 129.775 ;
        RECT 62.935 128.925 63.340 129.095 ;
        RECT 63.675 129.005 64.215 129.375 ;
        RECT 64.385 129.590 64.705 129.945 ;
        RECT 64.950 129.865 65.255 130.325 ;
        RECT 65.425 129.615 65.680 130.145 ;
        RECT 64.385 129.415 64.710 129.590 ;
        RECT 64.385 129.115 65.300 129.415 ;
        RECT 64.560 129.085 65.300 129.115 ;
        RECT 62.035 128.755 62.710 128.915 ;
        RECT 63.170 128.835 63.340 128.925 ;
        RECT 62.035 128.745 63.000 128.755 ;
        RECT 61.675 128.575 61.845 128.715 ;
        RECT 58.420 127.775 58.670 128.235 ;
        RECT 58.840 127.945 59.090 128.275 ;
        RECT 59.305 127.945 59.985 128.275 ;
        RECT 60.155 128.375 61.230 128.545 ;
        RECT 61.675 128.405 62.235 128.575 ;
        RECT 62.540 128.455 63.000 128.745 ;
        RECT 63.170 128.665 64.390 128.835 ;
        RECT 60.155 128.035 60.325 128.375 ;
        RECT 60.560 127.775 60.890 128.205 ;
        RECT 61.060 128.035 61.230 128.375 ;
        RECT 61.525 127.775 61.895 128.235 ;
        RECT 62.065 127.945 62.235 128.405 ;
        RECT 63.170 128.285 63.340 128.665 ;
        RECT 64.560 128.495 64.730 129.085 ;
        RECT 65.470 128.965 65.680 129.615 ;
        RECT 65.855 129.555 68.445 130.325 ;
        RECT 69.085 129.945 69.415 130.325 ;
        RECT 69.585 129.775 69.755 130.155 ;
        RECT 69.925 129.945 70.255 130.325 ;
        RECT 70.425 129.775 70.595 130.155 ;
        RECT 70.765 129.945 71.095 130.325 ;
        RECT 71.280 129.945 72.535 130.115 ;
        RECT 73.665 129.945 73.995 130.325 ;
        RECT 69.080 129.605 70.595 129.775 ;
        RECT 71.280 129.755 71.450 129.945 ;
        RECT 74.165 129.785 74.420 130.115 ;
        RECT 65.855 129.035 67.065 129.555 ;
        RECT 62.470 127.945 63.340 128.285 ;
        RECT 63.930 128.325 64.730 128.495 ;
        RECT 63.510 127.775 63.760 128.235 ;
        RECT 63.930 128.035 64.100 128.325 ;
        RECT 64.280 127.775 64.610 128.155 ;
        RECT 64.950 127.775 65.255 128.915 ;
        RECT 65.425 128.085 65.680 128.965 ;
        RECT 67.235 128.865 68.445 129.385 ;
        RECT 65.855 127.775 68.445 128.865 ;
        RECT 69.080 128.835 69.310 129.605 ;
        RECT 70.775 129.585 71.450 129.755 ;
        RECT 71.660 129.605 73.940 129.775 ;
        RECT 70.775 129.335 70.945 129.585 ;
        RECT 71.660 129.415 71.830 129.605 ;
        RECT 73.770 129.415 73.940 129.605 ;
        RECT 69.480 129.165 70.945 129.335 ;
        RECT 69.080 128.665 70.595 128.835 ;
        RECT 69.085 127.775 69.415 128.495 ;
        RECT 69.585 127.945 69.755 128.665 ;
        RECT 69.925 127.775 70.255 128.495 ;
        RECT 70.425 127.945 70.595 128.665 ;
        RECT 70.775 128.815 70.945 129.165 ;
        RECT 71.115 129.085 71.830 129.415 ;
        RECT 72.075 129.085 72.545 129.415 ;
        RECT 70.775 128.645 72.530 128.815 ;
        RECT 72.760 128.795 73.030 129.415 ;
        RECT 73.430 128.915 73.600 129.415 ;
        RECT 73.770 129.085 74.080 129.415 ;
        RECT 74.250 128.915 74.420 129.785 ;
        RECT 73.430 128.745 74.420 128.915 ;
        RECT 70.775 128.625 70.945 128.645 ;
        RECT 71.265 128.305 72.980 128.475 ;
        RECT 70.765 127.775 71.095 128.155 ;
        RECT 71.265 127.945 71.435 128.305 ;
        RECT 73.170 128.135 73.520 128.475 ;
        RECT 71.740 127.965 73.520 128.135 ;
        RECT 73.690 127.775 73.995 128.575 ;
        RECT 74.165 127.945 74.420 128.745 ;
        RECT 74.595 129.585 74.915 130.065 ;
        RECT 75.085 129.755 75.315 130.155 ;
        RECT 75.485 129.935 75.835 130.325 ;
        RECT 75.085 129.675 75.595 129.755 ;
        RECT 76.005 129.675 76.335 130.155 ;
        RECT 75.085 129.585 76.335 129.675 ;
        RECT 74.595 128.655 74.765 129.585 ;
        RECT 75.425 129.505 76.335 129.585 ;
        RECT 76.505 129.505 76.675 130.325 ;
        RECT 77.180 129.585 77.645 130.130 ;
        RECT 74.935 128.995 75.105 129.415 ;
        RECT 75.335 129.165 75.935 129.335 ;
        RECT 74.935 128.825 75.595 128.995 ;
        RECT 74.595 128.455 75.255 128.655 ;
        RECT 75.425 128.625 75.595 128.825 ;
        RECT 75.765 128.965 75.935 129.165 ;
        RECT 76.105 129.135 76.800 129.335 ;
        RECT 77.060 128.965 77.305 129.415 ;
        RECT 75.765 128.795 77.305 128.965 ;
        RECT 77.475 128.625 77.645 129.585 ;
        RECT 77.815 129.555 79.485 130.325 ;
        RECT 80.115 129.600 80.405 130.325 ;
        RECT 81.035 129.585 81.355 130.065 ;
        RECT 81.525 129.755 81.755 130.155 ;
        RECT 81.925 129.935 82.275 130.325 ;
        RECT 81.525 129.675 82.035 129.755 ;
        RECT 82.445 129.675 82.775 130.155 ;
        RECT 81.525 129.585 82.775 129.675 ;
        RECT 77.815 129.035 78.565 129.555 ;
        RECT 78.735 128.865 79.485 129.385 ;
        RECT 75.425 128.455 77.645 128.625 ;
        RECT 75.085 128.285 75.255 128.455 ;
        RECT 74.615 127.775 74.915 128.285 ;
        RECT 75.085 128.115 75.465 128.285 ;
        RECT 76.045 127.775 76.675 128.285 ;
        RECT 76.845 127.945 77.175 128.455 ;
        RECT 77.345 127.775 77.645 128.285 ;
        RECT 77.815 127.775 79.485 128.865 ;
        RECT 80.115 127.775 80.405 128.940 ;
        RECT 81.035 128.655 81.205 129.585 ;
        RECT 81.865 129.505 82.775 129.585 ;
        RECT 82.945 129.505 83.115 130.325 ;
        RECT 83.620 129.585 84.085 130.130 ;
        RECT 81.375 128.995 81.545 129.415 ;
        RECT 81.775 129.165 82.375 129.335 ;
        RECT 81.375 128.825 82.035 128.995 ;
        RECT 81.035 128.455 81.695 128.655 ;
        RECT 81.865 128.625 82.035 128.825 ;
        RECT 82.205 128.965 82.375 129.165 ;
        RECT 82.545 129.135 83.240 129.335 ;
        RECT 83.500 128.965 83.745 129.415 ;
        RECT 82.205 128.795 83.745 128.965 ;
        RECT 83.915 128.625 84.085 129.585 ;
        RECT 84.255 129.575 85.465 130.325 ;
        RECT 85.835 129.695 86.165 130.055 ;
        RECT 86.785 129.865 87.035 130.325 ;
        RECT 87.205 129.865 87.765 130.155 ;
        RECT 84.255 129.035 84.775 129.575 ;
        RECT 85.835 129.505 87.225 129.695 ;
        RECT 87.055 129.415 87.225 129.505 ;
        RECT 84.945 128.865 85.465 129.405 ;
        RECT 81.865 128.455 84.085 128.625 ;
        RECT 81.525 128.285 81.695 128.455 ;
        RECT 81.055 127.775 81.355 128.285 ;
        RECT 81.525 128.115 81.905 128.285 ;
        RECT 82.485 127.775 83.115 128.285 ;
        RECT 83.285 127.945 83.615 128.455 ;
        RECT 83.785 127.775 84.085 128.285 ;
        RECT 84.255 127.775 85.465 128.865 ;
        RECT 85.650 129.085 86.325 129.335 ;
        RECT 86.545 129.085 86.885 129.335 ;
        RECT 87.055 129.085 87.345 129.415 ;
        RECT 85.650 128.725 85.915 129.085 ;
        RECT 87.055 128.835 87.225 129.085 ;
        RECT 86.285 128.665 87.225 128.835 ;
        RECT 85.835 127.775 86.115 128.445 ;
        RECT 86.285 128.115 86.585 128.665 ;
        RECT 87.515 128.495 87.765 129.865 ;
        RECT 88.100 129.815 88.340 130.325 ;
        RECT 88.520 129.815 88.800 130.145 ;
        RECT 89.030 129.815 89.245 130.325 ;
        RECT 87.995 129.085 88.350 129.645 ;
        RECT 88.520 128.915 88.690 129.815 ;
        RECT 88.860 129.085 89.125 129.645 ;
        RECT 89.415 129.585 90.030 130.155 ;
        RECT 89.375 128.915 89.545 129.415 ;
        RECT 88.120 128.745 89.545 128.915 ;
        RECT 88.120 128.570 88.510 128.745 ;
        RECT 86.785 127.775 87.115 128.495 ;
        RECT 87.305 127.945 87.765 128.495 ;
        RECT 88.995 127.775 89.325 128.575 ;
        RECT 89.715 128.565 90.030 129.585 ;
        RECT 90.245 129.515 90.515 130.325 ;
        RECT 90.685 129.515 91.015 130.155 ;
        RECT 91.185 129.515 91.425 130.325 ;
        RECT 91.615 129.865 92.175 130.155 ;
        RECT 92.345 129.865 92.595 130.325 ;
        RECT 90.235 129.085 90.585 129.335 ;
        RECT 90.755 128.915 90.925 129.515 ;
        RECT 91.095 129.085 91.445 129.335 ;
        RECT 89.495 127.945 90.030 128.565 ;
        RECT 90.245 127.775 90.575 128.915 ;
        RECT 90.755 128.745 91.435 128.915 ;
        RECT 91.105 127.960 91.435 128.745 ;
        RECT 91.615 128.495 91.865 129.865 ;
        RECT 93.215 129.695 93.545 130.055 ;
        RECT 94.000 129.935 96.010 130.155 ;
        RECT 92.155 129.505 93.545 129.695 ;
        RECT 93.915 129.505 95.590 129.765 ;
        RECT 95.760 129.685 96.010 129.935 ;
        RECT 96.180 129.855 96.350 130.325 ;
        RECT 96.520 129.685 96.850 130.155 ;
        RECT 97.020 129.855 97.190 130.325 ;
        RECT 97.360 129.685 97.690 130.155 ;
        RECT 95.760 129.505 97.690 129.685 ;
        RECT 97.865 129.505 98.140 130.325 ;
        RECT 98.310 129.685 98.640 130.155 ;
        RECT 98.810 129.855 98.980 130.325 ;
        RECT 99.150 129.685 99.480 130.155 ;
        RECT 99.650 129.855 99.820 130.325 ;
        RECT 99.990 129.685 100.320 130.155 ;
        RECT 100.490 129.855 100.660 130.325 ;
        RECT 100.830 129.685 101.160 130.155 ;
        RECT 101.330 129.855 101.600 130.325 ;
        RECT 101.790 129.935 103.800 130.105 ;
        RECT 98.310 129.675 101.260 129.685 ;
        RECT 101.790 129.675 102.040 129.935 ;
        RECT 98.310 129.505 102.040 129.675 ;
        RECT 102.210 129.505 103.865 129.765 ;
        RECT 104.055 129.515 104.295 130.325 ;
        RECT 104.465 129.515 104.795 130.155 ;
        RECT 104.965 129.515 105.235 130.325 ;
        RECT 105.875 129.600 106.165 130.325 ;
        RECT 106.425 129.675 106.595 130.155 ;
        RECT 106.765 129.845 107.095 130.325 ;
        RECT 107.320 129.905 108.855 130.155 ;
        RECT 107.320 129.675 107.490 129.905 ;
        RECT 92.155 129.415 92.325 129.505 ;
        RECT 92.035 129.085 92.325 129.415 ;
        RECT 92.495 129.085 92.835 129.335 ;
        RECT 93.055 129.085 93.730 129.335 ;
        RECT 92.155 128.835 92.325 129.085 ;
        RECT 92.155 128.665 93.095 128.835 ;
        RECT 93.465 128.725 93.730 129.085 ;
        RECT 93.915 128.965 94.150 129.505 ;
        RECT 94.320 129.135 95.685 129.335 ;
        RECT 96.005 129.135 99.220 129.335 ;
        RECT 99.390 129.135 101.260 129.335 ;
        RECT 101.430 129.135 103.475 129.335 ;
        RECT 95.515 128.965 95.685 129.135 ;
        RECT 99.390 128.965 99.560 129.135 ;
        RECT 101.430 128.965 101.600 129.135 ;
        RECT 103.645 128.965 103.865 129.505 ;
        RECT 104.035 129.085 104.385 129.335 ;
        RECT 93.915 128.795 95.130 128.965 ;
        RECT 95.515 128.795 99.560 128.965 ;
        RECT 99.730 128.795 101.600 128.965 ;
        RECT 91.615 127.945 92.075 128.495 ;
        RECT 92.265 127.775 92.595 128.495 ;
        RECT 92.795 128.115 93.095 128.665 ;
        RECT 93.265 127.775 93.545 128.445 ;
        RECT 93.915 127.945 94.290 128.795 ;
        RECT 94.880 128.625 95.130 128.795 ;
        RECT 101.790 128.745 103.865 128.965 ;
        RECT 104.555 128.915 104.725 129.515 ;
        RECT 106.425 129.505 107.490 129.675 ;
        RECT 107.670 129.335 107.950 129.735 ;
        RECT 104.895 129.085 105.245 129.335 ;
        RECT 106.340 129.125 106.690 129.335 ;
        RECT 106.860 129.135 107.305 129.335 ;
        RECT 107.475 129.135 107.950 129.335 ;
        RECT 108.220 129.335 108.505 129.735 ;
        RECT 108.685 129.675 108.855 129.905 ;
        RECT 109.025 129.845 109.355 130.325 ;
        RECT 109.570 129.825 109.825 130.155 ;
        RECT 109.640 129.745 109.825 129.825 ;
        RECT 108.685 129.505 109.485 129.675 ;
        RECT 108.220 129.135 108.550 129.335 ;
        RECT 108.720 129.135 109.085 129.335 ;
        RECT 109.315 128.955 109.485 129.505 ;
        RECT 101.790 128.625 102.080 128.745 ;
        RECT 94.460 127.775 94.710 128.575 ;
        RECT 94.880 128.405 97.650 128.625 ;
        RECT 94.880 127.945 95.130 128.405 ;
        RECT 95.300 127.775 95.550 128.235 ;
        RECT 95.720 127.945 95.970 128.405 ;
        RECT 96.140 127.775 96.390 128.235 ;
        RECT 96.560 127.945 96.810 128.405 ;
        RECT 96.980 127.775 97.230 128.235 ;
        RECT 97.400 127.945 97.650 128.405 ;
        RECT 97.865 128.405 99.820 128.625 ;
        RECT 97.865 127.945 98.180 128.405 ;
        RECT 98.350 127.775 98.600 128.235 ;
        RECT 98.770 127.945 99.020 128.405 ;
        RECT 99.190 127.775 99.440 128.235 ;
        RECT 99.610 128.195 99.820 128.405 ;
        RECT 99.990 128.365 102.080 128.625 ;
        RECT 99.610 127.945 101.580 128.195 ;
        RECT 101.790 127.945 102.080 128.365 ;
        RECT 102.250 127.775 102.500 128.575 ;
        RECT 102.670 127.945 102.920 128.745 ;
        RECT 103.090 127.775 103.340 128.575 ;
        RECT 103.510 127.945 103.865 128.745 ;
        RECT 104.045 128.745 104.725 128.915 ;
        RECT 104.045 127.960 104.375 128.745 ;
        RECT 104.905 127.775 105.235 128.915 ;
        RECT 105.875 127.775 106.165 128.940 ;
        RECT 106.425 128.785 109.485 128.955 ;
        RECT 106.425 127.945 106.595 128.785 ;
        RECT 109.655 128.625 109.825 129.745 ;
        RECT 109.615 128.615 109.825 128.625 ;
        RECT 106.765 128.115 107.095 128.615 ;
        RECT 107.265 128.375 108.900 128.615 ;
        RECT 107.265 128.285 107.495 128.375 ;
        RECT 107.605 128.115 107.935 128.155 ;
        RECT 106.765 127.945 107.935 128.115 ;
        RECT 108.125 127.775 108.480 128.195 ;
        RECT 108.650 127.945 108.900 128.375 ;
        RECT 109.070 127.775 109.400 128.535 ;
        RECT 109.570 127.945 109.825 128.615 ;
        RECT 110.015 129.865 110.575 130.155 ;
        RECT 110.745 129.865 110.995 130.325 ;
        RECT 110.015 128.495 110.265 129.865 ;
        RECT 111.615 129.695 111.945 130.055 ;
        RECT 110.555 129.505 111.945 129.695 ;
        RECT 112.315 129.555 114.905 130.325 ;
        RECT 115.545 129.600 115.875 130.110 ;
        RECT 116.045 129.925 116.375 130.325 ;
        RECT 117.425 129.755 117.755 130.095 ;
        RECT 117.925 129.925 118.255 130.325 ;
        RECT 110.555 129.415 110.725 129.505 ;
        RECT 110.435 129.085 110.725 129.415 ;
        RECT 110.895 129.085 111.235 129.335 ;
        RECT 111.455 129.085 112.130 129.335 ;
        RECT 110.555 128.835 110.725 129.085 ;
        RECT 110.555 128.665 111.495 128.835 ;
        RECT 111.865 128.725 112.130 129.085 ;
        RECT 112.315 129.035 113.525 129.555 ;
        RECT 113.695 128.865 114.905 129.385 ;
        RECT 110.015 127.945 110.475 128.495 ;
        RECT 110.665 127.775 110.995 128.495 ;
        RECT 111.195 128.115 111.495 128.665 ;
        RECT 111.665 127.775 111.945 128.445 ;
        RECT 112.315 127.775 114.905 128.865 ;
        RECT 115.545 128.835 115.735 129.600 ;
        RECT 116.045 129.585 118.410 129.755 ;
        RECT 119.685 129.595 119.985 130.325 ;
        RECT 116.045 129.415 116.215 129.585 ;
        RECT 115.905 129.085 116.215 129.415 ;
        RECT 116.385 129.085 116.690 129.415 ;
        RECT 115.545 127.985 115.875 128.835 ;
        RECT 116.045 127.775 116.295 128.915 ;
        RECT 116.475 128.755 116.690 129.085 ;
        RECT 116.865 128.755 117.150 129.415 ;
        RECT 117.345 128.755 117.610 129.415 ;
        RECT 117.825 128.755 118.070 129.415 ;
        RECT 118.240 128.585 118.410 129.585 ;
        RECT 120.165 129.415 120.395 130.035 ;
        RECT 120.595 129.765 120.820 130.145 ;
        RECT 120.990 129.935 121.320 130.325 ;
        RECT 121.555 129.815 121.955 130.325 ;
        RECT 120.595 129.585 120.925 129.765 ;
        RECT 119.690 129.085 119.985 129.415 ;
        RECT 120.165 129.085 120.580 129.415 ;
        RECT 120.750 128.915 120.925 129.585 ;
        RECT 121.095 129.085 121.335 129.735 ;
        RECT 122.530 129.710 122.700 130.155 ;
        RECT 122.870 129.925 123.590 130.325 ;
        RECT 123.760 129.755 123.930 130.155 ;
        RECT 124.165 129.880 124.595 130.325 ;
        RECT 116.485 128.415 117.775 128.585 ;
        RECT 116.485 127.995 116.735 128.415 ;
        RECT 116.965 127.775 117.295 128.245 ;
        RECT 117.525 127.995 117.775 128.415 ;
        RECT 117.955 128.415 118.410 128.585 ;
        RECT 119.685 128.555 120.580 128.885 ;
        RECT 120.750 128.725 121.335 128.915 ;
        RECT 121.570 128.755 121.830 129.645 ;
        RECT 122.030 129.055 122.290 129.645 ;
        RECT 122.530 129.540 122.880 129.710 ;
        RECT 122.030 128.755 122.510 129.055 ;
        RECT 117.955 127.985 118.285 128.415 ;
        RECT 119.685 128.385 120.890 128.555 ;
        RECT 119.685 127.955 120.015 128.385 ;
        RECT 120.195 127.775 120.390 128.215 ;
        RECT 120.560 127.955 120.890 128.385 ;
        RECT 121.060 127.955 121.335 128.725 ;
        RECT 121.595 128.405 122.535 128.575 ;
        RECT 121.595 127.945 121.775 128.405 ;
        RECT 121.945 127.775 122.195 128.235 ;
        RECT 122.365 128.155 122.535 128.405 ;
        RECT 122.710 128.515 122.880 129.540 ;
        RECT 123.050 129.585 123.930 129.755 ;
        RECT 124.765 129.600 125.025 130.155 ;
        RECT 123.050 128.865 123.220 129.585 ;
        RECT 123.410 129.035 123.700 129.415 ;
        RECT 123.050 128.695 123.570 128.865 ;
        RECT 123.870 128.795 124.200 129.415 ;
        RECT 124.425 129.085 124.680 129.415 ;
        RECT 122.710 128.345 123.120 128.515 ;
        RECT 123.400 128.505 123.570 128.695 ;
        RECT 124.425 128.605 124.595 129.085 ;
        RECT 124.850 128.885 125.025 129.600 ;
        RECT 125.195 129.555 128.705 130.325 ;
        RECT 128.875 129.575 130.085 130.325 ;
        RECT 125.195 129.035 126.845 129.555 ;
        RECT 122.865 128.210 123.120 128.345 ;
        RECT 123.835 128.435 124.595 128.605 ;
        RECT 123.835 128.210 124.005 128.435 ;
        RECT 122.365 127.985 122.695 128.155 ;
        RECT 122.865 128.040 124.005 128.210 ;
        RECT 122.865 127.945 123.120 128.040 ;
        RECT 124.265 127.775 124.595 128.175 ;
        RECT 124.765 127.945 125.025 128.885 ;
        RECT 127.015 128.865 128.705 129.385 ;
        RECT 128.875 129.035 129.395 129.575 ;
        RECT 130.255 129.525 130.565 130.325 ;
        RECT 130.770 129.525 131.465 130.155 ;
        RECT 131.635 129.600 131.925 130.325 ;
        RECT 133.015 129.935 134.325 130.105 ;
        RECT 129.565 128.865 130.085 129.405 ;
        RECT 130.265 129.085 130.600 129.355 ;
        RECT 130.770 128.925 130.940 129.525 ;
        RECT 131.110 129.085 131.445 129.335 ;
        RECT 133.015 128.995 133.405 129.935 ;
        RECT 134.595 129.855 134.765 130.325 ;
        RECT 133.575 129.685 133.905 129.765 ;
        RECT 134.935 129.685 135.300 130.155 ;
        RECT 135.470 129.855 135.640 130.325 ;
        RECT 135.810 129.685 136.140 130.155 ;
        RECT 133.575 129.505 136.140 129.685 ;
        RECT 136.310 129.505 136.480 130.325 ;
        RECT 136.790 129.685 137.120 130.155 ;
        RECT 137.290 129.855 137.460 130.325 ;
        RECT 137.630 129.935 138.805 130.155 ;
        RECT 137.630 129.685 137.880 129.935 ;
        RECT 136.790 129.505 137.880 129.685 ;
        RECT 138.050 129.515 138.825 129.765 ;
        RECT 133.615 129.165 134.275 129.335 ;
        RECT 125.195 127.775 128.705 128.865 ;
        RECT 128.875 127.775 130.085 128.865 ;
        RECT 130.255 127.775 130.535 128.915 ;
        RECT 130.705 127.945 131.035 128.925 ;
        RECT 131.205 127.775 131.465 128.915 ;
        RECT 131.635 127.775 131.925 128.940 ;
        RECT 133.015 128.785 133.865 128.995 ;
        RECT 134.105 128.955 134.275 129.165 ;
        RECT 134.955 129.125 135.980 129.335 ;
        RECT 136.205 129.135 137.655 129.335 ;
        RECT 135.810 128.965 135.980 129.125 ;
        RECT 137.950 129.125 138.425 129.335 ;
        RECT 137.950 128.965 138.120 129.125 ;
        RECT 134.105 128.785 135.600 128.955 ;
        RECT 135.810 128.795 138.120 128.965 ;
        RECT 133.615 128.615 133.865 128.785 ;
        RECT 135.430 128.625 135.600 128.785 ;
        RECT 138.595 128.625 138.825 129.515 ;
        RECT 139.035 129.505 139.265 130.325 ;
        RECT 139.435 129.525 139.765 130.155 ;
        RECT 139.015 129.085 139.345 129.335 ;
        RECT 139.515 128.925 139.765 129.525 ;
        RECT 139.935 129.505 140.145 130.325 ;
        RECT 140.375 129.780 145.720 130.325 ;
        RECT 145.895 129.780 151.240 130.325 ;
        RECT 151.415 129.780 156.760 130.325 ;
        RECT 141.960 128.950 142.300 129.780 ;
        RECT 133.015 127.775 133.445 128.615 ;
        RECT 133.615 128.445 135.185 128.615 ;
        RECT 135.430 128.455 138.825 128.625 ;
        RECT 133.615 128.285 133.865 128.445 ;
        RECT 134.975 128.285 135.185 128.445 ;
        RECT 136.830 128.445 138.825 128.455 ;
        RECT 134.035 127.775 134.285 128.275 ;
        RECT 134.555 128.115 134.805 128.275 ;
        RECT 135.355 128.115 135.680 128.285 ;
        RECT 134.555 127.945 135.680 128.115 ;
        RECT 135.850 127.775 136.100 128.275 ;
        RECT 136.270 127.945 136.520 128.285 ;
        RECT 136.830 127.945 137.080 128.445 ;
        RECT 137.250 127.775 137.500 128.275 ;
        RECT 137.670 127.945 137.920 128.445 ;
        RECT 138.090 127.775 138.340 128.275 ;
        RECT 138.510 127.945 138.825 128.445 ;
        RECT 139.035 127.775 139.265 128.915 ;
        RECT 139.435 127.945 139.765 128.925 ;
        RECT 139.935 127.775 140.145 128.915 ;
        RECT 143.780 128.210 144.130 129.460 ;
        RECT 147.480 128.950 147.820 129.780 ;
        RECT 149.300 128.210 149.650 129.460 ;
        RECT 153.000 128.950 153.340 129.780 ;
        RECT 156.935 129.575 158.145 130.325 ;
        RECT 154.820 128.210 155.170 129.460 ;
        RECT 156.935 128.865 157.455 129.405 ;
        RECT 157.625 129.035 158.145 129.575 ;
        RECT 140.375 127.775 145.720 128.210 ;
        RECT 145.895 127.775 151.240 128.210 ;
        RECT 151.415 127.775 156.760 128.210 ;
        RECT 156.935 127.775 158.145 128.865 ;
        RECT 2.750 127.605 158.230 127.775 ;
        RECT 2.835 126.515 4.045 127.605 ;
        RECT 4.215 126.515 7.725 127.605 ;
        RECT 7.895 126.515 9.105 127.605 ;
        RECT 2.835 125.805 3.355 126.345 ;
        RECT 3.525 125.975 4.045 126.515 ;
        RECT 4.215 125.825 5.865 126.345 ;
        RECT 6.035 125.995 7.725 126.515 ;
        RECT 2.835 125.055 4.045 125.805 ;
        RECT 4.215 125.055 7.725 125.825 ;
        RECT 7.895 125.805 8.415 126.345 ;
        RECT 8.585 125.975 9.105 126.515 ;
        RECT 9.280 126.465 9.615 127.435 ;
        RECT 9.785 126.465 9.955 127.605 ;
        RECT 10.125 127.265 12.155 127.435 ;
        RECT 7.895 125.055 9.105 125.805 ;
        RECT 9.280 125.795 9.450 126.465 ;
        RECT 10.125 126.295 10.295 127.265 ;
        RECT 9.620 125.965 9.875 126.295 ;
        RECT 10.100 125.965 10.295 126.295 ;
        RECT 10.465 126.925 11.590 127.095 ;
        RECT 9.705 125.795 9.875 125.965 ;
        RECT 10.465 125.795 10.635 126.925 ;
        RECT 9.280 125.225 9.535 125.795 ;
        RECT 9.705 125.625 10.635 125.795 ;
        RECT 10.805 126.585 11.815 126.755 ;
        RECT 10.805 125.785 10.975 126.585 ;
        RECT 11.180 125.905 11.455 126.385 ;
        RECT 11.175 125.735 11.455 125.905 ;
        RECT 10.460 125.590 10.635 125.625 ;
        RECT 9.705 125.055 10.035 125.455 ;
        RECT 10.460 125.225 10.990 125.590 ;
        RECT 11.180 125.225 11.455 125.735 ;
        RECT 11.625 125.225 11.815 126.585 ;
        RECT 11.985 126.600 12.155 127.265 ;
        RECT 12.325 126.845 12.495 127.605 ;
        RECT 12.730 126.845 13.245 127.255 ;
        RECT 11.985 126.410 12.735 126.600 ;
        RECT 12.905 126.035 13.245 126.845 ;
        RECT 12.015 125.865 13.245 126.035 ;
        RECT 13.875 126.530 14.145 127.435 ;
        RECT 14.315 126.845 14.645 127.605 ;
        RECT 14.825 126.675 14.995 127.435 ;
        RECT 11.995 125.055 12.505 125.590 ;
        RECT 12.725 125.260 12.970 125.865 ;
        RECT 13.875 125.730 14.045 126.530 ;
        RECT 14.330 126.505 14.995 126.675 ;
        RECT 14.330 126.360 14.500 126.505 ;
        RECT 15.715 126.440 16.005 127.605 ;
        RECT 16.175 126.515 18.765 127.605 ;
        RECT 14.215 126.030 14.500 126.360 ;
        RECT 14.330 125.775 14.500 126.030 ;
        RECT 14.735 125.955 15.065 126.325 ;
        RECT 16.175 125.825 17.385 126.345 ;
        RECT 17.555 125.995 18.765 126.515 ;
        RECT 18.935 126.465 19.320 127.435 ;
        RECT 19.490 127.145 19.815 127.605 ;
        RECT 20.335 126.975 20.615 127.435 ;
        RECT 19.490 126.755 20.615 126.975 ;
        RECT 13.875 125.225 14.135 125.730 ;
        RECT 14.330 125.605 14.995 125.775 ;
        RECT 14.315 125.055 14.645 125.435 ;
        RECT 14.825 125.225 14.995 125.605 ;
        RECT 15.715 125.055 16.005 125.780 ;
        RECT 16.175 125.055 18.765 125.825 ;
        RECT 18.935 125.795 19.215 126.465 ;
        RECT 19.490 126.295 19.940 126.755 ;
        RECT 20.805 126.585 21.205 127.435 ;
        RECT 21.605 127.145 21.875 127.605 ;
        RECT 22.045 126.975 22.330 127.435 ;
        RECT 22.615 127.170 27.960 127.605 ;
        RECT 19.385 125.965 19.940 126.295 ;
        RECT 20.110 126.025 21.205 126.585 ;
        RECT 19.490 125.855 19.940 125.965 ;
        RECT 18.935 125.225 19.320 125.795 ;
        RECT 19.490 125.685 20.615 125.855 ;
        RECT 19.490 125.055 19.815 125.515 ;
        RECT 20.335 125.225 20.615 125.685 ;
        RECT 20.805 125.225 21.205 126.025 ;
        RECT 21.375 126.755 22.330 126.975 ;
        RECT 21.375 125.855 21.585 126.755 ;
        RECT 21.755 126.025 22.445 126.585 ;
        RECT 21.375 125.685 22.330 125.855 ;
        RECT 21.605 125.055 21.875 125.515 ;
        RECT 22.045 125.225 22.330 125.685 ;
        RECT 24.200 125.600 24.540 126.430 ;
        RECT 26.020 125.920 26.370 127.170 ;
        RECT 29.055 126.465 29.440 127.435 ;
        RECT 29.610 127.145 29.935 127.605 ;
        RECT 30.455 126.975 30.735 127.435 ;
        RECT 29.610 126.755 30.735 126.975 ;
        RECT 29.055 125.795 29.335 126.465 ;
        RECT 29.610 126.295 30.060 126.755 ;
        RECT 30.925 126.585 31.325 127.435 ;
        RECT 31.725 127.145 31.995 127.605 ;
        RECT 32.165 126.975 32.450 127.435 ;
        RECT 29.505 125.965 30.060 126.295 ;
        RECT 30.230 126.025 31.325 126.585 ;
        RECT 29.610 125.855 30.060 125.965 ;
        RECT 22.615 125.055 27.960 125.600 ;
        RECT 29.055 125.225 29.440 125.795 ;
        RECT 29.610 125.685 30.735 125.855 ;
        RECT 29.610 125.055 29.935 125.515 ;
        RECT 30.455 125.225 30.735 125.685 ;
        RECT 30.925 125.225 31.325 126.025 ;
        RECT 31.495 126.755 32.450 126.975 ;
        RECT 31.495 125.855 31.705 126.755 ;
        RECT 31.875 126.025 32.565 126.585 ;
        RECT 33.655 126.530 33.925 127.435 ;
        RECT 34.095 126.845 34.425 127.605 ;
        RECT 34.605 126.675 34.775 127.435 ;
        RECT 31.495 125.685 32.450 125.855 ;
        RECT 31.725 125.055 31.995 125.515 ;
        RECT 32.165 125.225 32.450 125.685 ;
        RECT 33.655 125.730 33.825 126.530 ;
        RECT 34.110 126.505 34.775 126.675 ;
        RECT 34.110 126.360 34.280 126.505 ;
        RECT 33.995 126.030 34.280 126.360 ;
        RECT 35.040 126.465 35.375 127.435 ;
        RECT 35.545 126.465 35.715 127.605 ;
        RECT 35.885 127.265 37.915 127.435 ;
        RECT 34.110 125.775 34.280 126.030 ;
        RECT 34.515 125.955 34.845 126.325 ;
        RECT 35.040 125.795 35.210 126.465 ;
        RECT 35.885 126.295 36.055 127.265 ;
        RECT 35.380 125.965 35.635 126.295 ;
        RECT 35.860 125.965 36.055 126.295 ;
        RECT 36.225 126.925 37.350 127.095 ;
        RECT 35.465 125.795 35.635 125.965 ;
        RECT 36.225 125.795 36.395 126.925 ;
        RECT 33.655 125.225 33.915 125.730 ;
        RECT 34.110 125.605 34.775 125.775 ;
        RECT 34.095 125.055 34.425 125.435 ;
        RECT 34.605 125.225 34.775 125.605 ;
        RECT 35.040 125.225 35.295 125.795 ;
        RECT 35.465 125.625 36.395 125.795 ;
        RECT 36.565 126.585 37.575 126.755 ;
        RECT 36.565 125.785 36.735 126.585 ;
        RECT 36.940 126.245 37.215 126.385 ;
        RECT 36.935 126.075 37.215 126.245 ;
        RECT 36.220 125.590 36.395 125.625 ;
        RECT 35.465 125.055 35.795 125.455 ;
        RECT 36.220 125.225 36.750 125.590 ;
        RECT 36.940 125.225 37.215 126.075 ;
        RECT 37.385 125.225 37.575 126.585 ;
        RECT 37.745 126.600 37.915 127.265 ;
        RECT 38.085 126.845 38.255 127.605 ;
        RECT 38.490 126.845 39.005 127.255 ;
        RECT 37.745 126.410 38.495 126.600 ;
        RECT 38.665 126.035 39.005 126.845 ;
        RECT 37.775 125.865 39.005 126.035 ;
        RECT 40.095 126.530 40.365 127.435 ;
        RECT 40.535 126.845 40.865 127.605 ;
        RECT 41.045 126.675 41.215 127.435 ;
        RECT 37.755 125.055 38.265 125.590 ;
        RECT 38.485 125.260 38.730 125.865 ;
        RECT 40.095 125.730 40.265 126.530 ;
        RECT 40.550 126.505 41.215 126.675 ;
        RECT 40.550 126.360 40.720 126.505 ;
        RECT 41.475 126.440 41.765 127.605 ;
        RECT 42.395 126.530 42.665 127.435 ;
        RECT 42.835 126.845 43.165 127.605 ;
        RECT 43.345 126.675 43.515 127.435 ;
        RECT 40.435 126.030 40.720 126.360 ;
        RECT 40.550 125.775 40.720 126.030 ;
        RECT 40.955 125.955 41.285 126.325 ;
        RECT 40.095 125.225 40.355 125.730 ;
        RECT 40.550 125.605 41.215 125.775 ;
        RECT 40.535 125.055 40.865 125.435 ;
        RECT 41.045 125.225 41.215 125.605 ;
        RECT 41.475 125.055 41.765 125.780 ;
        RECT 42.395 125.730 42.565 126.530 ;
        RECT 42.850 126.505 43.515 126.675 ;
        RECT 42.850 126.360 43.020 126.505 ;
        RECT 42.735 126.030 43.020 126.360 ;
        RECT 43.780 126.465 44.115 127.435 ;
        RECT 44.285 126.465 44.455 127.605 ;
        RECT 44.625 127.265 46.655 127.435 ;
        RECT 42.850 125.775 43.020 126.030 ;
        RECT 43.255 125.955 43.585 126.325 ;
        RECT 43.780 125.795 43.950 126.465 ;
        RECT 44.625 126.295 44.795 127.265 ;
        RECT 44.120 125.965 44.375 126.295 ;
        RECT 44.600 125.965 44.795 126.295 ;
        RECT 44.965 126.925 46.090 127.095 ;
        RECT 44.205 125.795 44.375 125.965 ;
        RECT 44.965 125.795 45.135 126.925 ;
        RECT 42.395 125.225 42.655 125.730 ;
        RECT 42.850 125.605 43.515 125.775 ;
        RECT 42.835 125.055 43.165 125.435 ;
        RECT 43.345 125.225 43.515 125.605 ;
        RECT 43.780 125.225 44.035 125.795 ;
        RECT 44.205 125.625 45.135 125.795 ;
        RECT 45.305 126.585 46.315 126.755 ;
        RECT 45.305 125.785 45.475 126.585 ;
        RECT 45.680 126.245 45.955 126.385 ;
        RECT 45.675 126.075 45.955 126.245 ;
        RECT 44.960 125.590 45.135 125.625 ;
        RECT 44.205 125.055 44.535 125.455 ;
        RECT 44.960 125.225 45.490 125.590 ;
        RECT 45.680 125.225 45.955 126.075 ;
        RECT 46.125 125.225 46.315 126.585 ;
        RECT 46.485 126.600 46.655 127.265 ;
        RECT 46.825 126.845 46.995 127.605 ;
        RECT 47.230 126.845 47.745 127.255 ;
        RECT 46.485 126.410 47.235 126.600 ;
        RECT 47.405 126.035 47.745 126.845 ;
        RECT 47.915 126.515 49.125 127.605 ;
        RECT 49.300 126.935 49.555 127.435 ;
        RECT 49.725 127.105 50.055 127.605 ;
        RECT 49.300 126.765 50.050 126.935 ;
        RECT 46.515 125.865 47.745 126.035 ;
        RECT 46.495 125.055 47.005 125.590 ;
        RECT 47.225 125.260 47.470 125.865 ;
        RECT 47.915 125.805 48.435 126.345 ;
        RECT 48.605 125.975 49.125 126.515 ;
        RECT 49.300 125.945 49.650 126.595 ;
        RECT 47.915 125.055 49.125 125.805 ;
        RECT 49.820 125.775 50.050 126.765 ;
        RECT 49.300 125.605 50.050 125.775 ;
        RECT 49.300 125.315 49.555 125.605 ;
        RECT 49.725 125.055 50.055 125.435 ;
        RECT 50.225 125.315 50.395 127.435 ;
        RECT 50.565 126.635 50.890 127.420 ;
        RECT 51.060 127.145 51.310 127.605 ;
        RECT 51.480 127.105 51.730 127.435 ;
        RECT 51.945 127.105 52.625 127.435 ;
        RECT 51.480 126.975 51.650 127.105 ;
        RECT 51.255 126.805 51.650 126.975 ;
        RECT 50.625 125.585 51.085 126.635 ;
        RECT 51.255 125.445 51.425 126.805 ;
        RECT 51.820 126.545 52.285 126.935 ;
        RECT 51.595 125.735 51.945 126.355 ;
        RECT 52.115 125.955 52.285 126.545 ;
        RECT 52.455 126.325 52.625 127.105 ;
        RECT 52.795 127.005 52.965 127.345 ;
        RECT 53.200 127.175 53.530 127.605 ;
        RECT 53.700 127.005 53.870 127.345 ;
        RECT 54.165 127.145 54.535 127.605 ;
        RECT 52.795 126.835 53.870 127.005 ;
        RECT 54.705 126.975 54.875 127.435 ;
        RECT 55.110 127.095 55.980 127.435 ;
        RECT 56.150 127.145 56.400 127.605 ;
        RECT 54.315 126.805 54.875 126.975 ;
        RECT 54.315 126.665 54.485 126.805 ;
        RECT 52.985 126.495 54.485 126.665 ;
        RECT 55.180 126.635 55.640 126.925 ;
        RECT 52.455 126.155 54.145 126.325 ;
        RECT 52.115 125.735 52.470 125.955 ;
        RECT 52.640 125.445 52.810 126.155 ;
        RECT 53.015 125.735 53.805 125.985 ;
        RECT 53.975 125.975 54.145 126.155 ;
        RECT 54.315 125.805 54.485 126.495 ;
        RECT 50.755 125.055 51.085 125.415 ;
        RECT 51.255 125.275 51.750 125.445 ;
        RECT 51.955 125.275 52.810 125.445 ;
        RECT 53.685 125.055 54.015 125.515 ;
        RECT 54.225 125.415 54.485 125.805 ;
        RECT 54.675 126.625 55.640 126.635 ;
        RECT 55.810 126.715 55.980 127.095 ;
        RECT 56.570 127.055 56.740 127.345 ;
        RECT 56.920 127.225 57.250 127.605 ;
        RECT 56.570 126.885 57.370 127.055 ;
        RECT 54.675 126.465 55.350 126.625 ;
        RECT 55.810 126.545 57.030 126.715 ;
        RECT 54.675 125.675 54.885 126.465 ;
        RECT 55.810 126.455 55.980 126.545 ;
        RECT 55.055 125.675 55.405 126.295 ;
        RECT 55.575 126.285 55.980 126.455 ;
        RECT 55.575 125.505 55.745 126.285 ;
        RECT 55.915 125.835 56.135 126.115 ;
        RECT 56.315 126.005 56.855 126.375 ;
        RECT 57.200 126.295 57.370 126.885 ;
        RECT 57.590 126.465 57.895 127.605 ;
        RECT 58.065 126.415 58.320 127.295 ;
        RECT 57.200 126.265 57.940 126.295 ;
        RECT 55.915 125.665 56.445 125.835 ;
        RECT 54.225 125.245 54.575 125.415 ;
        RECT 54.795 125.225 55.745 125.505 ;
        RECT 55.915 125.055 56.105 125.495 ;
        RECT 56.275 125.435 56.445 125.665 ;
        RECT 56.615 125.605 56.855 126.005 ;
        RECT 57.025 125.965 57.940 126.265 ;
        RECT 57.025 125.790 57.350 125.965 ;
        RECT 57.025 125.435 57.345 125.790 ;
        RECT 58.110 125.765 58.320 126.415 ;
        RECT 56.275 125.265 57.345 125.435 ;
        RECT 57.590 125.055 57.895 125.515 ;
        RECT 58.065 125.235 58.320 125.765 ;
        RECT 58.500 126.465 58.835 127.435 ;
        RECT 59.005 126.465 59.175 127.605 ;
        RECT 59.345 127.265 61.375 127.435 ;
        RECT 58.500 125.795 58.670 126.465 ;
        RECT 59.345 126.295 59.515 127.265 ;
        RECT 58.840 125.965 59.095 126.295 ;
        RECT 59.320 125.965 59.515 126.295 ;
        RECT 59.685 126.925 60.810 127.095 ;
        RECT 58.925 125.795 59.095 125.965 ;
        RECT 59.685 125.795 59.855 126.925 ;
        RECT 58.500 125.225 58.755 125.795 ;
        RECT 58.925 125.625 59.855 125.795 ;
        RECT 60.025 126.585 61.035 126.755 ;
        RECT 60.025 125.785 60.195 126.585 ;
        RECT 60.400 125.905 60.675 126.385 ;
        RECT 60.395 125.735 60.675 125.905 ;
        RECT 59.680 125.590 59.855 125.625 ;
        RECT 58.925 125.055 59.255 125.455 ;
        RECT 59.680 125.225 60.210 125.590 ;
        RECT 60.400 125.225 60.675 125.735 ;
        RECT 60.845 125.225 61.035 126.585 ;
        RECT 61.205 126.600 61.375 127.265 ;
        RECT 61.545 126.845 61.715 127.605 ;
        RECT 61.950 126.845 62.465 127.255 ;
        RECT 61.205 126.410 61.955 126.600 ;
        RECT 62.125 126.035 62.465 126.845 ;
        RECT 62.635 126.515 66.145 127.605 ;
        RECT 61.235 125.865 62.465 126.035 ;
        RECT 61.215 125.055 61.725 125.590 ;
        RECT 61.945 125.260 62.190 125.865 ;
        RECT 62.635 125.825 64.285 126.345 ;
        RECT 64.455 125.995 66.145 126.515 ;
        RECT 67.235 126.440 67.525 127.605 ;
        RECT 67.705 126.885 68.035 127.605 ;
        RECT 68.205 126.715 68.375 127.435 ;
        RECT 68.545 126.885 68.875 127.605 ;
        RECT 69.045 126.715 69.215 127.435 ;
        RECT 69.385 127.225 69.715 127.605 ;
        RECT 69.885 127.075 70.055 127.435 ;
        RECT 70.360 127.245 72.140 127.415 ;
        RECT 69.885 126.905 71.600 127.075 ;
        RECT 71.790 126.905 72.140 127.245 ;
        RECT 72.310 126.805 72.615 127.605 ;
        RECT 67.700 126.545 69.215 126.715 ;
        RECT 69.395 126.735 69.565 126.755 ;
        RECT 69.395 126.565 71.150 126.735 ;
        RECT 72.785 126.635 73.040 127.435 ;
        RECT 62.635 125.055 66.145 125.825 ;
        RECT 67.235 125.055 67.525 125.780 ;
        RECT 67.700 125.775 67.930 126.545 ;
        RECT 69.395 126.215 69.565 126.565 ;
        RECT 68.100 126.045 69.565 126.215 ;
        RECT 69.395 125.795 69.565 126.045 ;
        RECT 69.735 125.965 70.450 126.295 ;
        RECT 70.695 125.965 71.165 126.295 ;
        RECT 71.380 125.965 71.650 126.585 ;
        RECT 72.050 126.465 73.040 126.635 ;
        RECT 73.215 126.515 74.425 127.605 ;
        RECT 72.050 125.965 72.220 126.465 ;
        RECT 72.390 125.965 72.700 126.295 ;
        RECT 67.700 125.605 69.215 125.775 ;
        RECT 69.395 125.625 70.070 125.795 ;
        RECT 67.705 125.055 68.035 125.435 ;
        RECT 68.205 125.225 68.375 125.605 ;
        RECT 68.545 125.055 68.875 125.435 ;
        RECT 69.045 125.225 69.215 125.605 ;
        RECT 69.900 125.435 70.070 125.625 ;
        RECT 70.280 125.775 70.450 125.965 ;
        RECT 72.390 125.775 72.560 125.965 ;
        RECT 70.280 125.605 72.560 125.775 ;
        RECT 72.870 125.595 73.040 126.465 ;
        RECT 69.385 125.055 69.715 125.435 ;
        RECT 69.900 125.265 71.155 125.435 ;
        RECT 72.285 125.055 72.615 125.435 ;
        RECT 72.785 125.265 73.040 125.595 ;
        RECT 73.215 125.805 73.735 126.345 ;
        RECT 73.905 125.975 74.425 126.515 ;
        RECT 74.595 126.465 74.865 127.435 ;
        RECT 75.075 126.805 75.355 127.605 ;
        RECT 75.535 127.055 76.730 127.385 ;
        RECT 75.860 126.635 76.280 126.885 ;
        RECT 75.035 126.465 76.280 126.635 ;
        RECT 73.215 125.055 74.425 125.805 ;
        RECT 74.595 125.730 74.765 126.465 ;
        RECT 75.035 126.295 75.205 126.465 ;
        RECT 76.505 126.295 76.675 126.855 ;
        RECT 76.925 126.465 77.180 127.605 ;
        RECT 74.975 125.965 75.205 126.295 ;
        RECT 75.935 125.965 76.675 126.295 ;
        RECT 76.845 126.045 77.180 126.295 ;
        RECT 75.035 125.795 75.205 125.965 ;
        RECT 76.425 125.875 76.675 125.965 ;
        RECT 77.355 126.000 77.635 127.435 ;
        RECT 77.805 126.830 78.515 127.605 ;
        RECT 78.685 126.660 79.015 127.435 ;
        RECT 77.865 126.445 79.015 126.660 ;
        RECT 74.595 125.385 74.865 125.730 ;
        RECT 75.035 125.625 75.775 125.795 ;
        RECT 76.425 125.705 77.160 125.875 ;
        RECT 75.055 125.055 75.435 125.455 ;
        RECT 75.605 125.275 75.775 125.625 ;
        RECT 75.945 125.055 76.680 125.535 ;
        RECT 76.850 125.235 77.160 125.705 ;
        RECT 77.355 125.225 77.695 126.000 ;
        RECT 77.865 125.875 78.150 126.445 ;
        RECT 78.335 126.045 78.805 126.275 ;
        RECT 79.210 126.245 79.425 127.360 ;
        RECT 79.605 126.885 79.935 127.605 ;
        RECT 79.715 126.245 79.945 126.585 ;
        RECT 80.115 126.515 82.705 127.605 ;
        RECT 78.975 126.065 79.425 126.245 ;
        RECT 78.975 126.045 79.305 126.065 ;
        RECT 79.615 126.045 79.945 126.245 ;
        RECT 77.865 125.685 78.575 125.875 ;
        RECT 78.275 125.545 78.575 125.685 ;
        RECT 78.765 125.685 79.945 125.875 ;
        RECT 78.765 125.605 79.095 125.685 ;
        RECT 78.275 125.535 78.590 125.545 ;
        RECT 78.275 125.525 78.600 125.535 ;
        RECT 78.275 125.520 78.610 125.525 ;
        RECT 77.865 125.055 78.035 125.515 ;
        RECT 78.275 125.510 78.615 125.520 ;
        RECT 78.275 125.505 78.620 125.510 ;
        RECT 78.275 125.495 78.625 125.505 ;
        RECT 78.275 125.490 78.630 125.495 ;
        RECT 78.275 125.225 78.635 125.490 ;
        RECT 79.265 125.055 79.435 125.515 ;
        RECT 79.605 125.225 79.945 125.685 ;
        RECT 80.115 125.825 81.325 126.345 ;
        RECT 81.495 125.995 82.705 126.515 ;
        RECT 80.115 125.055 82.705 125.825 ;
        RECT 83.345 125.235 83.605 127.425 ;
        RECT 83.775 126.875 84.115 127.605 ;
        RECT 84.295 126.695 84.565 127.425 ;
        RECT 83.795 126.475 84.565 126.695 ;
        RECT 84.745 126.715 84.975 127.425 ;
        RECT 85.145 126.895 85.475 127.605 ;
        RECT 85.645 126.715 85.905 127.425 ;
        RECT 84.745 126.475 85.905 126.715 ;
        RECT 83.795 125.805 84.085 126.475 ;
        RECT 86.100 126.465 86.355 127.605 ;
        RECT 86.550 127.055 87.745 127.385 ;
        RECT 86.605 126.295 86.775 126.855 ;
        RECT 87.000 126.635 87.420 126.885 ;
        RECT 87.925 126.805 88.205 127.605 ;
        RECT 87.000 126.465 88.245 126.635 ;
        RECT 88.415 126.465 88.685 127.435 ;
        RECT 88.075 126.295 88.245 126.465 ;
        RECT 84.265 125.985 84.730 126.295 ;
        RECT 84.910 125.985 85.435 126.295 ;
        RECT 83.795 125.605 85.025 125.805 ;
        RECT 83.865 125.055 84.535 125.425 ;
        RECT 84.715 125.235 85.025 125.605 ;
        RECT 85.205 125.345 85.435 125.985 ;
        RECT 85.615 125.965 85.915 126.295 ;
        RECT 86.100 126.045 86.435 126.295 ;
        RECT 86.605 125.965 87.345 126.295 ;
        RECT 88.075 125.965 88.305 126.295 ;
        RECT 86.605 125.875 86.855 125.965 ;
        RECT 85.615 125.055 85.905 125.785 ;
        RECT 86.120 125.705 86.855 125.875 ;
        RECT 88.075 125.795 88.245 125.965 ;
        RECT 86.120 125.235 86.430 125.705 ;
        RECT 87.505 125.625 88.245 125.795 ;
        RECT 88.515 125.730 88.685 126.465 ;
        RECT 86.600 125.055 87.335 125.535 ;
        RECT 87.505 125.275 87.675 125.625 ;
        RECT 87.845 125.055 88.225 125.455 ;
        RECT 88.415 125.385 88.685 125.730 ;
        RECT 88.855 126.885 89.315 127.435 ;
        RECT 89.505 126.885 89.835 127.605 ;
        RECT 88.855 125.515 89.105 126.885 ;
        RECT 90.035 126.715 90.335 127.265 ;
        RECT 90.505 126.935 90.785 127.605 ;
        RECT 89.395 126.545 90.335 126.715 ;
        RECT 89.395 126.295 89.565 126.545 ;
        RECT 90.705 126.295 90.970 126.655 ;
        RECT 91.155 126.515 92.825 127.605 ;
        RECT 89.275 125.965 89.565 126.295 ;
        RECT 89.735 126.045 90.075 126.295 ;
        RECT 90.295 126.045 90.970 126.295 ;
        RECT 89.395 125.875 89.565 125.965 ;
        RECT 89.395 125.685 90.785 125.875 ;
        RECT 88.855 125.225 89.415 125.515 ;
        RECT 89.585 125.055 89.835 125.515 ;
        RECT 90.455 125.325 90.785 125.685 ;
        RECT 91.155 125.825 91.905 126.345 ;
        RECT 92.075 125.995 92.825 126.515 ;
        RECT 92.995 126.440 93.285 127.605 ;
        RECT 93.455 127.050 94.060 127.605 ;
        RECT 94.235 127.095 94.715 127.435 ;
        RECT 94.885 127.060 95.140 127.605 ;
        RECT 93.455 126.950 94.070 127.050 ;
        RECT 93.885 126.925 94.070 126.950 ;
        RECT 93.455 126.330 93.715 126.780 ;
        RECT 93.885 126.680 94.215 126.925 ;
        RECT 94.385 126.605 95.140 126.855 ;
        RECT 95.310 126.735 95.585 127.435 ;
        RECT 94.370 126.570 95.140 126.605 ;
        RECT 94.355 126.560 95.140 126.570 ;
        RECT 94.350 126.545 95.245 126.560 ;
        RECT 94.330 126.530 95.245 126.545 ;
        RECT 94.310 126.520 95.245 126.530 ;
        RECT 94.285 126.510 95.245 126.520 ;
        RECT 94.215 126.480 95.245 126.510 ;
        RECT 94.195 126.450 95.245 126.480 ;
        RECT 94.175 126.420 95.245 126.450 ;
        RECT 94.145 126.395 95.245 126.420 ;
        RECT 94.110 126.360 95.245 126.395 ;
        RECT 94.080 126.355 95.245 126.360 ;
        RECT 94.080 126.350 94.470 126.355 ;
        RECT 94.080 126.340 94.445 126.350 ;
        RECT 94.080 126.335 94.430 126.340 ;
        RECT 94.080 126.330 94.415 126.335 ;
        RECT 93.455 126.325 94.415 126.330 ;
        RECT 93.455 126.315 94.405 126.325 ;
        RECT 93.455 126.310 94.395 126.315 ;
        RECT 93.455 126.300 94.385 126.310 ;
        RECT 93.455 126.290 94.380 126.300 ;
        RECT 93.455 126.285 94.375 126.290 ;
        RECT 93.455 126.270 94.365 126.285 ;
        RECT 93.455 126.255 94.360 126.270 ;
        RECT 93.455 126.230 94.350 126.255 ;
        RECT 93.455 126.160 94.345 126.230 ;
        RECT 91.155 125.055 92.825 125.825 ;
        RECT 92.995 125.055 93.285 125.780 ;
        RECT 93.455 125.605 94.005 125.990 ;
        RECT 94.175 125.435 94.345 126.160 ;
        RECT 93.455 125.265 94.345 125.435 ;
        RECT 94.515 125.760 94.845 126.185 ;
        RECT 95.015 125.960 95.245 126.355 ;
        RECT 94.515 125.275 94.735 125.760 ;
        RECT 95.415 125.705 95.585 126.735 ;
        RECT 94.905 125.055 95.155 125.595 ;
        RECT 95.325 125.225 95.585 125.705 ;
        RECT 96.215 126.765 96.475 127.435 ;
        RECT 96.645 127.205 96.975 127.605 ;
        RECT 97.845 127.205 98.245 127.605 ;
        RECT 98.535 127.025 98.865 127.260 ;
        RECT 96.785 126.855 98.865 127.025 ;
        RECT 96.215 125.795 96.390 126.765 ;
        RECT 96.785 126.585 96.955 126.855 ;
        RECT 96.560 126.415 96.955 126.585 ;
        RECT 97.125 126.465 98.140 126.685 ;
        RECT 96.560 125.965 96.730 126.415 ;
        RECT 97.865 126.325 98.140 126.465 ;
        RECT 98.310 126.465 98.865 126.855 ;
        RECT 96.900 126.045 97.350 126.245 ;
        RECT 97.520 125.875 97.695 126.070 ;
        RECT 96.215 125.225 96.555 125.795 ;
        RECT 96.750 125.055 96.920 125.720 ;
        RECT 97.200 125.705 97.695 125.875 ;
        RECT 97.200 125.565 97.420 125.705 ;
        RECT 97.195 125.395 97.420 125.565 ;
        RECT 97.865 125.535 98.035 126.325 ;
        RECT 98.310 126.215 98.480 126.465 ;
        RECT 99.035 126.295 99.210 127.395 ;
        RECT 99.380 126.785 99.725 127.605 ;
        RECT 99.905 126.635 100.235 127.420 ;
        RECT 98.285 126.045 98.480 126.215 ;
        RECT 98.650 126.045 99.210 126.295 ;
        RECT 99.380 126.045 99.725 126.615 ;
        RECT 99.905 126.465 100.585 126.635 ;
        RECT 100.765 126.465 101.095 127.605 ;
        RECT 102.200 126.465 102.535 127.435 ;
        RECT 102.705 126.465 102.875 127.605 ;
        RECT 103.045 127.265 105.075 127.435 ;
        RECT 99.895 126.045 100.245 126.295 ;
        RECT 98.285 125.660 98.455 126.045 ;
        RECT 97.200 125.350 97.420 125.395 ;
        RECT 97.590 125.365 98.035 125.535 ;
        RECT 98.205 125.290 98.455 125.660 ;
        RECT 98.625 125.695 99.725 125.875 ;
        RECT 100.415 125.865 100.585 126.465 ;
        RECT 100.755 126.045 101.105 126.295 ;
        RECT 98.625 125.290 98.875 125.695 ;
        RECT 99.045 125.055 99.215 125.525 ;
        RECT 99.385 125.290 99.725 125.695 ;
        RECT 99.915 125.055 100.155 125.865 ;
        RECT 100.325 125.225 100.655 125.865 ;
        RECT 100.825 125.055 101.095 125.865 ;
        RECT 102.200 125.795 102.370 126.465 ;
        RECT 103.045 126.295 103.215 127.265 ;
        RECT 102.540 125.965 102.795 126.295 ;
        RECT 103.020 125.965 103.215 126.295 ;
        RECT 103.385 126.925 104.510 127.095 ;
        RECT 102.625 125.795 102.795 125.965 ;
        RECT 103.385 125.795 103.555 126.925 ;
        RECT 102.200 125.225 102.455 125.795 ;
        RECT 102.625 125.625 103.555 125.795 ;
        RECT 103.725 126.585 104.735 126.755 ;
        RECT 103.725 125.785 103.895 126.585 ;
        RECT 104.100 125.905 104.375 126.385 ;
        RECT 104.095 125.735 104.375 125.905 ;
        RECT 103.380 125.590 103.555 125.625 ;
        RECT 102.625 125.055 102.955 125.455 ;
        RECT 103.380 125.225 103.910 125.590 ;
        RECT 104.100 125.225 104.375 125.735 ;
        RECT 104.545 125.225 104.735 126.585 ;
        RECT 104.905 126.600 105.075 127.265 ;
        RECT 105.245 126.845 105.415 127.605 ;
        RECT 105.650 126.845 106.165 127.255 ;
        RECT 104.905 126.410 105.655 126.600 ;
        RECT 105.825 126.035 106.165 126.845 ;
        RECT 104.935 125.865 106.165 126.035 ;
        RECT 107.290 126.815 107.825 127.435 ;
        RECT 104.915 125.055 105.425 125.590 ;
        RECT 105.645 125.260 105.890 125.865 ;
        RECT 107.290 125.795 107.605 126.815 ;
        RECT 107.995 126.805 108.325 127.605 ;
        RECT 110.050 126.815 110.585 127.435 ;
        RECT 108.810 126.635 109.200 126.810 ;
        RECT 107.775 126.465 109.200 126.635 ;
        RECT 107.775 125.965 107.945 126.465 ;
        RECT 107.290 125.225 107.905 125.795 ;
        RECT 108.195 125.735 108.460 126.295 ;
        RECT 108.630 125.565 108.800 126.465 ;
        RECT 108.970 125.735 109.325 126.295 ;
        RECT 110.050 125.795 110.365 126.815 ;
        RECT 110.755 126.805 111.085 127.605 ;
        RECT 111.570 126.635 111.960 126.810 ;
        RECT 110.535 126.465 111.960 126.635 ;
        RECT 110.535 125.965 110.705 126.465 ;
        RECT 108.075 125.055 108.290 125.565 ;
        RECT 108.520 125.235 108.800 125.565 ;
        RECT 108.980 125.055 109.220 125.565 ;
        RECT 110.050 125.225 110.665 125.795 ;
        RECT 110.955 125.735 111.220 126.295 ;
        RECT 111.390 125.565 111.560 126.465 ;
        RECT 111.730 125.735 112.085 126.295 ;
        RECT 110.835 125.055 111.050 125.565 ;
        RECT 111.280 125.235 111.560 125.565 ;
        RECT 111.740 125.055 111.980 125.565 ;
        RECT 113.235 125.335 113.515 127.435 ;
        RECT 113.705 126.845 114.490 127.605 ;
        RECT 114.885 126.775 115.270 127.435 ;
        RECT 114.885 126.675 115.295 126.775 ;
        RECT 113.685 126.465 115.295 126.675 ;
        RECT 115.595 126.585 115.795 127.375 ;
        RECT 113.685 125.865 113.960 126.465 ;
        RECT 115.465 126.415 115.795 126.585 ;
        RECT 115.965 126.425 116.285 127.605 ;
        RECT 116.490 126.815 117.025 127.435 ;
        RECT 115.465 126.295 115.645 126.415 ;
        RECT 114.130 126.045 114.485 126.295 ;
        RECT 114.680 126.245 115.145 126.295 ;
        RECT 114.675 126.075 115.145 126.245 ;
        RECT 114.680 126.045 115.145 126.075 ;
        RECT 115.315 126.045 115.645 126.295 ;
        RECT 115.820 126.045 116.285 126.245 ;
        RECT 113.685 125.685 114.935 125.865 ;
        RECT 114.570 125.615 114.935 125.685 ;
        RECT 115.105 125.665 116.285 125.835 ;
        RECT 113.745 125.055 113.915 125.515 ;
        RECT 115.105 125.445 115.435 125.665 ;
        RECT 114.185 125.265 115.435 125.445 ;
        RECT 115.605 125.055 115.775 125.495 ;
        RECT 115.945 125.250 116.285 125.665 ;
        RECT 116.490 125.795 116.805 126.815 ;
        RECT 117.195 126.805 117.525 127.605 ;
        RECT 118.010 126.635 118.400 126.810 ;
        RECT 116.975 126.465 118.400 126.635 ;
        RECT 116.975 125.965 117.145 126.465 ;
        RECT 116.490 125.225 117.105 125.795 ;
        RECT 117.395 125.735 117.660 126.295 ;
        RECT 117.830 125.565 118.000 126.465 ;
        RECT 118.755 126.440 119.045 127.605 ;
        RECT 119.225 126.465 119.555 127.605 ;
        RECT 120.085 126.635 120.415 127.420 ;
        RECT 119.735 126.465 120.415 126.635 ;
        RECT 120.595 126.465 120.855 127.605 ;
        RECT 118.170 125.735 118.525 126.295 ;
        RECT 119.215 126.045 119.565 126.295 ;
        RECT 119.735 125.865 119.905 126.465 ;
        RECT 121.025 126.455 121.355 127.435 ;
        RECT 121.525 126.465 121.805 127.605 ;
        RECT 122.065 126.595 122.235 127.435 ;
        RECT 122.405 127.265 123.575 127.435 ;
        RECT 122.405 126.765 122.735 127.265 ;
        RECT 123.245 127.225 123.575 127.265 ;
        RECT 123.765 127.185 124.120 127.605 ;
        RECT 122.905 127.005 123.135 127.095 ;
        RECT 124.290 127.005 124.540 127.435 ;
        RECT 122.905 126.765 124.540 127.005 ;
        RECT 124.710 126.845 125.040 127.605 ;
        RECT 125.210 126.765 125.465 127.435 ;
        RECT 125.255 126.755 125.465 126.765 ;
        RECT 120.075 126.045 120.425 126.295 ;
        RECT 120.615 126.045 120.950 126.295 ;
        RECT 117.275 125.055 117.490 125.565 ;
        RECT 117.720 125.235 118.000 125.565 ;
        RECT 118.180 125.055 118.420 125.565 ;
        RECT 118.755 125.055 119.045 125.780 ;
        RECT 119.225 125.055 119.495 125.865 ;
        RECT 119.665 125.225 119.995 125.865 ;
        RECT 120.165 125.055 120.405 125.865 ;
        RECT 121.120 125.855 121.290 126.455 ;
        RECT 122.065 126.425 125.125 126.595 ;
        RECT 121.460 126.025 121.795 126.295 ;
        RECT 121.980 126.045 122.330 126.255 ;
        RECT 122.500 126.045 122.945 126.245 ;
        RECT 123.115 126.045 123.590 126.245 ;
        RECT 120.595 125.225 121.290 125.855 ;
        RECT 121.495 125.055 121.805 125.855 ;
        RECT 122.065 125.705 123.130 125.875 ;
        RECT 122.065 125.225 122.235 125.705 ;
        RECT 122.405 125.055 122.735 125.535 ;
        RECT 122.960 125.475 123.130 125.705 ;
        RECT 123.310 125.645 123.590 126.045 ;
        RECT 123.860 126.045 124.190 126.245 ;
        RECT 124.360 126.075 124.735 126.245 ;
        RECT 124.360 126.045 124.725 126.075 ;
        RECT 123.860 125.645 124.145 126.045 ;
        RECT 124.955 125.875 125.125 126.425 ;
        RECT 124.325 125.705 125.125 125.875 ;
        RECT 124.325 125.475 124.495 125.705 ;
        RECT 125.295 125.635 125.465 126.755 ;
        RECT 125.695 126.655 125.985 127.425 ;
        RECT 126.555 127.065 126.815 127.425 ;
        RECT 126.985 127.235 127.315 127.605 ;
        RECT 127.485 127.065 127.745 127.425 ;
        RECT 126.555 126.835 127.745 127.065 ;
        RECT 127.935 126.885 128.265 127.605 ;
        RECT 128.435 126.655 128.700 127.425 ;
        RECT 125.695 126.475 128.190 126.655 ;
        RECT 125.665 125.965 125.935 126.295 ;
        RECT 126.115 125.965 126.550 126.295 ;
        RECT 126.730 125.965 127.305 126.295 ;
        RECT 127.485 125.965 127.765 126.295 ;
        RECT 127.965 125.785 128.190 126.475 ;
        RECT 125.280 125.555 125.465 125.635 ;
        RECT 122.960 125.225 124.495 125.475 ;
        RECT 124.665 125.055 124.995 125.535 ;
        RECT 125.210 125.225 125.465 125.555 ;
        RECT 125.705 125.595 128.190 125.785 ;
        RECT 125.705 125.235 125.930 125.595 ;
        RECT 126.110 125.055 126.440 125.425 ;
        RECT 126.620 125.235 126.875 125.595 ;
        RECT 127.440 125.055 128.185 125.425 ;
        RECT 128.365 125.235 128.700 126.655 ;
        RECT 128.875 126.515 131.465 127.605 ;
        RECT 128.875 125.825 130.085 126.345 ;
        RECT 130.255 125.995 131.465 126.515 ;
        RECT 132.095 126.000 132.375 127.435 ;
        RECT 132.545 126.830 133.255 127.605 ;
        RECT 133.425 126.660 133.755 127.435 ;
        RECT 132.605 126.445 133.755 126.660 ;
        RECT 128.875 125.055 131.465 125.825 ;
        RECT 132.095 125.225 132.435 126.000 ;
        RECT 132.605 125.875 132.890 126.445 ;
        RECT 133.075 126.045 133.545 126.275 ;
        RECT 133.950 126.245 134.165 127.360 ;
        RECT 134.345 126.885 134.675 127.605 ;
        RECT 134.855 127.095 136.045 127.385 ;
        RECT 134.875 126.755 136.045 126.925 ;
        RECT 136.215 126.805 136.495 127.605 ;
        RECT 134.455 126.245 134.685 126.585 ;
        RECT 134.875 126.465 135.200 126.755 ;
        RECT 135.875 126.635 136.045 126.755 ;
        RECT 135.370 126.295 135.565 126.585 ;
        RECT 135.875 126.465 136.535 126.635 ;
        RECT 136.705 126.465 136.980 127.435 ;
        RECT 137.155 127.170 142.500 127.605 ;
        RECT 136.365 126.295 136.535 126.465 ;
        RECT 133.715 126.065 134.165 126.245 ;
        RECT 133.715 126.045 134.045 126.065 ;
        RECT 134.355 126.045 134.685 126.245 ;
        RECT 134.855 125.965 135.200 126.295 ;
        RECT 135.370 125.965 136.195 126.295 ;
        RECT 136.365 125.965 136.640 126.295 ;
        RECT 132.605 125.685 133.315 125.875 ;
        RECT 133.015 125.545 133.315 125.685 ;
        RECT 133.505 125.685 134.685 125.875 ;
        RECT 136.365 125.795 136.535 125.965 ;
        RECT 133.505 125.605 133.835 125.685 ;
        RECT 133.015 125.535 133.330 125.545 ;
        RECT 133.015 125.525 133.340 125.535 ;
        RECT 133.015 125.520 133.350 125.525 ;
        RECT 132.605 125.055 132.775 125.515 ;
        RECT 133.015 125.510 133.355 125.520 ;
        RECT 133.015 125.505 133.360 125.510 ;
        RECT 133.015 125.495 133.365 125.505 ;
        RECT 133.015 125.490 133.370 125.495 ;
        RECT 133.015 125.225 133.375 125.490 ;
        RECT 134.005 125.055 134.175 125.515 ;
        RECT 134.345 125.225 134.685 125.685 ;
        RECT 134.870 125.625 136.535 125.795 ;
        RECT 136.810 125.730 136.980 126.465 ;
        RECT 134.870 125.275 135.125 125.625 ;
        RECT 135.295 125.055 135.625 125.455 ;
        RECT 135.795 125.275 135.965 125.625 ;
        RECT 136.135 125.055 136.515 125.455 ;
        RECT 136.705 125.385 136.980 125.730 ;
        RECT 138.740 125.600 139.080 126.430 ;
        RECT 140.560 125.920 140.910 127.170 ;
        RECT 142.675 126.515 144.345 127.605 ;
        RECT 142.675 125.825 143.425 126.345 ;
        RECT 143.595 125.995 144.345 126.515 ;
        RECT 144.515 126.440 144.805 127.605 ;
        RECT 144.975 127.170 150.320 127.605 ;
        RECT 150.495 127.170 155.840 127.605 ;
        RECT 137.155 125.055 142.500 125.600 ;
        RECT 142.675 125.055 144.345 125.825 ;
        RECT 144.515 125.055 144.805 125.780 ;
        RECT 146.560 125.600 146.900 126.430 ;
        RECT 148.380 125.920 148.730 127.170 ;
        RECT 152.080 125.600 152.420 126.430 ;
        RECT 153.900 125.920 154.250 127.170 ;
        RECT 156.935 126.515 158.145 127.605 ;
        RECT 156.935 125.975 157.455 126.515 ;
        RECT 157.625 125.805 158.145 126.345 ;
        RECT 144.975 125.055 150.320 125.600 ;
        RECT 150.495 125.055 155.840 125.600 ;
        RECT 156.935 125.055 158.145 125.805 ;
        RECT 2.750 124.885 158.230 125.055 ;
        RECT 2.835 124.135 4.045 124.885 ;
        RECT 4.215 124.340 9.560 124.885 ;
        RECT 9.735 124.340 15.080 124.885 ;
        RECT 15.255 124.340 20.600 124.885 ;
        RECT 20.775 124.340 26.120 124.885 ;
        RECT 2.835 123.595 3.355 124.135 ;
        RECT 3.525 123.425 4.045 123.965 ;
        RECT 5.800 123.510 6.140 124.340 ;
        RECT 2.835 122.335 4.045 123.425 ;
        RECT 7.620 122.770 7.970 124.020 ;
        RECT 11.320 123.510 11.660 124.340 ;
        RECT 13.140 122.770 13.490 124.020 ;
        RECT 16.840 123.510 17.180 124.340 ;
        RECT 18.660 122.770 19.010 124.020 ;
        RECT 22.360 123.510 22.700 124.340 ;
        RECT 26.295 124.115 27.965 124.885 ;
        RECT 28.595 124.160 28.885 124.885 ;
        RECT 29.055 124.340 34.400 124.885 ;
        RECT 24.180 122.770 24.530 124.020 ;
        RECT 26.295 123.595 27.045 124.115 ;
        RECT 27.215 123.425 27.965 123.945 ;
        RECT 30.640 123.510 30.980 124.340 ;
        RECT 34.575 124.115 38.085 124.885 ;
        RECT 38.715 124.145 39.100 124.715 ;
        RECT 39.270 124.425 39.595 124.885 ;
        RECT 40.115 124.255 40.395 124.715 ;
        RECT 4.215 122.335 9.560 122.770 ;
        RECT 9.735 122.335 15.080 122.770 ;
        RECT 15.255 122.335 20.600 122.770 ;
        RECT 20.775 122.335 26.120 122.770 ;
        RECT 26.295 122.335 27.965 123.425 ;
        RECT 28.595 122.335 28.885 123.500 ;
        RECT 32.460 122.770 32.810 124.020 ;
        RECT 34.575 123.595 36.225 124.115 ;
        RECT 36.395 123.425 38.085 123.945 ;
        RECT 29.055 122.335 34.400 122.770 ;
        RECT 34.575 122.335 38.085 123.425 ;
        RECT 38.715 123.475 38.995 124.145 ;
        RECT 39.270 124.085 40.395 124.255 ;
        RECT 39.270 123.975 39.720 124.085 ;
        RECT 39.165 123.645 39.720 123.975 ;
        RECT 40.585 123.915 40.985 124.715 ;
        RECT 41.385 124.425 41.655 124.885 ;
        RECT 41.825 124.255 42.110 124.715 ;
        RECT 42.395 124.340 47.740 124.885 ;
        RECT 38.715 122.505 39.100 123.475 ;
        RECT 39.270 123.185 39.720 123.645 ;
        RECT 39.890 123.355 40.985 123.915 ;
        RECT 39.270 122.965 40.395 123.185 ;
        RECT 39.270 122.335 39.595 122.795 ;
        RECT 40.115 122.505 40.395 122.965 ;
        RECT 40.585 122.505 40.985 123.355 ;
        RECT 41.155 124.085 42.110 124.255 ;
        RECT 41.155 123.185 41.365 124.085 ;
        RECT 41.535 123.355 42.225 123.915 ;
        RECT 43.980 123.510 44.320 124.340 ;
        RECT 47.915 124.145 48.300 124.715 ;
        RECT 48.470 124.425 48.795 124.885 ;
        RECT 49.315 124.255 49.595 124.715 ;
        RECT 41.155 122.965 42.110 123.185 ;
        RECT 41.385 122.335 41.655 122.795 ;
        RECT 41.825 122.505 42.110 122.965 ;
        RECT 45.800 122.770 46.150 124.020 ;
        RECT 47.915 123.475 48.195 124.145 ;
        RECT 48.470 124.085 49.595 124.255 ;
        RECT 48.470 123.975 48.920 124.085 ;
        RECT 48.365 123.645 48.920 123.975 ;
        RECT 49.785 123.915 50.185 124.715 ;
        RECT 50.585 124.425 50.855 124.885 ;
        RECT 51.025 124.255 51.310 124.715 ;
        RECT 42.395 122.335 47.740 122.770 ;
        RECT 47.915 122.505 48.300 123.475 ;
        RECT 48.470 123.185 48.920 123.645 ;
        RECT 49.090 123.355 50.185 123.915 ;
        RECT 48.470 122.965 49.595 123.185 ;
        RECT 48.470 122.335 48.795 122.795 ;
        RECT 49.315 122.505 49.595 122.965 ;
        RECT 49.785 122.505 50.185 123.355 ;
        RECT 50.355 124.085 51.310 124.255 ;
        RECT 51.595 124.115 54.185 124.885 ;
        RECT 54.355 124.160 54.645 124.885 ;
        RECT 54.815 124.340 60.160 124.885 ;
        RECT 60.335 124.340 65.680 124.885 ;
        RECT 50.355 123.185 50.565 124.085 ;
        RECT 50.735 123.355 51.425 123.915 ;
        RECT 51.595 123.595 52.805 124.115 ;
        RECT 52.975 123.425 54.185 123.945 ;
        RECT 56.400 123.510 56.740 124.340 ;
        RECT 50.355 122.965 51.310 123.185 ;
        RECT 50.585 122.335 50.855 122.795 ;
        RECT 51.025 122.505 51.310 122.965 ;
        RECT 51.595 122.335 54.185 123.425 ;
        RECT 54.355 122.335 54.645 123.500 ;
        RECT 58.220 122.770 58.570 124.020 ;
        RECT 61.920 123.510 62.260 124.340 ;
        RECT 65.855 124.115 67.525 124.885 ;
        RECT 67.705 124.505 68.035 124.885 ;
        RECT 68.205 124.335 68.375 124.715 ;
        RECT 68.545 124.505 68.875 124.885 ;
        RECT 69.045 124.335 69.215 124.715 ;
        RECT 69.385 124.505 69.715 124.885 ;
        RECT 69.900 124.505 71.155 124.675 ;
        RECT 72.285 124.505 72.615 124.885 ;
        RECT 67.700 124.165 69.215 124.335 ;
        RECT 69.900 124.315 70.070 124.505 ;
        RECT 72.785 124.345 73.040 124.675 ;
        RECT 63.740 122.770 64.090 124.020 ;
        RECT 65.855 123.595 66.605 124.115 ;
        RECT 66.775 123.425 67.525 123.945 ;
        RECT 54.815 122.335 60.160 122.770 ;
        RECT 60.335 122.335 65.680 122.770 ;
        RECT 65.855 122.335 67.525 123.425 ;
        RECT 67.700 123.395 67.930 124.165 ;
        RECT 69.395 124.145 70.070 124.315 ;
        RECT 70.280 124.165 72.560 124.335 ;
        RECT 69.395 123.895 69.565 124.145 ;
        RECT 70.280 123.975 70.450 124.165 ;
        RECT 72.390 123.975 72.560 124.165 ;
        RECT 68.100 123.725 69.565 123.895 ;
        RECT 67.700 123.225 69.215 123.395 ;
        RECT 67.705 122.335 68.035 123.055 ;
        RECT 68.205 122.505 68.375 123.225 ;
        RECT 68.545 122.335 68.875 123.055 ;
        RECT 69.045 122.505 69.215 123.225 ;
        RECT 69.395 123.375 69.565 123.725 ;
        RECT 69.735 123.645 70.450 123.975 ;
        RECT 70.695 123.645 71.165 123.975 ;
        RECT 69.395 123.205 71.150 123.375 ;
        RECT 71.380 123.355 71.650 123.975 ;
        RECT 72.050 123.475 72.220 123.975 ;
        RECT 72.390 123.645 72.700 123.975 ;
        RECT 72.870 123.475 73.040 124.345 ;
        RECT 73.215 124.115 74.885 124.885 ;
        RECT 75.385 124.485 75.715 124.885 ;
        RECT 75.885 124.315 76.215 124.655 ;
        RECT 77.265 124.485 77.595 124.885 ;
        RECT 75.230 124.145 77.595 124.315 ;
        RECT 77.765 124.160 78.095 124.670 ;
        RECT 73.215 123.595 73.965 124.115 ;
        RECT 72.050 123.305 73.040 123.475 ;
        RECT 74.135 123.425 74.885 123.945 ;
        RECT 69.395 123.185 69.565 123.205 ;
        RECT 69.885 122.865 71.600 123.035 ;
        RECT 69.385 122.335 69.715 122.715 ;
        RECT 69.885 122.505 70.055 122.865 ;
        RECT 71.790 122.695 72.140 123.035 ;
        RECT 70.360 122.525 72.140 122.695 ;
        RECT 72.310 122.335 72.615 123.135 ;
        RECT 72.785 122.505 73.040 123.305 ;
        RECT 73.215 122.335 74.885 123.425 ;
        RECT 75.230 123.145 75.400 124.145 ;
        RECT 77.425 123.975 77.595 124.145 ;
        RECT 75.570 123.315 75.815 123.975 ;
        RECT 76.030 123.315 76.295 123.975 ;
        RECT 76.490 123.315 76.775 123.975 ;
        RECT 76.950 123.645 77.255 123.975 ;
        RECT 77.425 123.645 77.735 123.975 ;
        RECT 76.950 123.315 77.165 123.645 ;
        RECT 75.230 122.975 75.685 123.145 ;
        RECT 75.355 122.545 75.685 122.975 ;
        RECT 75.865 122.975 77.155 123.145 ;
        RECT 75.865 122.555 76.115 122.975 ;
        RECT 76.345 122.335 76.675 122.805 ;
        RECT 76.905 122.555 77.155 122.975 ;
        RECT 77.345 122.335 77.595 123.475 ;
        RECT 77.905 123.395 78.095 124.160 ;
        RECT 78.275 124.085 78.970 124.715 ;
        RECT 79.175 124.085 79.485 124.885 ;
        RECT 80.115 124.160 80.405 124.885 ;
        RECT 80.575 124.495 81.885 124.665 ;
        RECT 78.795 124.035 78.970 124.085 ;
        RECT 78.295 123.645 78.630 123.895 ;
        RECT 78.800 123.485 78.970 124.035 ;
        RECT 79.140 123.645 79.475 123.915 ;
        RECT 80.575 123.555 80.965 124.495 ;
        RECT 82.155 124.415 82.325 124.885 ;
        RECT 81.135 124.245 81.465 124.325 ;
        RECT 82.495 124.245 82.860 124.715 ;
        RECT 83.030 124.415 83.200 124.885 ;
        RECT 83.370 124.245 83.700 124.715 ;
        RECT 81.135 124.065 83.700 124.245 ;
        RECT 83.870 124.065 84.040 124.885 ;
        RECT 84.350 124.245 84.680 124.715 ;
        RECT 84.850 124.415 85.020 124.885 ;
        RECT 85.190 124.495 86.365 124.715 ;
        RECT 85.190 124.245 85.440 124.495 ;
        RECT 84.350 124.065 85.440 124.245 ;
        RECT 85.610 124.075 86.385 124.325 ;
        RECT 86.565 124.315 86.895 124.675 ;
        RECT 87.065 124.505 87.395 124.885 ;
        RECT 87.645 124.315 87.815 124.715 ;
        RECT 87.995 124.505 89.715 124.675 ;
        RECT 90.225 124.505 90.555 124.885 ;
        RECT 86.565 124.145 88.775 124.315 ;
        RECT 88.965 124.145 90.975 124.315 ;
        RECT 91.155 124.165 91.495 124.675 ;
        RECT 81.175 123.725 81.835 123.895 ;
        RECT 77.765 122.545 78.095 123.395 ;
        RECT 78.275 122.335 78.535 123.475 ;
        RECT 78.705 122.505 79.035 123.485 ;
        RECT 79.205 122.335 79.485 123.475 ;
        RECT 80.115 122.335 80.405 123.500 ;
        RECT 80.575 123.345 81.425 123.555 ;
        RECT 81.665 123.515 81.835 123.725 ;
        RECT 82.515 123.865 83.540 123.895 ;
        RECT 82.515 123.695 83.565 123.865 ;
        RECT 83.765 123.695 85.215 123.895 ;
        RECT 82.515 123.685 83.540 123.695 ;
        RECT 83.370 123.525 83.540 123.685 ;
        RECT 85.510 123.685 85.985 123.895 ;
        RECT 85.510 123.525 85.680 123.685 ;
        RECT 81.665 123.345 83.160 123.515 ;
        RECT 83.370 123.355 85.680 123.525 ;
        RECT 81.175 123.175 81.425 123.345 ;
        RECT 82.990 123.185 83.160 123.345 ;
        RECT 86.155 123.185 86.385 124.075 ;
        RECT 86.580 123.695 87.250 123.895 ;
        RECT 86.580 123.345 86.805 123.695 ;
        RECT 87.500 123.525 87.815 124.145 ;
        RECT 87.995 123.645 88.165 123.975 ;
        RECT 86.985 123.355 87.815 123.525 ;
        RECT 88.405 123.355 89.115 123.975 ;
        RECT 89.315 123.355 90.020 123.975 ;
        RECT 90.250 123.355 90.925 123.975 ;
        RECT 80.575 122.335 81.005 123.175 ;
        RECT 81.175 123.005 82.745 123.175 ;
        RECT 82.990 123.015 86.385 123.185 ;
        RECT 81.175 122.845 81.425 123.005 ;
        RECT 82.535 122.845 82.745 123.005 ;
        RECT 84.390 123.005 86.385 123.015 ;
        RECT 81.595 122.335 81.845 122.835 ;
        RECT 82.115 122.675 82.365 122.835 ;
        RECT 82.915 122.675 83.240 122.845 ;
        RECT 82.115 122.505 83.240 122.675 ;
        RECT 83.410 122.335 83.660 122.835 ;
        RECT 83.830 122.505 84.080 122.845 ;
        RECT 84.390 122.505 84.640 123.005 ;
        RECT 84.810 122.335 85.060 122.835 ;
        RECT 85.230 122.505 85.480 123.005 ;
        RECT 85.650 122.335 85.900 122.835 ;
        RECT 86.070 122.505 86.385 123.005 ;
        RECT 86.645 122.675 86.815 123.175 ;
        RECT 86.985 122.855 87.315 123.355 ;
        RECT 87.565 123.015 90.895 123.185 ;
        RECT 87.565 122.675 87.735 123.015 ;
        RECT 86.645 122.505 87.735 122.675 ;
        RECT 88.090 122.335 88.760 122.845 ;
        RECT 89.045 122.505 89.215 123.015 ;
        RECT 89.385 122.335 89.715 122.845 ;
        RECT 89.885 122.505 90.055 123.015 ;
        RECT 90.225 122.335 90.555 122.845 ;
        RECT 90.725 122.505 90.895 123.015 ;
        RECT 91.155 122.765 91.415 124.165 ;
        RECT 91.665 124.085 91.935 124.885 ;
        RECT 91.590 123.645 91.920 123.895 ;
        RECT 92.115 123.645 92.395 124.615 ;
        RECT 92.575 123.645 92.875 124.615 ;
        RECT 93.055 123.645 93.405 124.610 ;
        RECT 93.625 124.385 94.120 124.715 ;
        RECT 91.605 123.475 91.920 123.645 ;
        RECT 93.625 123.475 93.795 124.385 ;
        RECT 91.605 123.305 93.795 123.475 ;
        RECT 91.155 122.505 91.495 122.765 ;
        RECT 91.665 122.335 91.995 123.135 ;
        RECT 92.460 122.505 92.710 123.305 ;
        RECT 92.895 122.335 93.225 123.055 ;
        RECT 93.445 122.505 93.695 123.305 ;
        RECT 93.965 122.895 94.205 124.205 ;
        RECT 94.380 123.285 94.715 124.705 ;
        RECT 94.895 124.515 95.640 124.885 ;
        RECT 96.205 124.345 96.460 124.705 ;
        RECT 96.640 124.515 96.970 124.885 ;
        RECT 97.150 124.345 97.375 124.705 ;
        RECT 94.890 124.155 97.375 124.345 ;
        RECT 94.890 123.465 95.115 124.155 ;
        RECT 98.115 124.065 98.325 124.885 ;
        RECT 98.495 124.085 98.825 124.715 ;
        RECT 95.315 123.645 95.595 123.975 ;
        RECT 95.775 123.645 96.350 123.975 ;
        RECT 96.530 123.645 96.965 123.975 ;
        RECT 97.145 123.645 97.415 123.975 ;
        RECT 98.495 123.485 98.745 124.085 ;
        RECT 98.995 124.065 99.225 124.885 ;
        RECT 99.435 124.115 102.945 124.885 ;
        RECT 98.915 123.645 99.245 123.895 ;
        RECT 99.435 123.595 101.085 124.115 ;
        RECT 94.890 123.285 97.385 123.465 ;
        RECT 93.865 122.335 94.200 122.715 ;
        RECT 94.380 122.515 94.645 123.285 ;
        RECT 94.815 122.335 95.145 123.055 ;
        RECT 95.335 122.875 96.525 123.105 ;
        RECT 95.335 122.515 95.595 122.875 ;
        RECT 95.765 122.335 96.095 122.705 ;
        RECT 96.265 122.515 96.525 122.875 ;
        RECT 97.095 122.515 97.385 123.285 ;
        RECT 98.115 122.335 98.325 123.475 ;
        RECT 98.495 122.505 98.825 123.485 ;
        RECT 98.995 122.335 99.225 123.475 ;
        RECT 101.255 123.425 102.945 123.945 ;
        RECT 99.435 122.335 102.945 123.425 ;
        RECT 103.125 122.515 103.385 124.705 ;
        RECT 103.645 124.515 104.315 124.885 ;
        RECT 104.495 124.335 104.805 124.705 ;
        RECT 103.575 124.135 104.805 124.335 ;
        RECT 103.575 123.465 103.865 124.135 ;
        RECT 104.985 123.955 105.215 124.595 ;
        RECT 105.395 124.155 105.685 124.885 ;
        RECT 105.875 124.160 106.165 124.885 ;
        RECT 106.345 124.155 106.645 124.885 ;
        RECT 106.825 123.975 107.055 124.595 ;
        RECT 107.255 124.325 107.480 124.705 ;
        RECT 107.650 124.495 107.980 124.885 ;
        RECT 107.255 124.145 107.585 124.325 ;
        RECT 104.045 123.645 104.510 123.955 ;
        RECT 104.690 123.645 105.215 123.955 ;
        RECT 105.395 123.645 105.695 123.975 ;
        RECT 106.350 123.645 106.645 123.975 ;
        RECT 106.825 123.645 107.240 123.975 ;
        RECT 103.575 123.245 104.345 123.465 ;
        RECT 103.555 122.335 103.895 123.065 ;
        RECT 104.075 122.515 104.345 123.245 ;
        RECT 104.525 123.225 105.685 123.465 ;
        RECT 104.525 122.515 104.755 123.225 ;
        RECT 104.925 122.335 105.255 123.045 ;
        RECT 105.425 122.515 105.685 123.225 ;
        RECT 105.875 122.335 106.165 123.500 ;
        RECT 107.410 123.475 107.585 124.145 ;
        RECT 107.755 123.645 107.995 124.295 ;
        RECT 108.645 124.290 108.895 124.715 ;
        RECT 109.065 124.460 109.395 124.885 ;
        RECT 109.565 124.465 110.655 124.715 ;
        RECT 110.845 124.465 111.935 124.715 ;
        RECT 109.565 124.290 109.735 124.465 ;
        RECT 108.645 124.120 109.735 124.290 ;
        RECT 109.905 124.125 111.595 124.295 ;
        RECT 111.765 124.290 111.935 124.465 ;
        RECT 112.105 124.460 112.435 124.885 ;
        RECT 112.605 124.290 112.925 124.715 ;
        RECT 108.700 123.865 109.330 123.895 ;
        RECT 108.695 123.695 109.330 123.865 ;
        RECT 109.620 123.695 110.250 123.895 ;
        RECT 110.420 123.485 110.710 124.125 ;
        RECT 111.765 124.120 112.925 124.290 ;
        RECT 110.995 123.695 111.650 123.895 ;
        RECT 111.940 123.865 113.050 123.895 ;
        RECT 111.915 123.695 113.050 123.865 ;
        RECT 106.345 123.115 107.240 123.445 ;
        RECT 107.410 123.285 107.995 123.475 ;
        RECT 106.345 122.945 107.550 123.115 ;
        RECT 106.345 122.515 106.675 122.945 ;
        RECT 106.855 122.335 107.050 122.775 ;
        RECT 107.220 122.515 107.550 122.945 ;
        RECT 107.720 122.515 107.995 123.285 ;
        RECT 108.645 123.315 110.710 123.485 ;
        RECT 108.645 122.505 108.895 123.315 ;
        RECT 109.065 122.675 109.315 123.145 ;
        RECT 109.485 122.845 109.815 123.315 ;
        RECT 109.985 122.675 110.155 123.145 ;
        RECT 110.325 122.845 110.710 123.315 ;
        RECT 110.925 123.315 112.855 123.485 ;
        RECT 110.925 122.675 111.175 123.315 ;
        RECT 109.065 122.505 111.175 122.675 ;
        RECT 111.345 122.335 111.515 123.145 ;
        RECT 111.685 122.505 112.015 123.315 ;
        RECT 112.185 122.335 112.355 123.145 ;
        RECT 112.525 122.505 112.855 123.315 ;
        RECT 113.250 122.515 113.530 124.705 ;
        RECT 113.730 124.515 114.460 124.885 ;
        RECT 115.040 124.345 115.470 124.705 ;
        RECT 113.730 124.155 115.470 124.345 ;
        RECT 113.730 123.645 113.990 124.155 ;
        RECT 113.720 122.335 114.005 123.475 ;
        RECT 114.200 123.355 114.460 123.975 ;
        RECT 114.655 123.355 115.080 123.975 ;
        RECT 115.250 123.925 115.470 124.155 ;
        RECT 115.640 124.105 115.885 124.885 ;
        RECT 115.250 123.625 115.795 123.925 ;
        RECT 116.085 123.805 116.315 124.705 ;
        RECT 114.270 122.985 115.295 123.185 ;
        RECT 114.270 122.515 114.440 122.985 ;
        RECT 114.615 122.335 114.945 122.815 ;
        RECT 115.115 122.515 115.295 122.985 ;
        RECT 115.465 122.515 115.795 123.625 ;
        RECT 115.975 123.125 116.315 123.805 ;
        RECT 116.495 123.305 116.725 124.645 ;
        RECT 116.935 124.075 117.175 124.885 ;
        RECT 117.345 124.075 117.675 124.715 ;
        RECT 117.845 124.075 118.115 124.885 ;
        RECT 116.915 123.645 117.265 123.895 ;
        RECT 117.435 123.475 117.605 124.075 ;
        RECT 117.775 123.645 118.125 123.895 ;
        RECT 116.925 123.305 117.605 123.475 ;
        RECT 115.975 122.925 116.725 123.125 ;
        RECT 115.965 122.335 116.315 122.745 ;
        RECT 116.485 122.535 116.725 122.925 ;
        RECT 116.925 122.520 117.255 123.305 ;
        RECT 117.785 122.335 118.115 123.475 ;
        RECT 118.765 122.515 119.025 124.705 ;
        RECT 119.285 124.515 119.955 124.885 ;
        RECT 120.135 124.335 120.445 124.705 ;
        RECT 119.215 124.135 120.445 124.335 ;
        RECT 119.215 123.465 119.505 124.135 ;
        RECT 120.625 123.955 120.855 124.595 ;
        RECT 121.035 124.155 121.325 124.885 ;
        RECT 121.535 124.495 122.710 124.715 ;
        RECT 121.515 124.075 122.290 124.325 ;
        RECT 122.460 124.245 122.710 124.495 ;
        RECT 122.880 124.415 123.050 124.885 ;
        RECT 123.220 124.245 123.550 124.715 ;
        RECT 119.685 123.645 120.150 123.955 ;
        RECT 120.330 123.645 120.855 123.955 ;
        RECT 121.035 123.645 121.335 123.975 ;
        RECT 119.215 123.245 119.985 123.465 ;
        RECT 119.195 122.335 119.535 123.065 ;
        RECT 119.715 122.515 119.985 123.245 ;
        RECT 120.165 123.225 121.325 123.465 ;
        RECT 120.165 122.515 120.395 123.225 ;
        RECT 120.565 122.335 120.895 123.045 ;
        RECT 121.065 122.515 121.325 123.225 ;
        RECT 121.515 123.185 121.745 124.075 ;
        RECT 122.460 124.065 123.550 124.245 ;
        RECT 123.860 124.065 124.030 124.885 ;
        RECT 124.200 124.245 124.530 124.715 ;
        RECT 124.700 124.415 124.870 124.885 ;
        RECT 125.040 124.245 125.405 124.715 ;
        RECT 125.575 124.415 125.745 124.885 ;
        RECT 126.015 124.495 127.325 124.665 ;
        RECT 126.435 124.245 126.765 124.325 ;
        RECT 124.200 124.065 126.765 124.245 ;
        RECT 121.915 123.685 122.390 123.895 ;
        RECT 122.685 123.695 124.135 123.895 ;
        RECT 122.220 123.525 122.390 123.685 ;
        RECT 124.360 123.685 125.385 123.895 ;
        RECT 126.065 123.725 126.725 123.895 ;
        RECT 124.360 123.525 124.530 123.685 ;
        RECT 122.220 123.355 124.530 123.525 ;
        RECT 126.065 123.515 126.235 123.725 ;
        RECT 126.935 123.555 127.325 124.495 ;
        RECT 127.515 124.075 127.755 124.885 ;
        RECT 127.925 124.075 128.255 124.715 ;
        RECT 128.425 124.075 128.695 124.885 ;
        RECT 129.820 124.495 130.150 124.885 ;
        RECT 130.320 124.325 130.545 124.705 ;
        RECT 127.495 123.645 127.845 123.895 ;
        RECT 124.740 123.345 126.235 123.515 ;
        RECT 126.475 123.345 127.325 123.555 ;
        RECT 128.015 123.475 128.185 124.075 ;
        RECT 128.355 123.645 128.705 123.895 ;
        RECT 129.805 123.645 130.045 124.295 ;
        RECT 130.215 124.145 130.545 124.325 ;
        RECT 130.215 123.475 130.390 124.145 ;
        RECT 130.745 123.975 130.975 124.595 ;
        RECT 131.155 124.155 131.455 124.885 ;
        RECT 131.635 124.160 131.925 124.885 ;
        RECT 132.105 124.145 132.435 124.885 ;
        RECT 132.615 124.355 132.935 124.715 ;
        RECT 133.140 124.525 133.470 124.885 ;
        RECT 133.930 124.355 134.275 124.715 ;
        RECT 132.615 124.185 134.275 124.355 ;
        RECT 130.560 123.645 130.975 123.975 ;
        RECT 131.155 123.645 131.450 123.975 ;
        RECT 124.740 123.185 124.910 123.345 ;
        RECT 121.515 123.015 124.910 123.185 ;
        RECT 126.475 123.175 126.725 123.345 ;
        RECT 127.505 123.305 128.185 123.475 ;
        RECT 121.515 123.005 123.510 123.015 ;
        RECT 121.515 122.505 121.830 123.005 ;
        RECT 122.000 122.335 122.250 122.835 ;
        RECT 122.420 122.505 122.670 123.005 ;
        RECT 122.840 122.335 123.090 122.835 ;
        RECT 123.260 122.505 123.510 123.005 ;
        RECT 125.155 123.005 126.725 123.175 ;
        RECT 125.155 122.845 125.365 123.005 ;
        RECT 126.475 122.845 126.725 123.005 ;
        RECT 123.820 122.505 124.070 122.845 ;
        RECT 124.240 122.335 124.490 122.835 ;
        RECT 124.660 122.675 124.985 122.845 ;
        RECT 125.535 122.675 125.785 122.835 ;
        RECT 124.660 122.505 125.785 122.675 ;
        RECT 126.055 122.335 126.305 122.835 ;
        RECT 126.895 122.335 127.325 123.175 ;
        RECT 127.505 122.520 127.835 123.305 ;
        RECT 128.365 122.335 128.695 123.475 ;
        RECT 129.805 123.285 130.390 123.475 ;
        RECT 129.805 122.515 130.080 123.285 ;
        RECT 130.560 123.115 131.455 123.445 ;
        RECT 130.250 122.945 131.455 123.115 ;
        RECT 130.250 122.515 130.580 122.945 ;
        RECT 130.750 122.335 130.945 122.775 ;
        RECT 131.125 122.515 131.455 122.945 ;
        RECT 131.635 122.335 131.925 123.500 ;
        RECT 132.155 123.345 132.430 123.975 ;
        RECT 132.140 122.685 132.445 123.175 ;
        RECT 132.615 122.855 132.915 124.185 ;
        RECT 134.835 124.105 135.130 124.885 ;
        RECT 135.335 124.195 135.575 124.715 ;
        RECT 135.745 124.390 136.140 124.885 ;
        RECT 136.705 124.555 136.875 124.700 ;
        RECT 136.500 124.360 136.875 124.555 ;
        RECT 133.295 123.725 133.625 123.895 ;
        RECT 133.300 123.475 133.625 123.725 ;
        RECT 133.805 123.645 134.415 123.975 ;
        RECT 134.585 123.475 135.085 123.935 ;
        RECT 133.300 123.295 135.085 123.475 ;
        RECT 135.335 123.390 135.510 124.195 ;
        RECT 136.500 124.025 136.670 124.360 ;
        RECT 137.155 124.315 137.395 124.690 ;
        RECT 137.565 124.380 137.900 124.885 ;
        RECT 138.075 124.340 143.420 124.885 ;
        RECT 143.595 124.340 148.940 124.885 ;
        RECT 149.115 124.340 154.460 124.885 ;
        RECT 137.155 124.165 137.375 124.315 ;
        RECT 135.685 123.665 136.670 124.025 ;
        RECT 136.840 123.835 137.375 124.165 ;
        RECT 135.685 123.645 136.970 123.665 ;
        RECT 136.110 123.495 136.970 123.645 ;
        RECT 133.085 122.945 135.120 123.115 ;
        RECT 133.085 122.685 133.415 122.945 ;
        RECT 134.010 122.865 135.120 122.945 ;
        RECT 132.140 122.505 133.415 122.685 ;
        RECT 133.585 122.335 133.755 122.775 ;
        RECT 134.010 122.505 134.180 122.865 ;
        RECT 134.360 122.335 134.690 122.695 ;
        RECT 134.860 122.505 135.120 122.865 ;
        RECT 135.335 122.605 135.640 123.390 ;
        RECT 135.815 123.015 136.510 123.325 ;
        RECT 135.820 122.335 136.505 122.805 ;
        RECT 136.685 122.550 136.970 123.495 ;
        RECT 137.140 123.185 137.375 123.835 ;
        RECT 137.545 123.355 137.845 124.205 ;
        RECT 139.660 123.510 140.000 124.340 ;
        RECT 137.140 122.955 137.815 123.185 ;
        RECT 137.145 122.335 137.475 122.785 ;
        RECT 137.645 122.525 137.815 122.955 ;
        RECT 141.480 122.770 141.830 124.020 ;
        RECT 145.180 123.510 145.520 124.340 ;
        RECT 147.000 122.770 147.350 124.020 ;
        RECT 150.700 123.510 151.040 124.340 ;
        RECT 154.635 124.115 156.305 124.885 ;
        RECT 156.935 124.135 158.145 124.885 ;
        RECT 152.520 122.770 152.870 124.020 ;
        RECT 154.635 123.595 155.385 124.115 ;
        RECT 155.555 123.425 156.305 123.945 ;
        RECT 138.075 122.335 143.420 122.770 ;
        RECT 143.595 122.335 148.940 122.770 ;
        RECT 149.115 122.335 154.460 122.770 ;
        RECT 154.635 122.335 156.305 123.425 ;
        RECT 156.935 123.425 157.455 123.965 ;
        RECT 157.625 123.595 158.145 124.135 ;
        RECT 156.935 122.335 158.145 123.425 ;
        RECT 2.750 122.165 158.230 122.335 ;
        RECT 2.835 121.075 4.045 122.165 ;
        RECT 4.215 121.730 9.560 122.165 ;
        RECT 9.735 121.730 15.080 122.165 ;
        RECT 2.835 120.365 3.355 120.905 ;
        RECT 3.525 120.535 4.045 121.075 ;
        RECT 2.835 119.615 4.045 120.365 ;
        RECT 5.800 120.160 6.140 120.990 ;
        RECT 7.620 120.480 7.970 121.730 ;
        RECT 11.320 120.160 11.660 120.990 ;
        RECT 13.140 120.480 13.490 121.730 ;
        RECT 15.715 121.000 16.005 122.165 ;
        RECT 16.175 121.730 21.520 122.165 ;
        RECT 21.695 121.730 27.040 122.165 ;
        RECT 27.215 121.730 32.560 122.165 ;
        RECT 32.735 121.730 38.080 122.165 ;
        RECT 4.215 119.615 9.560 120.160 ;
        RECT 9.735 119.615 15.080 120.160 ;
        RECT 15.715 119.615 16.005 120.340 ;
        RECT 17.760 120.160 18.100 120.990 ;
        RECT 19.580 120.480 19.930 121.730 ;
        RECT 23.280 120.160 23.620 120.990 ;
        RECT 25.100 120.480 25.450 121.730 ;
        RECT 28.800 120.160 29.140 120.990 ;
        RECT 30.620 120.480 30.970 121.730 ;
        RECT 34.320 120.160 34.660 120.990 ;
        RECT 36.140 120.480 36.490 121.730 ;
        RECT 38.255 121.075 40.845 122.165 ;
        RECT 38.255 120.385 39.465 120.905 ;
        RECT 39.635 120.555 40.845 121.075 ;
        RECT 41.475 121.000 41.765 122.165 ;
        RECT 41.935 121.730 47.280 122.165 ;
        RECT 47.455 121.730 52.800 122.165 ;
        RECT 52.975 121.730 58.320 122.165 ;
        RECT 58.495 121.730 63.840 122.165 ;
        RECT 16.175 119.615 21.520 120.160 ;
        RECT 21.695 119.615 27.040 120.160 ;
        RECT 27.215 119.615 32.560 120.160 ;
        RECT 32.735 119.615 38.080 120.160 ;
        RECT 38.255 119.615 40.845 120.385 ;
        RECT 41.475 119.615 41.765 120.340 ;
        RECT 43.520 120.160 43.860 120.990 ;
        RECT 45.340 120.480 45.690 121.730 ;
        RECT 49.040 120.160 49.380 120.990 ;
        RECT 50.860 120.480 51.210 121.730 ;
        RECT 54.560 120.160 54.900 120.990 ;
        RECT 56.380 120.480 56.730 121.730 ;
        RECT 60.080 120.160 60.420 120.990 ;
        RECT 61.900 120.480 62.250 121.730 ;
        RECT 64.015 121.075 66.605 122.165 ;
        RECT 64.015 120.385 65.225 120.905 ;
        RECT 65.395 120.555 66.605 121.075 ;
        RECT 67.235 121.000 67.525 122.165 ;
        RECT 67.695 121.075 71.205 122.165 ;
        RECT 71.375 121.075 72.585 122.165 ;
        RECT 67.695 120.385 69.345 120.905 ;
        RECT 69.515 120.555 71.205 121.075 ;
        RECT 41.935 119.615 47.280 120.160 ;
        RECT 47.455 119.615 52.800 120.160 ;
        RECT 52.975 119.615 58.320 120.160 ;
        RECT 58.495 119.615 63.840 120.160 ;
        RECT 64.015 119.615 66.605 120.385 ;
        RECT 67.235 119.615 67.525 120.340 ;
        RECT 67.695 119.615 71.205 120.385 ;
        RECT 71.375 120.365 71.895 120.905 ;
        RECT 72.065 120.535 72.585 121.075 ;
        RECT 72.790 121.375 73.325 121.995 ;
        RECT 71.375 119.615 72.585 120.365 ;
        RECT 72.790 120.355 73.105 121.375 ;
        RECT 73.495 121.365 73.825 122.165 ;
        RECT 74.310 121.195 74.700 121.370 ;
        RECT 73.275 121.025 74.700 121.195 ;
        RECT 75.515 121.065 75.835 121.995 ;
        RECT 76.015 121.485 76.415 121.995 ;
        RECT 76.585 121.655 76.755 122.165 ;
        RECT 76.925 121.485 77.255 121.995 ;
        RECT 76.015 121.315 77.255 121.485 ;
        RECT 77.425 121.315 77.595 122.165 ;
        RECT 78.185 121.315 78.565 121.995 ;
        RECT 78.735 121.730 84.080 122.165 ;
        RECT 73.275 120.525 73.445 121.025 ;
        RECT 72.790 119.785 73.405 120.355 ;
        RECT 73.695 120.295 73.960 120.855 ;
        RECT 74.130 120.125 74.300 121.025 ;
        RECT 75.515 120.895 76.145 121.065 ;
        RECT 74.470 120.295 74.825 120.855 ;
        RECT 73.575 119.615 73.790 120.125 ;
        RECT 74.020 119.795 74.300 120.125 ;
        RECT 74.480 119.615 74.720 120.125 ;
        RECT 75.515 119.615 75.805 120.450 ;
        RECT 75.975 120.015 76.145 120.895 ;
        RECT 76.920 120.975 78.225 121.145 ;
        RECT 76.315 120.355 76.545 120.855 ;
        RECT 76.920 120.775 77.090 120.975 ;
        RECT 76.715 120.605 77.090 120.775 ;
        RECT 77.260 120.605 77.810 120.805 ;
        RECT 77.980 120.525 78.225 120.975 ;
        RECT 78.395 120.355 78.565 121.315 ;
        RECT 76.315 120.185 78.565 120.355 ;
        RECT 75.975 119.845 76.930 120.015 ;
        RECT 77.345 119.615 77.675 120.005 ;
        RECT 77.845 119.865 78.015 120.185 ;
        RECT 80.320 120.160 80.660 120.990 ;
        RECT 82.140 120.480 82.490 121.730 ;
        RECT 84.255 121.315 84.635 121.995 ;
        RECT 85.225 121.315 85.395 122.165 ;
        RECT 85.565 121.485 85.895 121.995 ;
        RECT 86.065 121.655 86.235 122.165 ;
        RECT 86.405 121.485 86.805 121.995 ;
        RECT 85.565 121.315 86.805 121.485 ;
        RECT 84.255 120.355 84.425 121.315 ;
        RECT 84.595 120.975 85.900 121.145 ;
        RECT 86.985 121.065 87.305 121.995 ;
        RECT 87.475 121.075 90.065 122.165 ;
        RECT 84.595 120.525 84.840 120.975 ;
        RECT 85.010 120.605 85.560 120.805 ;
        RECT 85.730 120.775 85.900 120.975 ;
        RECT 86.675 120.895 87.305 121.065 ;
        RECT 85.730 120.605 86.105 120.775 ;
        RECT 86.275 120.355 86.505 120.855 ;
        RECT 84.255 120.185 86.505 120.355 ;
        RECT 78.185 119.615 78.515 120.005 ;
        RECT 78.735 119.615 84.080 120.160 ;
        RECT 84.305 119.615 84.635 120.005 ;
        RECT 84.805 119.865 84.975 120.185 ;
        RECT 86.675 120.015 86.845 120.895 ;
        RECT 85.145 119.615 85.475 120.005 ;
        RECT 85.890 119.845 86.845 120.015 ;
        RECT 87.015 119.615 87.305 120.450 ;
        RECT 87.475 120.385 88.685 120.905 ;
        RECT 88.855 120.555 90.065 121.075 ;
        RECT 90.730 121.375 91.265 121.995 ;
        RECT 87.475 119.615 90.065 120.385 ;
        RECT 90.730 120.355 91.045 121.375 ;
        RECT 91.435 121.365 91.765 122.165 ;
        RECT 92.250 121.195 92.640 121.370 ;
        RECT 91.215 121.025 92.640 121.195 ;
        RECT 91.215 120.525 91.385 121.025 ;
        RECT 90.730 119.785 91.345 120.355 ;
        RECT 91.635 120.295 91.900 120.855 ;
        RECT 92.070 120.125 92.240 121.025 ;
        RECT 92.995 121.000 93.285 122.165 ;
        RECT 94.375 121.025 94.650 121.995 ;
        RECT 94.860 121.365 95.140 122.165 ;
        RECT 95.310 121.655 96.925 121.985 ;
        RECT 95.310 121.315 96.485 121.485 ;
        RECT 95.310 121.195 95.480 121.315 ;
        RECT 94.820 121.025 95.480 121.195 ;
        RECT 92.410 120.295 92.765 120.855 ;
        RECT 91.515 119.615 91.730 120.125 ;
        RECT 91.960 119.795 92.240 120.125 ;
        RECT 92.420 119.615 92.660 120.125 ;
        RECT 92.995 119.615 93.285 120.340 ;
        RECT 94.375 120.290 94.545 121.025 ;
        RECT 94.820 120.855 94.990 121.025 ;
        RECT 95.740 120.855 95.985 121.145 ;
        RECT 96.155 121.025 96.485 121.315 ;
        RECT 96.745 120.855 96.915 121.415 ;
        RECT 97.165 121.025 97.425 122.165 ;
        RECT 97.595 121.025 97.875 122.165 ;
        RECT 98.045 121.015 98.375 121.995 ;
        RECT 98.545 121.025 98.805 122.165 ;
        RECT 99.895 121.065 100.215 121.995 ;
        RECT 100.395 121.485 100.795 121.995 ;
        RECT 100.965 121.655 101.135 122.165 ;
        RECT 101.305 121.485 101.635 121.995 ;
        RECT 100.395 121.315 101.635 121.485 ;
        RECT 101.805 121.315 101.975 122.165 ;
        RECT 102.565 121.315 102.945 121.995 ;
        RECT 103.115 121.655 103.415 122.165 ;
        RECT 103.585 121.485 103.915 121.995 ;
        RECT 104.085 121.655 104.715 122.165 ;
        RECT 105.295 121.655 105.675 121.825 ;
        RECT 105.845 121.655 106.145 122.165 ;
        RECT 105.505 121.485 105.675 121.655 ;
        RECT 94.715 120.525 94.990 120.855 ;
        RECT 95.160 120.525 95.985 120.855 ;
        RECT 96.200 120.525 96.915 120.855 ;
        RECT 97.085 120.605 97.420 120.855 ;
        RECT 97.605 120.585 97.940 120.855 ;
        RECT 94.820 120.355 94.990 120.525 ;
        RECT 96.665 120.435 96.915 120.525 ;
        RECT 94.375 119.945 94.650 120.290 ;
        RECT 94.820 120.185 96.485 120.355 ;
        RECT 94.840 119.615 95.215 120.015 ;
        RECT 95.385 119.835 95.555 120.185 ;
        RECT 95.725 119.615 96.055 120.015 ;
        RECT 96.225 119.785 96.485 120.185 ;
        RECT 96.665 120.015 96.995 120.435 ;
        RECT 97.165 119.615 97.425 120.435 ;
        RECT 98.110 120.415 98.280 121.015 ;
        RECT 99.895 120.895 100.525 121.065 ;
        RECT 98.450 120.605 98.785 120.855 ;
        RECT 97.595 119.615 97.905 120.415 ;
        RECT 98.110 119.785 98.805 120.415 ;
        RECT 99.895 119.615 100.185 120.450 ;
        RECT 100.355 120.015 100.525 120.895 ;
        RECT 101.300 120.975 102.605 121.145 ;
        RECT 100.695 120.355 100.925 120.855 ;
        RECT 101.300 120.775 101.470 120.975 ;
        RECT 101.095 120.605 101.470 120.775 ;
        RECT 101.640 120.605 102.190 120.805 ;
        RECT 102.360 120.525 102.605 120.975 ;
        RECT 102.775 120.355 102.945 121.315 ;
        RECT 100.695 120.185 102.945 120.355 ;
        RECT 103.115 121.315 105.335 121.485 ;
        RECT 103.115 120.355 103.285 121.315 ;
        RECT 103.455 120.975 104.995 121.145 ;
        RECT 103.455 120.525 103.700 120.975 ;
        RECT 103.960 120.605 104.655 120.805 ;
        RECT 104.825 120.775 104.995 120.975 ;
        RECT 105.165 121.115 105.335 121.315 ;
        RECT 105.505 121.285 106.165 121.485 ;
        RECT 105.165 120.945 105.825 121.115 ;
        RECT 104.825 120.605 105.425 120.775 ;
        RECT 105.655 120.525 105.825 120.945 ;
        RECT 100.355 119.845 101.310 120.015 ;
        RECT 101.725 119.615 102.055 120.005 ;
        RECT 102.225 119.865 102.395 120.185 ;
        RECT 102.565 119.615 102.895 120.005 ;
        RECT 103.115 119.810 103.580 120.355 ;
        RECT 104.085 119.615 104.255 120.435 ;
        RECT 104.425 120.355 105.335 120.435 ;
        RECT 105.995 120.355 106.165 121.285 ;
        RECT 106.335 121.025 106.615 122.165 ;
        RECT 106.785 121.015 107.115 121.995 ;
        RECT 107.285 121.025 107.545 122.165 ;
        RECT 107.715 121.075 108.925 122.165 ;
        RECT 109.095 121.655 109.395 122.165 ;
        RECT 109.565 121.485 109.895 121.995 ;
        RECT 110.065 121.655 110.695 122.165 ;
        RECT 111.275 121.655 111.655 121.825 ;
        RECT 111.825 121.655 112.125 122.165 ;
        RECT 112.315 121.730 117.660 122.165 ;
        RECT 111.485 121.485 111.655 121.655 ;
        RECT 106.345 120.585 106.680 120.855 ;
        RECT 106.850 120.465 107.020 121.015 ;
        RECT 107.190 120.605 107.525 120.855 ;
        RECT 106.850 120.415 107.025 120.465 ;
        RECT 104.425 120.265 105.675 120.355 ;
        RECT 104.425 119.785 104.755 120.265 ;
        RECT 105.165 120.185 105.675 120.265 ;
        RECT 104.925 119.615 105.275 120.005 ;
        RECT 105.445 119.785 105.675 120.185 ;
        RECT 105.845 119.875 106.165 120.355 ;
        RECT 106.335 119.615 106.645 120.415 ;
        RECT 106.850 119.785 107.545 120.415 ;
        RECT 107.715 120.365 108.235 120.905 ;
        RECT 108.405 120.535 108.925 121.075 ;
        RECT 109.095 121.315 111.315 121.485 ;
        RECT 107.715 119.615 108.925 120.365 ;
        RECT 109.095 120.355 109.265 121.315 ;
        RECT 109.435 120.975 110.975 121.145 ;
        RECT 109.435 120.525 109.680 120.975 ;
        RECT 109.940 120.605 110.635 120.805 ;
        RECT 110.805 120.775 110.975 120.975 ;
        RECT 111.145 121.115 111.315 121.315 ;
        RECT 111.485 121.285 112.145 121.485 ;
        RECT 111.145 120.945 111.805 121.115 ;
        RECT 110.805 120.605 111.405 120.775 ;
        RECT 111.635 120.525 111.805 120.945 ;
        RECT 109.095 119.810 109.560 120.355 ;
        RECT 110.065 119.615 110.235 120.435 ;
        RECT 110.405 120.355 111.315 120.435 ;
        RECT 111.975 120.355 112.145 121.285 ;
        RECT 110.405 120.265 111.655 120.355 ;
        RECT 110.405 119.785 110.735 120.265 ;
        RECT 111.145 120.185 111.655 120.265 ;
        RECT 110.905 119.615 111.255 120.005 ;
        RECT 111.425 119.785 111.655 120.185 ;
        RECT 111.825 119.875 112.145 120.355 ;
        RECT 113.900 120.160 114.240 120.990 ;
        RECT 115.720 120.480 116.070 121.730 ;
        RECT 118.755 121.000 119.045 122.165 ;
        RECT 119.215 121.075 121.805 122.165 ;
        RECT 119.215 120.385 120.425 120.905 ;
        RECT 120.595 120.555 121.805 121.075 ;
        RECT 121.975 121.065 122.295 121.995 ;
        RECT 122.475 121.485 122.875 121.995 ;
        RECT 123.045 121.655 123.215 122.165 ;
        RECT 123.385 121.485 123.715 121.995 ;
        RECT 122.475 121.315 123.715 121.485 ;
        RECT 123.885 121.315 124.055 122.165 ;
        RECT 124.645 121.315 125.025 121.995 ;
        RECT 121.975 120.895 122.605 121.065 ;
        RECT 112.315 119.615 117.660 120.160 ;
        RECT 118.755 119.615 119.045 120.340 ;
        RECT 119.215 119.615 121.805 120.385 ;
        RECT 121.975 119.615 122.265 120.450 ;
        RECT 122.435 120.015 122.605 120.895 ;
        RECT 123.380 120.975 124.685 121.145 ;
        RECT 122.775 120.355 123.005 120.855 ;
        RECT 123.380 120.775 123.550 120.975 ;
        RECT 123.175 120.605 123.550 120.775 ;
        RECT 123.720 120.605 124.270 120.805 ;
        RECT 124.440 120.525 124.685 120.975 ;
        RECT 124.855 120.355 125.025 121.315 ;
        RECT 125.195 121.025 125.455 122.165 ;
        RECT 125.625 121.015 125.955 121.995 ;
        RECT 126.125 121.025 126.405 122.165 ;
        RECT 126.615 121.025 126.845 122.165 ;
        RECT 127.015 121.015 127.345 121.995 ;
        RECT 127.515 121.025 127.725 122.165 ;
        RECT 127.955 121.075 131.465 122.165 ;
        RECT 132.100 121.365 132.355 122.165 ;
        RECT 132.555 121.315 132.885 121.995 ;
        RECT 125.215 120.605 125.550 120.855 ;
        RECT 125.720 120.415 125.890 121.015 ;
        RECT 126.060 120.585 126.395 120.855 ;
        RECT 126.595 120.605 126.925 120.855 ;
        RECT 122.775 120.185 125.025 120.355 ;
        RECT 122.435 119.845 123.390 120.015 ;
        RECT 123.805 119.615 124.135 120.005 ;
        RECT 124.305 119.865 124.475 120.185 ;
        RECT 124.645 119.615 124.975 120.005 ;
        RECT 125.195 119.785 125.890 120.415 ;
        RECT 126.095 119.615 126.405 120.415 ;
        RECT 126.615 119.615 126.845 120.435 ;
        RECT 127.095 120.415 127.345 121.015 ;
        RECT 127.015 119.785 127.345 120.415 ;
        RECT 127.515 119.615 127.725 120.435 ;
        RECT 127.955 120.385 129.605 120.905 ;
        RECT 129.775 120.555 131.465 121.075 ;
        RECT 132.100 120.825 132.345 121.185 ;
        RECT 132.535 121.035 132.885 121.315 ;
        RECT 132.535 120.655 132.705 121.035 ;
        RECT 133.065 120.855 133.260 121.905 ;
        RECT 133.440 121.025 133.760 122.165 ;
        RECT 133.935 121.730 139.280 122.165 ;
        RECT 132.185 120.485 132.705 120.655 ;
        RECT 132.875 120.525 133.260 120.855 ;
        RECT 133.440 120.805 133.700 120.855 ;
        RECT 133.440 120.635 133.705 120.805 ;
        RECT 133.440 120.525 133.700 120.635 ;
        RECT 127.955 119.615 131.465 120.385 ;
        RECT 132.185 119.920 132.355 120.485 ;
        RECT 132.545 120.145 133.760 120.315 ;
        RECT 135.520 120.160 135.860 120.990 ;
        RECT 137.340 120.480 137.690 121.730 ;
        RECT 139.455 121.075 142.965 122.165 ;
        RECT 143.135 121.075 144.345 122.165 ;
        RECT 139.455 120.385 141.105 120.905 ;
        RECT 141.275 120.555 142.965 121.075 ;
        RECT 132.545 119.840 132.775 120.145 ;
        RECT 132.945 119.615 133.275 119.975 ;
        RECT 133.470 119.795 133.760 120.145 ;
        RECT 133.935 119.615 139.280 120.160 ;
        RECT 139.455 119.615 142.965 120.385 ;
        RECT 143.135 120.365 143.655 120.905 ;
        RECT 143.825 120.535 144.345 121.075 ;
        RECT 144.515 121.000 144.805 122.165 ;
        RECT 144.975 121.730 150.320 122.165 ;
        RECT 150.495 121.730 155.840 122.165 ;
        RECT 143.135 119.615 144.345 120.365 ;
        RECT 144.515 119.615 144.805 120.340 ;
        RECT 146.560 120.160 146.900 120.990 ;
        RECT 148.380 120.480 148.730 121.730 ;
        RECT 152.080 120.160 152.420 120.990 ;
        RECT 153.900 120.480 154.250 121.730 ;
        RECT 156.935 121.075 158.145 122.165 ;
        RECT 156.935 120.535 157.455 121.075 ;
        RECT 157.625 120.365 158.145 120.905 ;
        RECT 144.975 119.615 150.320 120.160 ;
        RECT 150.495 119.615 155.840 120.160 ;
        RECT 156.935 119.615 158.145 120.365 ;
        RECT 2.750 119.445 158.230 119.615 ;
        RECT 2.835 118.695 4.045 119.445 ;
        RECT 4.215 118.900 9.560 119.445 ;
        RECT 9.735 118.900 15.080 119.445 ;
        RECT 15.255 118.900 20.600 119.445 ;
        RECT 20.775 118.900 26.120 119.445 ;
        RECT 2.835 118.155 3.355 118.695 ;
        RECT 3.525 117.985 4.045 118.525 ;
        RECT 5.800 118.070 6.140 118.900 ;
        RECT 2.835 116.895 4.045 117.985 ;
        RECT 7.620 117.330 7.970 118.580 ;
        RECT 11.320 118.070 11.660 118.900 ;
        RECT 13.140 117.330 13.490 118.580 ;
        RECT 16.840 118.070 17.180 118.900 ;
        RECT 18.660 117.330 19.010 118.580 ;
        RECT 22.360 118.070 22.700 118.900 ;
        RECT 26.295 118.675 27.965 119.445 ;
        RECT 28.595 118.720 28.885 119.445 ;
        RECT 29.055 118.900 34.400 119.445 ;
        RECT 34.575 118.900 39.920 119.445 ;
        RECT 40.095 118.900 45.440 119.445 ;
        RECT 45.615 118.900 50.960 119.445 ;
        RECT 24.180 117.330 24.530 118.580 ;
        RECT 26.295 118.155 27.045 118.675 ;
        RECT 27.215 117.985 27.965 118.505 ;
        RECT 30.640 118.070 30.980 118.900 ;
        RECT 4.215 116.895 9.560 117.330 ;
        RECT 9.735 116.895 15.080 117.330 ;
        RECT 15.255 116.895 20.600 117.330 ;
        RECT 20.775 116.895 26.120 117.330 ;
        RECT 26.295 116.895 27.965 117.985 ;
        RECT 28.595 116.895 28.885 118.060 ;
        RECT 32.460 117.330 32.810 118.580 ;
        RECT 36.160 118.070 36.500 118.900 ;
        RECT 37.980 117.330 38.330 118.580 ;
        RECT 41.680 118.070 42.020 118.900 ;
        RECT 43.500 117.330 43.850 118.580 ;
        RECT 47.200 118.070 47.540 118.900 ;
        RECT 51.135 118.675 53.725 119.445 ;
        RECT 54.355 118.720 54.645 119.445 ;
        RECT 54.815 118.900 60.160 119.445 ;
        RECT 60.335 118.900 65.680 119.445 ;
        RECT 65.855 118.900 71.200 119.445 ;
        RECT 71.375 118.900 76.720 119.445 ;
        RECT 49.020 117.330 49.370 118.580 ;
        RECT 51.135 118.155 52.345 118.675 ;
        RECT 52.515 117.985 53.725 118.505 ;
        RECT 56.400 118.070 56.740 118.900 ;
        RECT 29.055 116.895 34.400 117.330 ;
        RECT 34.575 116.895 39.920 117.330 ;
        RECT 40.095 116.895 45.440 117.330 ;
        RECT 45.615 116.895 50.960 117.330 ;
        RECT 51.135 116.895 53.725 117.985 ;
        RECT 54.355 116.895 54.645 118.060 ;
        RECT 58.220 117.330 58.570 118.580 ;
        RECT 61.920 118.070 62.260 118.900 ;
        RECT 63.740 117.330 64.090 118.580 ;
        RECT 67.440 118.070 67.780 118.900 ;
        RECT 69.260 117.330 69.610 118.580 ;
        RECT 72.960 118.070 73.300 118.900 ;
        RECT 76.895 118.675 79.485 119.445 ;
        RECT 80.115 118.720 80.405 119.445 ;
        RECT 80.575 118.900 85.920 119.445 ;
        RECT 86.095 118.900 91.440 119.445 ;
        RECT 74.780 117.330 75.130 118.580 ;
        RECT 76.895 118.155 78.105 118.675 ;
        RECT 78.275 117.985 79.485 118.505 ;
        RECT 82.160 118.070 82.500 118.900 ;
        RECT 54.815 116.895 60.160 117.330 ;
        RECT 60.335 116.895 65.680 117.330 ;
        RECT 65.855 116.895 71.200 117.330 ;
        RECT 71.375 116.895 76.720 117.330 ;
        RECT 76.895 116.895 79.485 117.985 ;
        RECT 80.115 116.895 80.405 118.060 ;
        RECT 83.980 117.330 84.330 118.580 ;
        RECT 87.680 118.070 88.020 118.900 ;
        RECT 91.615 118.675 94.205 119.445 ;
        RECT 94.375 118.685 95.085 119.275 ;
        RECT 95.595 118.915 95.925 119.275 ;
        RECT 96.125 119.085 96.455 119.445 ;
        RECT 96.625 118.915 96.955 119.275 ;
        RECT 95.595 118.705 96.955 118.915 ;
        RECT 89.500 117.330 89.850 118.580 ;
        RECT 91.615 118.155 92.825 118.675 ;
        RECT 92.995 117.985 94.205 118.505 ;
        RECT 80.575 116.895 85.920 117.330 ;
        RECT 86.095 116.895 91.440 117.330 ;
        RECT 91.615 116.895 94.205 117.985 ;
        RECT 94.375 117.715 94.580 118.685 ;
        RECT 97.615 118.635 97.855 119.445 ;
        RECT 98.025 118.635 98.355 119.275 ;
        RECT 98.525 118.635 98.795 119.445 ;
        RECT 98.975 118.900 104.320 119.445 ;
        RECT 94.750 117.915 95.080 118.455 ;
        RECT 95.255 118.205 95.750 118.535 ;
        RECT 96.070 118.205 96.445 118.535 ;
        RECT 96.655 118.205 96.965 118.535 ;
        RECT 97.595 118.205 97.945 118.455 ;
        RECT 95.255 117.915 95.580 118.205 ;
        RECT 95.775 117.715 96.105 117.935 ;
        RECT 94.375 117.485 96.105 117.715 ;
        RECT 94.375 117.065 95.075 117.485 ;
        RECT 95.275 116.895 95.605 117.255 ;
        RECT 95.775 117.085 96.105 117.485 ;
        RECT 96.275 117.235 96.445 118.205 ;
        RECT 98.115 118.035 98.285 118.635 ;
        RECT 98.455 118.205 98.805 118.455 ;
        RECT 100.560 118.070 100.900 118.900 ;
        RECT 104.495 118.695 105.705 119.445 ;
        RECT 105.875 118.720 106.165 119.445 ;
        RECT 106.335 118.900 111.680 119.445 ;
        RECT 111.855 118.900 117.200 119.445 ;
        RECT 117.375 118.900 122.720 119.445 ;
        RECT 122.895 118.900 128.240 119.445 ;
        RECT 96.625 116.895 96.955 117.955 ;
        RECT 97.605 117.865 98.285 118.035 ;
        RECT 97.605 117.080 97.935 117.865 ;
        RECT 98.465 116.895 98.795 118.035 ;
        RECT 102.380 117.330 102.730 118.580 ;
        RECT 104.495 118.155 105.015 118.695 ;
        RECT 105.185 117.985 105.705 118.525 ;
        RECT 107.920 118.070 108.260 118.900 ;
        RECT 98.975 116.895 104.320 117.330 ;
        RECT 104.495 116.895 105.705 117.985 ;
        RECT 105.875 116.895 106.165 118.060 ;
        RECT 109.740 117.330 110.090 118.580 ;
        RECT 113.440 118.070 113.780 118.900 ;
        RECT 115.260 117.330 115.610 118.580 ;
        RECT 118.960 118.070 119.300 118.900 ;
        RECT 120.780 117.330 121.130 118.580 ;
        RECT 124.480 118.070 124.820 118.900 ;
        RECT 128.415 118.675 131.005 119.445 ;
        RECT 131.635 118.720 131.925 119.445 ;
        RECT 132.095 118.900 137.440 119.445 ;
        RECT 137.615 118.900 142.960 119.445 ;
        RECT 143.135 118.900 148.480 119.445 ;
        RECT 148.655 118.900 154.000 119.445 ;
        RECT 126.300 117.330 126.650 118.580 ;
        RECT 128.415 118.155 129.625 118.675 ;
        RECT 129.795 117.985 131.005 118.505 ;
        RECT 133.680 118.070 134.020 118.900 ;
        RECT 106.335 116.895 111.680 117.330 ;
        RECT 111.855 116.895 117.200 117.330 ;
        RECT 117.375 116.895 122.720 117.330 ;
        RECT 122.895 116.895 128.240 117.330 ;
        RECT 128.415 116.895 131.005 117.985 ;
        RECT 131.635 116.895 131.925 118.060 ;
        RECT 135.500 117.330 135.850 118.580 ;
        RECT 139.200 118.070 139.540 118.900 ;
        RECT 141.020 117.330 141.370 118.580 ;
        RECT 144.720 118.070 145.060 118.900 ;
        RECT 146.540 117.330 146.890 118.580 ;
        RECT 150.240 118.070 150.580 118.900 ;
        RECT 154.175 118.675 156.765 119.445 ;
        RECT 156.935 118.695 158.145 119.445 ;
        RECT 152.060 117.330 152.410 118.580 ;
        RECT 154.175 118.155 155.385 118.675 ;
        RECT 155.555 117.985 156.765 118.505 ;
        RECT 132.095 116.895 137.440 117.330 ;
        RECT 137.615 116.895 142.960 117.330 ;
        RECT 143.135 116.895 148.480 117.330 ;
        RECT 148.655 116.895 154.000 117.330 ;
        RECT 154.175 116.895 156.765 117.985 ;
        RECT 156.935 117.985 157.455 118.525 ;
        RECT 157.625 118.155 158.145 118.695 ;
        RECT 156.935 116.895 158.145 117.985 ;
        RECT 2.750 116.725 158.230 116.895 ;
        RECT 2.835 115.635 4.045 116.725 ;
        RECT 4.215 116.290 9.560 116.725 ;
        RECT 9.735 116.290 15.080 116.725 ;
        RECT 2.835 114.925 3.355 115.465 ;
        RECT 3.525 115.095 4.045 115.635 ;
        RECT 2.835 114.175 4.045 114.925 ;
        RECT 5.800 114.720 6.140 115.550 ;
        RECT 7.620 115.040 7.970 116.290 ;
        RECT 11.320 114.720 11.660 115.550 ;
        RECT 13.140 115.040 13.490 116.290 ;
        RECT 15.715 115.560 16.005 116.725 ;
        RECT 16.175 116.290 21.520 116.725 ;
        RECT 21.695 116.290 27.040 116.725 ;
        RECT 4.215 114.175 9.560 114.720 ;
        RECT 9.735 114.175 15.080 114.720 ;
        RECT 15.715 114.175 16.005 114.900 ;
        RECT 17.760 114.720 18.100 115.550 ;
        RECT 19.580 115.040 19.930 116.290 ;
        RECT 23.280 114.720 23.620 115.550 ;
        RECT 25.100 115.040 25.450 116.290 ;
        RECT 27.215 115.635 28.425 116.725 ;
        RECT 27.215 114.925 27.735 115.465 ;
        RECT 27.905 115.095 28.425 115.635 ;
        RECT 28.595 115.560 28.885 116.725 ;
        RECT 29.055 116.290 34.400 116.725 ;
        RECT 34.575 116.290 39.920 116.725 ;
        RECT 16.175 114.175 21.520 114.720 ;
        RECT 21.695 114.175 27.040 114.720 ;
        RECT 27.215 114.175 28.425 114.925 ;
        RECT 28.595 114.175 28.885 114.900 ;
        RECT 30.640 114.720 30.980 115.550 ;
        RECT 32.460 115.040 32.810 116.290 ;
        RECT 36.160 114.720 36.500 115.550 ;
        RECT 37.980 115.040 38.330 116.290 ;
        RECT 40.095 115.635 41.305 116.725 ;
        RECT 40.095 114.925 40.615 115.465 ;
        RECT 40.785 115.095 41.305 115.635 ;
        RECT 41.475 115.560 41.765 116.725 ;
        RECT 41.935 116.290 47.280 116.725 ;
        RECT 47.455 116.290 52.800 116.725 ;
        RECT 29.055 114.175 34.400 114.720 ;
        RECT 34.575 114.175 39.920 114.720 ;
        RECT 40.095 114.175 41.305 114.925 ;
        RECT 41.475 114.175 41.765 114.900 ;
        RECT 43.520 114.720 43.860 115.550 ;
        RECT 45.340 115.040 45.690 116.290 ;
        RECT 49.040 114.720 49.380 115.550 ;
        RECT 50.860 115.040 51.210 116.290 ;
        RECT 52.975 115.635 54.185 116.725 ;
        RECT 52.975 114.925 53.495 115.465 ;
        RECT 53.665 115.095 54.185 115.635 ;
        RECT 54.355 115.560 54.645 116.725 ;
        RECT 54.815 116.290 60.160 116.725 ;
        RECT 60.335 116.290 65.680 116.725 ;
        RECT 41.935 114.175 47.280 114.720 ;
        RECT 47.455 114.175 52.800 114.720 ;
        RECT 52.975 114.175 54.185 114.925 ;
        RECT 54.355 114.175 54.645 114.900 ;
        RECT 56.400 114.720 56.740 115.550 ;
        RECT 58.220 115.040 58.570 116.290 ;
        RECT 61.920 114.720 62.260 115.550 ;
        RECT 63.740 115.040 64.090 116.290 ;
        RECT 65.855 115.635 67.065 116.725 ;
        RECT 65.855 114.925 66.375 115.465 ;
        RECT 66.545 115.095 67.065 115.635 ;
        RECT 67.235 115.560 67.525 116.725 ;
        RECT 67.695 116.290 73.040 116.725 ;
        RECT 73.215 116.290 78.560 116.725 ;
        RECT 54.815 114.175 60.160 114.720 ;
        RECT 60.335 114.175 65.680 114.720 ;
        RECT 65.855 114.175 67.065 114.925 ;
        RECT 67.235 114.175 67.525 114.900 ;
        RECT 69.280 114.720 69.620 115.550 ;
        RECT 71.100 115.040 71.450 116.290 ;
        RECT 74.800 114.720 75.140 115.550 ;
        RECT 76.620 115.040 76.970 116.290 ;
        RECT 78.735 115.635 79.945 116.725 ;
        RECT 78.735 114.925 79.255 115.465 ;
        RECT 79.425 115.095 79.945 115.635 ;
        RECT 80.115 115.560 80.405 116.725 ;
        RECT 80.575 116.290 85.920 116.725 ;
        RECT 86.095 116.290 91.440 116.725 ;
        RECT 67.695 114.175 73.040 114.720 ;
        RECT 73.215 114.175 78.560 114.720 ;
        RECT 78.735 114.175 79.945 114.925 ;
        RECT 80.115 114.175 80.405 114.900 ;
        RECT 82.160 114.720 82.500 115.550 ;
        RECT 83.980 115.040 84.330 116.290 ;
        RECT 87.680 114.720 88.020 115.550 ;
        RECT 89.500 115.040 89.850 116.290 ;
        RECT 91.615 115.635 92.825 116.725 ;
        RECT 91.615 114.925 92.135 115.465 ;
        RECT 92.305 115.095 92.825 115.635 ;
        RECT 92.995 115.560 93.285 116.725 ;
        RECT 93.455 116.290 98.800 116.725 ;
        RECT 98.975 116.290 104.320 116.725 ;
        RECT 80.575 114.175 85.920 114.720 ;
        RECT 86.095 114.175 91.440 114.720 ;
        RECT 91.615 114.175 92.825 114.925 ;
        RECT 92.995 114.175 93.285 114.900 ;
        RECT 95.040 114.720 95.380 115.550 ;
        RECT 96.860 115.040 97.210 116.290 ;
        RECT 100.560 114.720 100.900 115.550 ;
        RECT 102.380 115.040 102.730 116.290 ;
        RECT 104.495 115.635 105.705 116.725 ;
        RECT 104.495 114.925 105.015 115.465 ;
        RECT 105.185 115.095 105.705 115.635 ;
        RECT 105.875 115.560 106.165 116.725 ;
        RECT 106.335 116.290 111.680 116.725 ;
        RECT 111.855 116.290 117.200 116.725 ;
        RECT 93.455 114.175 98.800 114.720 ;
        RECT 98.975 114.175 104.320 114.720 ;
        RECT 104.495 114.175 105.705 114.925 ;
        RECT 105.875 114.175 106.165 114.900 ;
        RECT 107.920 114.720 108.260 115.550 ;
        RECT 109.740 115.040 110.090 116.290 ;
        RECT 113.440 114.720 113.780 115.550 ;
        RECT 115.260 115.040 115.610 116.290 ;
        RECT 117.375 115.635 118.585 116.725 ;
        RECT 117.375 114.925 117.895 115.465 ;
        RECT 118.065 115.095 118.585 115.635 ;
        RECT 118.755 115.560 119.045 116.725 ;
        RECT 119.215 116.290 124.560 116.725 ;
        RECT 124.735 116.290 130.080 116.725 ;
        RECT 106.335 114.175 111.680 114.720 ;
        RECT 111.855 114.175 117.200 114.720 ;
        RECT 117.375 114.175 118.585 114.925 ;
        RECT 118.755 114.175 119.045 114.900 ;
        RECT 120.800 114.720 121.140 115.550 ;
        RECT 122.620 115.040 122.970 116.290 ;
        RECT 126.320 114.720 126.660 115.550 ;
        RECT 128.140 115.040 128.490 116.290 ;
        RECT 130.255 115.635 131.465 116.725 ;
        RECT 130.255 114.925 130.775 115.465 ;
        RECT 130.945 115.095 131.465 115.635 ;
        RECT 131.635 115.560 131.925 116.725 ;
        RECT 132.095 116.290 137.440 116.725 ;
        RECT 137.615 116.290 142.960 116.725 ;
        RECT 119.215 114.175 124.560 114.720 ;
        RECT 124.735 114.175 130.080 114.720 ;
        RECT 130.255 114.175 131.465 114.925 ;
        RECT 131.635 114.175 131.925 114.900 ;
        RECT 133.680 114.720 134.020 115.550 ;
        RECT 135.500 115.040 135.850 116.290 ;
        RECT 139.200 114.720 139.540 115.550 ;
        RECT 141.020 115.040 141.370 116.290 ;
        RECT 143.135 115.635 144.345 116.725 ;
        RECT 143.135 114.925 143.655 115.465 ;
        RECT 143.825 115.095 144.345 115.635 ;
        RECT 144.515 115.560 144.805 116.725 ;
        RECT 144.975 116.290 150.320 116.725 ;
        RECT 150.495 116.290 155.840 116.725 ;
        RECT 132.095 114.175 137.440 114.720 ;
        RECT 137.615 114.175 142.960 114.720 ;
        RECT 143.135 114.175 144.345 114.925 ;
        RECT 144.515 114.175 144.805 114.900 ;
        RECT 146.560 114.720 146.900 115.550 ;
        RECT 148.380 115.040 148.730 116.290 ;
        RECT 152.080 114.720 152.420 115.550 ;
        RECT 153.900 115.040 154.250 116.290 ;
        RECT 156.935 115.635 158.145 116.725 ;
        RECT 156.935 115.095 157.455 115.635 ;
        RECT 157.625 114.925 158.145 115.465 ;
        RECT 144.975 114.175 150.320 114.720 ;
        RECT 150.495 114.175 155.840 114.720 ;
        RECT 156.935 114.175 158.145 114.925 ;
        RECT 2.750 114.005 158.230 114.175 ;
        RECT 110.050 82.390 111.700 82.560 ;
        RECT 106.050 55.390 107.700 55.560 ;
        RECT 106.050 13.810 106.220 55.390 ;
        RECT 106.700 52.750 107.050 54.910 ;
        RECT 105.360 12.870 106.300 13.810 ;
        RECT 106.050 10.110 106.220 12.870 ;
        RECT 106.700 10.590 107.050 12.750 ;
        RECT 107.530 10.110 107.700 55.390 ;
        RECT 110.050 37.110 110.220 82.390 ;
        RECT 110.700 79.750 111.050 81.910 ;
        RECT 110.700 37.590 111.050 39.750 ;
        RECT 111.530 37.110 111.700 82.390 ;
        RECT 110.050 36.940 111.700 37.110 ;
        RECT 113.050 82.390 114.700 82.560 ;
        RECT 113.050 37.110 113.220 82.390 ;
        RECT 113.700 79.750 114.050 81.910 ;
        RECT 113.700 37.590 114.050 39.750 ;
        RECT 114.530 37.110 114.700 82.390 ;
        RECT 113.050 36.940 114.700 37.110 ;
        RECT 116.050 82.390 117.700 82.560 ;
        RECT 116.050 37.110 116.220 82.390 ;
        RECT 116.700 79.750 117.050 81.910 ;
        RECT 116.700 37.590 117.050 39.750 ;
        RECT 117.530 37.110 117.700 82.390 ;
        RECT 116.050 36.940 117.700 37.110 ;
        RECT 119.050 82.390 120.700 82.560 ;
        RECT 119.050 37.110 119.220 82.390 ;
        RECT 119.700 79.750 120.050 81.910 ;
        RECT 119.700 37.590 120.050 39.750 ;
        RECT 120.530 37.110 120.700 82.390 ;
        RECT 119.050 36.940 120.700 37.110 ;
        RECT 122.050 82.390 123.700 82.560 ;
        RECT 122.050 37.110 122.220 82.390 ;
        RECT 122.700 79.750 123.050 81.910 ;
        RECT 122.700 37.590 123.050 39.750 ;
        RECT 123.530 37.110 123.700 82.390 ;
        RECT 122.050 36.940 123.700 37.110 ;
        RECT 125.050 82.390 126.700 82.560 ;
        RECT 125.050 37.110 125.220 82.390 ;
        RECT 125.700 79.750 126.050 81.910 ;
        RECT 125.700 37.590 126.050 39.750 ;
        RECT 126.530 37.110 126.700 82.390 ;
        RECT 125.050 36.940 126.700 37.110 ;
        RECT 128.050 82.390 129.700 82.560 ;
        RECT 128.050 37.110 128.220 82.390 ;
        RECT 128.700 79.750 129.050 81.910 ;
        RECT 128.700 37.590 129.050 39.750 ;
        RECT 129.530 37.110 129.700 82.390 ;
        RECT 128.050 36.940 129.700 37.110 ;
        RECT 131.050 82.390 132.700 82.560 ;
        RECT 131.050 37.110 131.220 82.390 ;
        RECT 131.700 79.750 132.050 81.910 ;
        RECT 131.700 37.590 132.050 39.750 ;
        RECT 132.530 37.110 132.700 82.390 ;
        RECT 131.050 36.940 132.700 37.110 ;
        RECT 106.050 9.940 107.700 10.110 ;
        RECT 110.050 35.390 111.700 35.560 ;
        RECT 110.050 10.110 110.220 35.390 ;
        RECT 110.700 32.750 111.050 34.910 ;
        RECT 110.700 10.590 111.050 12.750 ;
        RECT 111.530 10.110 111.700 35.390 ;
        RECT 110.050 9.940 111.700 10.110 ;
        RECT 113.050 35.390 114.700 35.560 ;
        RECT 113.050 10.110 113.220 35.390 ;
        RECT 113.700 32.750 114.050 34.910 ;
        RECT 113.700 10.590 114.050 12.750 ;
        RECT 114.530 10.110 114.700 35.390 ;
        RECT 113.050 9.940 114.700 10.110 ;
        RECT 116.050 35.390 117.700 35.560 ;
        RECT 116.050 10.110 116.220 35.390 ;
        RECT 116.700 32.750 117.050 34.910 ;
        RECT 116.700 10.590 117.050 12.750 ;
        RECT 117.530 10.110 117.700 35.390 ;
        RECT 116.050 9.940 117.700 10.110 ;
        RECT 119.050 35.390 120.700 35.560 ;
        RECT 119.050 10.110 119.220 35.390 ;
        RECT 119.700 32.750 120.050 34.910 ;
        RECT 119.700 10.590 120.050 12.750 ;
        RECT 120.530 10.110 120.700 35.390 ;
        RECT 119.050 9.940 120.700 10.110 ;
        RECT 122.050 35.390 123.700 35.560 ;
        RECT 122.050 10.110 122.220 35.390 ;
        RECT 122.700 32.750 123.050 34.910 ;
        RECT 122.700 10.590 123.050 12.750 ;
        RECT 123.530 10.110 123.700 35.390 ;
        RECT 122.050 9.940 123.700 10.110 ;
        RECT 125.050 35.390 126.700 35.560 ;
        RECT 125.050 10.110 125.220 35.390 ;
        RECT 125.700 32.750 126.050 34.910 ;
        RECT 125.700 10.590 126.050 12.750 ;
        RECT 126.530 10.110 126.700 35.390 ;
        RECT 125.050 9.940 126.700 10.110 ;
        RECT 128.050 35.390 129.700 35.560 ;
        RECT 128.050 10.110 128.220 35.390 ;
        RECT 128.700 32.750 129.050 34.910 ;
        RECT 128.700 10.590 129.050 12.750 ;
        RECT 129.530 10.110 129.700 35.390 ;
        RECT 128.050 9.940 129.700 10.110 ;
      LAYER met1 ;
        RECT 25.360 221.430 25.680 221.490 ;
        RECT 75.960 221.430 76.280 221.490 ;
        RECT 122.880 221.430 123.200 221.490 ;
        RECT 134.380 221.430 134.700 221.490 ;
        RECT 151.860 221.430 152.180 221.490 ;
        RECT 25.360 221.290 51.810 221.430 ;
        RECT 25.360 221.230 25.680 221.290 ;
        RECT 51.670 221.150 51.810 221.290 ;
        RECT 75.960 221.290 152.180 221.430 ;
        RECT 75.960 221.230 76.280 221.290 ;
        RECT 122.880 221.230 123.200 221.290 ;
        RECT 134.380 221.230 134.700 221.290 ;
        RECT 151.860 221.230 152.180 221.290 ;
        RECT 20.300 221.090 20.620 221.150 ;
        RECT 50.660 221.090 50.980 221.150 ;
        RECT 20.300 220.950 50.980 221.090 ;
        RECT 20.300 220.890 20.620 220.950 ;
        RECT 50.660 220.890 50.980 220.950 ;
        RECT 51.580 220.890 51.900 221.150 ;
        RECT 17.540 220.750 17.860 220.810 ;
        RECT 79.180 220.750 79.500 220.810 ;
        RECT 17.540 220.610 79.500 220.750 ;
        RECT 17.540 220.550 17.860 220.610 ;
        RECT 79.180 220.550 79.500 220.610 ;
        RECT 126.560 220.750 126.880 220.810 ;
        RECT 154.160 220.750 154.480 220.810 ;
        RECT 126.560 220.610 154.480 220.750 ;
        RECT 126.560 220.550 126.880 220.610 ;
        RECT 154.160 220.550 154.480 220.610 ;
        RECT 2.750 219.930 158.230 220.410 ;
        RECT 31.800 219.530 32.120 219.790 ;
        RECT 35.020 219.530 35.340 219.790 ;
        RECT 44.220 219.730 44.540 219.790 ;
        RECT 51.135 219.730 51.425 219.775 ;
        RECT 40.630 219.590 43.530 219.730 ;
        RECT 10.195 219.390 10.485 219.435 ;
        RECT 12.955 219.390 13.245 219.435 ;
        RECT 14.785 219.390 15.075 219.435 ;
        RECT 10.195 219.250 15.075 219.390 ;
        RECT 10.195 219.205 10.485 219.250 ;
        RECT 12.955 219.205 13.245 219.250 ;
        RECT 14.785 219.205 15.075 219.250 ;
        RECT 18.885 219.390 19.175 219.435 ;
        RECT 20.775 219.390 21.065 219.435 ;
        RECT 23.895 219.390 24.185 219.435 ;
        RECT 18.885 219.250 24.185 219.390 ;
        RECT 18.885 219.205 19.175 219.250 ;
        RECT 20.775 219.205 21.065 219.250 ;
        RECT 23.895 219.205 24.185 219.250 ;
        RECT 24.900 219.390 25.220 219.450 ;
        RECT 31.890 219.390 32.030 219.530 ;
        RECT 40.630 219.390 40.770 219.590 ;
        RECT 24.900 219.250 28.350 219.390 ;
        RECT 31.890 219.250 40.770 219.390 ;
        RECT 24.900 219.190 25.220 219.250 ;
        RECT 6.500 218.850 6.820 219.110 ;
        RECT 18.015 219.050 18.305 219.095 ;
        RECT 27.660 219.050 27.980 219.110 ;
        RECT 28.210 219.095 28.350 219.250 ;
        RECT 41.015 219.205 41.305 219.435 ;
        RECT 18.015 218.910 27.980 219.050 ;
        RECT 18.015 218.865 18.305 218.910 ;
        RECT 27.660 218.850 27.980 218.910 ;
        RECT 28.135 218.865 28.425 219.095 ;
        RECT 31.340 219.050 31.660 219.110 ;
        RECT 31.815 219.050 32.105 219.095 ;
        RECT 37.795 219.050 38.085 219.095 ;
        RECT 31.340 218.910 38.085 219.050 ;
        RECT 31.340 218.850 31.660 218.910 ;
        RECT 31.815 218.865 32.105 218.910 ;
        RECT 37.795 218.865 38.085 218.910 ;
        RECT 10.175 218.710 10.465 218.755 ;
        RECT 10.175 218.570 12.710 218.710 ;
        RECT 10.175 218.525 10.465 218.570 ;
        RECT 8.355 218.370 8.645 218.415 ;
        RECT 11.100 218.370 11.420 218.430 ;
        RECT 12.495 218.415 12.710 218.570 ;
        RECT 13.400 218.510 13.720 218.770 ;
        RECT 15.255 218.525 15.545 218.755 ;
        RECT 11.575 218.370 11.865 218.415 ;
        RECT 8.355 218.230 11.865 218.370 ;
        RECT 8.355 218.185 8.645 218.230 ;
        RECT 11.100 218.170 11.420 218.230 ;
        RECT 11.575 218.185 11.865 218.230 ;
        RECT 12.495 218.370 12.785 218.415 ;
        RECT 14.335 218.370 14.625 218.415 ;
        RECT 12.495 218.230 14.625 218.370 ;
        RECT 15.330 218.370 15.470 218.525 ;
        RECT 17.540 218.510 17.860 218.770 ;
        RECT 18.480 218.710 18.770 218.755 ;
        RECT 20.315 218.710 20.605 218.755 ;
        RECT 23.895 218.710 24.185 218.755 ;
        RECT 18.480 218.570 24.185 218.710 ;
        RECT 18.480 218.525 18.770 218.570 ;
        RECT 20.315 218.525 20.605 218.570 ;
        RECT 23.895 218.525 24.185 218.570 ;
        RECT 18.000 218.370 18.320 218.430 ;
        RECT 15.330 218.230 18.320 218.370 ;
        RECT 12.495 218.185 12.785 218.230 ;
        RECT 14.335 218.185 14.625 218.230 ;
        RECT 18.000 218.170 18.320 218.230 ;
        RECT 19.380 218.170 19.700 218.430 ;
        RECT 24.975 218.415 25.265 218.730 ;
        RECT 33.180 218.510 33.500 218.770 ;
        RECT 39.175 218.710 39.465 218.755 ;
        RECT 35.110 218.570 39.465 218.710 ;
        RECT 41.090 218.710 41.230 219.205 ;
        RECT 43.390 219.050 43.530 219.590 ;
        RECT 44.220 219.590 51.425 219.730 ;
        RECT 44.220 219.530 44.540 219.590 ;
        RECT 51.135 219.545 51.425 219.590 ;
        RECT 62.620 219.530 62.940 219.790 ;
        RECT 69.060 219.530 69.380 219.790 ;
        RECT 70.455 219.730 70.745 219.775 ;
        RECT 71.835 219.730 72.125 219.775 ;
        RECT 70.455 219.590 72.125 219.730 ;
        RECT 70.455 219.545 70.745 219.590 ;
        RECT 71.835 219.545 72.125 219.590 ;
        RECT 82.860 219.530 83.180 219.790 ;
        RECT 102.180 219.730 102.500 219.790 ;
        RECT 103.115 219.730 103.405 219.775 ;
        RECT 103.560 219.730 103.880 219.790 ;
        RECT 84.790 219.590 102.870 219.730 ;
        RECT 43.775 219.390 44.065 219.435 ;
        RECT 61.700 219.390 62.020 219.450 ;
        RECT 43.775 219.250 49.510 219.390 ;
        RECT 43.775 219.205 44.065 219.250 ;
        RECT 45.140 219.050 45.460 219.110 ;
        RECT 43.390 218.910 45.460 219.050 ;
        RECT 45.140 218.850 45.460 218.910 ;
        RECT 46.995 218.865 47.285 219.095 ;
        RECT 47.455 219.050 47.745 219.095 ;
        RECT 48.820 219.050 49.140 219.110 ;
        RECT 47.455 218.910 49.140 219.050 ;
        RECT 49.370 219.050 49.510 219.250 ;
        RECT 55.350 219.250 62.020 219.390 ;
        RECT 55.350 219.050 55.490 219.250 ;
        RECT 61.700 219.190 62.020 219.250 ;
        RECT 67.695 219.390 67.985 219.435 ;
        RECT 68.140 219.390 68.460 219.450 ;
        RECT 67.695 219.250 68.460 219.390 ;
        RECT 69.150 219.390 69.290 219.530 ;
        RECT 74.135 219.390 74.425 219.435 ;
        RECT 84.790 219.390 84.930 219.590 ;
        RECT 102.180 219.530 102.500 219.590 ;
        RECT 69.150 219.250 74.425 219.390 ;
        RECT 67.695 219.205 67.985 219.250 ;
        RECT 68.140 219.190 68.460 219.250 ;
        RECT 74.135 219.205 74.425 219.250 ;
        RECT 82.720 219.250 84.930 219.390 ;
        RECT 49.370 218.910 55.490 219.050 ;
        RECT 55.735 219.050 56.025 219.095 ;
        RECT 65.840 219.050 66.160 219.110 ;
        RECT 69.520 219.050 69.840 219.110 ;
        RECT 82.720 219.050 82.860 219.250 ;
        RECT 85.175 219.205 85.465 219.435 ;
        RECT 94.835 219.390 95.125 219.435 ;
        RECT 101.260 219.390 101.580 219.450 ;
        RECT 94.835 219.250 101.580 219.390 ;
        RECT 102.730 219.390 102.870 219.590 ;
        RECT 103.115 219.590 103.880 219.730 ;
        RECT 103.115 219.545 103.405 219.590 ;
        RECT 103.560 219.530 103.880 219.590 ;
        RECT 110.000 219.730 110.320 219.790 ;
        RECT 133.475 219.730 133.765 219.775 ;
        RECT 110.000 219.590 133.765 219.730 ;
        RECT 110.000 219.530 110.320 219.590 ;
        RECT 133.475 219.545 133.765 219.590 ;
        RECT 142.200 219.730 142.520 219.790 ;
        RECT 149.115 219.730 149.405 219.775 ;
        RECT 142.200 219.590 149.405 219.730 ;
        RECT 142.200 219.530 142.520 219.590 ;
        RECT 149.115 219.545 149.405 219.590 ;
        RECT 107.240 219.390 107.560 219.450 ;
        RECT 102.730 219.250 107.560 219.390 ;
        RECT 94.835 219.205 95.125 219.250 ;
        RECT 55.735 218.910 66.160 219.050 ;
        RECT 47.455 218.865 47.745 218.910 ;
        RECT 45.615 218.710 45.905 218.755 ;
        RECT 41.090 218.570 45.905 218.710 ;
        RECT 47.070 218.710 47.210 218.865 ;
        RECT 48.820 218.850 49.140 218.910 ;
        RECT 55.735 218.865 56.025 218.910 ;
        RECT 65.840 218.850 66.160 218.910 ;
        RECT 66.390 218.910 69.290 219.050 ;
        RECT 48.360 218.710 48.680 218.770 ;
        RECT 52.500 218.710 52.820 218.770 ;
        RECT 62.175 218.710 62.465 218.755 ;
        RECT 47.070 218.570 48.680 218.710 ;
        RECT 35.110 218.430 35.250 218.570 ;
        RECT 39.175 218.525 39.465 218.570 ;
        RECT 45.615 218.525 45.905 218.570 ;
        RECT 48.360 218.510 48.680 218.570 ;
        RECT 49.370 218.570 51.350 218.710 ;
        RECT 21.675 218.370 22.325 218.415 ;
        RECT 24.975 218.370 25.565 218.415 ;
        RECT 34.560 218.370 34.880 218.430 ;
        RECT 21.675 218.230 34.880 218.370 ;
        RECT 21.675 218.185 22.325 218.230 ;
        RECT 25.275 218.185 25.565 218.230 ;
        RECT 34.560 218.170 34.880 218.230 ;
        RECT 35.020 218.170 35.340 218.430 ;
        RECT 36.400 218.170 36.720 218.430 ;
        RECT 36.860 218.370 37.180 218.430 ;
        RECT 42.395 218.370 42.685 218.415 ;
        RECT 49.370 218.370 49.510 218.570 ;
        RECT 36.860 218.230 42.685 218.370 ;
        RECT 36.860 218.170 37.180 218.230 ;
        RECT 42.395 218.185 42.685 218.230 ;
        RECT 44.310 218.230 49.510 218.370 ;
        RECT 14.780 218.030 15.100 218.090 ;
        RECT 16.635 218.030 16.925 218.075 ;
        RECT 18.920 218.030 19.240 218.090 ;
        RECT 14.780 217.890 19.240 218.030 ;
        RECT 14.780 217.830 15.100 217.890 ;
        RECT 16.635 217.845 16.925 217.890 ;
        RECT 18.920 217.830 19.240 217.890 ;
        RECT 23.060 218.030 23.380 218.090 ;
        RECT 29.055 218.030 29.345 218.075 ;
        RECT 23.060 217.890 29.345 218.030 ;
        RECT 23.060 217.830 23.380 217.890 ;
        RECT 29.055 217.845 29.345 217.890 ;
        RECT 30.880 217.830 31.200 218.090 ;
        RECT 31.355 218.030 31.645 218.075 ;
        RECT 31.800 218.030 32.120 218.090 ;
        RECT 31.355 217.890 32.120 218.030 ;
        RECT 31.355 217.845 31.645 217.890 ;
        RECT 31.800 217.830 32.120 217.890 ;
        RECT 34.115 218.030 34.405 218.075 ;
        RECT 35.940 218.030 36.260 218.090 ;
        RECT 34.115 217.890 36.260 218.030 ;
        RECT 34.115 217.845 34.405 217.890 ;
        RECT 35.940 217.830 36.260 217.890 ;
        RECT 38.715 218.030 39.005 218.075 ;
        RECT 44.310 218.030 44.450 218.230 ;
        RECT 50.675 218.185 50.965 218.415 ;
        RECT 51.210 218.370 51.350 218.570 ;
        RECT 52.500 218.570 62.465 218.710 ;
        RECT 52.500 218.510 52.820 218.570 ;
        RECT 62.175 218.525 62.465 218.570 ;
        RECT 64.475 218.710 64.765 218.755 ;
        RECT 66.390 218.710 66.530 218.910 ;
        RECT 64.475 218.570 66.530 218.710 ;
        RECT 67.680 218.710 68.000 218.770 ;
        RECT 68.615 218.720 68.905 218.755 ;
        RECT 68.230 218.710 68.905 218.720 ;
        RECT 67.680 218.580 68.905 218.710 ;
        RECT 67.680 218.570 68.370 218.580 ;
        RECT 64.475 218.525 64.765 218.570 ;
        RECT 67.680 218.510 68.000 218.570 ;
        RECT 68.615 218.525 68.905 218.580 ;
        RECT 69.150 218.710 69.290 218.910 ;
        RECT 69.520 218.910 82.860 219.050 ;
        RECT 85.250 219.050 85.390 219.205 ;
        RECT 101.260 219.190 101.580 219.250 ;
        RECT 107.240 219.190 107.560 219.250 ;
        RECT 107.715 219.390 108.005 219.435 ;
        RECT 122.435 219.390 122.725 219.435 ;
        RECT 107.715 219.250 122.725 219.390 ;
        RECT 107.715 219.205 108.005 219.250 ;
        RECT 122.435 219.205 122.725 219.250 ;
        RECT 127.495 219.390 127.785 219.435 ;
        RECT 132.095 219.390 132.385 219.435 ;
        RECT 127.495 219.250 132.385 219.390 ;
        RECT 127.495 219.205 127.785 219.250 ;
        RECT 132.095 219.205 132.385 219.250 ;
        RECT 134.395 219.390 134.685 219.435 ;
        RECT 137.615 219.390 137.905 219.435 ;
        RECT 147.735 219.390 148.025 219.435 ;
        RECT 134.395 219.250 137.905 219.390 ;
        RECT 134.395 219.205 134.685 219.250 ;
        RECT 137.615 219.205 137.905 219.250 ;
        RECT 138.150 219.250 148.025 219.390 ;
        RECT 129.320 219.050 129.640 219.110 ;
        RECT 85.250 218.910 120.350 219.050 ;
        RECT 69.520 218.850 69.840 218.910 ;
        RECT 73.215 218.710 73.505 218.755 ;
        RECT 69.150 218.570 73.505 218.710 ;
        RECT 73.215 218.525 73.505 218.570 ;
        RECT 76.420 218.710 76.740 218.770 ;
        RECT 82.415 218.710 82.705 218.755 ;
        RECT 76.420 218.570 82.705 218.710 ;
        RECT 76.420 218.510 76.740 218.570 ;
        RECT 82.415 218.525 82.705 218.570 ;
        RECT 84.255 218.710 84.545 218.755 ;
        RECT 93.455 218.710 93.745 218.755 ;
        RECT 84.255 218.570 93.745 218.710 ;
        RECT 84.255 218.525 84.545 218.570 ;
        RECT 93.455 218.525 93.745 218.570 ;
        RECT 94.375 218.525 94.665 218.755 ;
        RECT 56.180 218.370 56.500 218.430 ;
        RECT 51.210 218.230 56.500 218.370 ;
        RECT 38.715 217.890 44.450 218.030 ;
        RECT 38.715 217.845 39.005 217.890 ;
        RECT 44.680 217.830 45.000 218.090 ;
        RECT 45.600 218.030 45.920 218.090 ;
        RECT 47.915 218.030 48.205 218.075 ;
        RECT 45.600 217.890 48.205 218.030 ;
        RECT 45.600 217.830 45.920 217.890 ;
        RECT 47.915 217.845 48.205 217.890 ;
        RECT 49.755 218.030 50.045 218.075 ;
        RECT 50.750 218.030 50.890 218.185 ;
        RECT 56.180 218.170 56.500 218.230 ;
        RECT 56.640 218.370 56.960 218.430 ;
        RECT 57.115 218.370 57.405 218.415 ;
        RECT 56.640 218.230 57.405 218.370 ;
        RECT 56.640 218.170 56.960 218.230 ;
        RECT 57.115 218.185 57.405 218.230 ;
        RECT 58.480 218.370 58.800 218.430 ;
        RECT 59.415 218.370 59.705 218.415 ;
        RECT 58.480 218.230 59.705 218.370 ;
        RECT 58.480 218.170 58.800 218.230 ;
        RECT 59.415 218.185 59.705 218.230 ;
        RECT 61.700 218.170 62.020 218.430 ;
        RECT 64.920 218.370 65.240 218.430 ;
        RECT 65.395 218.370 65.685 218.415 ;
        RECT 64.920 218.230 65.685 218.370 ;
        RECT 64.920 218.170 65.240 218.230 ;
        RECT 65.395 218.185 65.685 218.230 ;
        RECT 66.300 218.170 66.620 218.430 ;
        RECT 72.740 218.370 73.060 218.430 ;
        RECT 75.500 218.370 75.820 218.430 ;
        RECT 70.990 218.230 72.510 218.370 ;
        RECT 49.755 217.890 50.890 218.030 ;
        RECT 60.795 218.030 61.085 218.075 ;
        RECT 61.240 218.030 61.560 218.090 ;
        RECT 60.795 217.890 61.560 218.030 ;
        RECT 61.790 218.030 61.930 218.170 ;
        RECT 70.990 218.090 71.130 218.230 ;
        RECT 66.760 218.030 67.080 218.090 ;
        RECT 69.075 218.030 69.365 218.075 ;
        RECT 61.790 217.890 69.365 218.030 ;
        RECT 49.755 217.845 50.045 217.890 ;
        RECT 60.795 217.845 61.085 217.890 ;
        RECT 61.240 217.830 61.560 217.890 ;
        RECT 66.760 217.830 67.080 217.890 ;
        RECT 69.075 217.845 69.365 217.890 ;
        RECT 69.520 217.830 69.840 218.090 ;
        RECT 70.900 217.830 71.220 218.090 ;
        RECT 71.820 218.075 72.140 218.090 ;
        RECT 71.755 217.845 72.140 218.075 ;
        RECT 72.370 218.030 72.510 218.230 ;
        RECT 72.740 218.230 75.820 218.370 ;
        RECT 72.740 218.170 73.060 218.230 ;
        RECT 75.500 218.170 75.820 218.230 ;
        RECT 83.320 218.030 83.640 218.090 ;
        RECT 72.370 217.890 83.640 218.030 ;
        RECT 94.450 218.030 94.590 218.525 ;
        RECT 95.280 218.510 95.600 218.770 ;
        RECT 95.740 218.510 96.060 218.770 ;
        RECT 96.675 218.525 96.965 218.755 ;
        RECT 97.580 218.710 97.900 218.770 ;
        RECT 102.195 218.710 102.485 218.755 ;
        RECT 97.580 218.570 102.485 218.710 ;
        RECT 96.750 218.370 96.890 218.525 ;
        RECT 97.580 218.510 97.900 218.570 ;
        RECT 102.195 218.525 102.485 218.570 ;
        RECT 102.640 218.710 102.960 218.770 ;
        RECT 103.115 218.710 103.405 218.755 ;
        RECT 102.640 218.570 103.405 218.710 ;
        RECT 102.640 218.510 102.960 218.570 ;
        RECT 103.115 218.525 103.405 218.570 ;
        RECT 107.240 218.710 107.560 218.770 ;
        RECT 109.095 218.710 109.385 218.755 ;
        RECT 119.660 218.710 119.980 218.770 ;
        RECT 120.210 218.755 120.350 218.910 ;
        RECT 121.130 218.910 129.640 219.050 ;
        RECT 107.240 218.570 119.980 218.710 ;
        RECT 107.240 218.510 107.560 218.570 ;
        RECT 109.095 218.525 109.385 218.570 ;
        RECT 119.660 218.510 119.980 218.570 ;
        RECT 120.135 218.525 120.425 218.755 ;
        RECT 104.940 218.370 105.260 218.430 ;
        RECT 121.130 218.370 121.270 218.910 ;
        RECT 129.320 218.850 129.640 218.910 ;
        RECT 123.340 218.510 123.660 218.770 ;
        RECT 124.260 218.710 124.580 218.770 ;
        RECT 128.875 218.710 129.165 218.755 ;
        RECT 124.260 218.570 129.165 218.710 ;
        RECT 124.260 218.510 124.580 218.570 ;
        RECT 128.875 218.525 129.165 218.570 ;
        RECT 130.240 218.510 130.560 218.770 ;
        RECT 133.000 218.510 133.320 218.770 ;
        RECT 137.140 218.510 137.460 218.770 ;
        RECT 137.600 218.710 137.920 218.770 ;
        RECT 138.150 218.710 138.290 219.250 ;
        RECT 147.735 219.205 148.025 219.250 ;
        RECT 144.040 219.050 144.360 219.110 ;
        RECT 146.355 219.050 146.645 219.095 ;
        RECT 144.040 218.910 146.645 219.050 ;
        RECT 144.040 218.850 144.360 218.910 ;
        RECT 146.355 218.865 146.645 218.910 ;
        RECT 137.600 218.570 138.290 218.710 ;
        RECT 137.600 218.510 137.920 218.570 ;
        RECT 138.520 218.510 138.840 218.770 ;
        RECT 140.360 218.510 140.680 218.770 ;
        RECT 144.960 218.510 145.280 218.770 ;
        RECT 145.880 218.755 146.200 218.770 ;
        RECT 145.665 218.525 146.200 218.755 ;
        RECT 147.275 218.525 147.565 218.755 ;
        RECT 145.880 218.510 146.200 218.525 ;
        RECT 96.750 218.230 105.260 218.370 ;
        RECT 104.940 218.170 105.260 218.230 ;
        RECT 119.750 218.230 121.270 218.370 ;
        RECT 121.975 218.370 122.265 218.415 ;
        RECT 131.620 218.370 131.940 218.430 ;
        RECT 135.775 218.370 136.065 218.415 ;
        RECT 147.350 218.370 147.490 218.525 ;
        RECT 148.640 218.510 148.960 218.770 ;
        RECT 150.020 218.510 150.340 218.770 ;
        RECT 151.400 218.710 151.720 218.770 ;
        RECT 152.335 218.710 152.625 218.755 ;
        RECT 151.400 218.570 152.625 218.710 ;
        RECT 151.400 218.510 151.720 218.570 ;
        RECT 152.335 218.525 152.625 218.570 ;
        RECT 148.180 218.370 148.500 218.430 ;
        RECT 121.975 218.230 126.790 218.370 ;
        RECT 98.040 218.030 98.360 218.090 ;
        RECT 94.450 217.890 98.360 218.030 ;
        RECT 71.820 217.830 72.140 217.845 ;
        RECT 83.320 217.830 83.640 217.890 ;
        RECT 98.040 217.830 98.360 217.890 ;
        RECT 103.100 218.030 103.420 218.090 ;
        RECT 119.750 218.075 119.890 218.230 ;
        RECT 121.975 218.185 122.265 218.230 ;
        RECT 106.795 218.030 107.085 218.075 ;
        RECT 103.100 217.890 107.085 218.030 ;
        RECT 103.100 217.830 103.420 217.890 ;
        RECT 106.795 217.845 107.085 217.890 ;
        RECT 119.675 217.845 119.965 218.075 ;
        RECT 120.580 217.830 120.900 218.090 ;
        RECT 121.040 218.030 121.360 218.090 ;
        RECT 124.260 218.030 124.580 218.090 ;
        RECT 126.650 218.075 126.790 218.230 ;
        RECT 131.620 218.230 148.500 218.370 ;
        RECT 131.620 218.170 131.940 218.230 ;
        RECT 135.775 218.185 136.065 218.230 ;
        RECT 148.180 218.170 148.500 218.230 ;
        RECT 121.040 217.890 124.580 218.030 ;
        RECT 121.040 217.830 121.360 217.890 ;
        RECT 124.260 217.830 124.580 217.890 ;
        RECT 126.575 217.845 126.865 218.075 ;
        RECT 129.320 217.830 129.640 218.090 ;
        RECT 136.220 217.830 136.540 218.090 ;
        RECT 141.295 218.030 141.585 218.075 ;
        RECT 144.960 218.030 145.280 218.090 ;
        RECT 141.295 217.890 145.280 218.030 ;
        RECT 141.295 217.845 141.585 217.890 ;
        RECT 144.960 217.830 145.280 217.890 ;
        RECT 146.800 217.830 147.120 218.090 ;
        RECT 151.400 217.830 151.720 218.090 ;
        RECT 2.750 217.210 159.030 217.690 ;
        RECT 10.640 217.010 10.960 217.070 ;
        RECT 17.555 217.010 17.845 217.055 ;
        RECT 19.380 217.010 19.700 217.070 ;
        RECT 10.640 216.870 12.250 217.010 ;
        RECT 10.640 216.810 10.960 216.870 ;
        RECT 7.875 216.670 8.525 216.715 ;
        RECT 11.475 216.670 11.765 216.715 ;
        RECT 7.875 216.530 11.765 216.670 ;
        RECT 12.110 216.670 12.250 216.870 ;
        RECT 17.555 216.870 19.700 217.010 ;
        RECT 17.555 216.825 17.845 216.870 ;
        RECT 19.380 216.810 19.700 216.870 ;
        RECT 19.840 216.810 20.160 217.070 ;
        RECT 20.300 216.810 20.620 217.070 ;
        RECT 23.075 216.825 23.365 217.055 ;
        RECT 14.335 216.670 14.625 216.715 ;
        RECT 23.150 216.670 23.290 216.825 ;
        RECT 24.900 216.810 25.220 217.070 ;
        RECT 25.360 216.810 25.680 217.070 ;
        RECT 32.260 216.810 32.580 217.070 ;
        RECT 33.180 217.010 33.500 217.070 ;
        RECT 34.115 217.010 34.405 217.055 ;
        RECT 44.680 217.010 45.000 217.070 ;
        RECT 33.180 216.870 34.405 217.010 ;
        RECT 33.180 216.810 33.500 216.870 ;
        RECT 34.115 216.825 34.405 216.870 ;
        RECT 43.850 216.870 45.000 217.010 ;
        RECT 12.110 216.530 14.625 216.670 ;
        RECT 7.875 216.485 8.525 216.530 ;
        RECT 11.175 216.485 11.765 216.530 ;
        RECT 14.335 216.485 14.625 216.530 ;
        RECT 16.710 216.530 23.290 216.670 ;
        RECT 23.520 216.670 23.840 216.730 ;
        RECT 35.020 216.670 35.340 216.730 ;
        RECT 43.850 216.715 43.990 216.870 ;
        RECT 44.680 216.810 45.000 216.870 ;
        RECT 45.140 216.810 45.460 217.070 ;
        RECT 46.980 217.010 47.300 217.070 ;
        RECT 50.215 217.010 50.505 217.055 ;
        RECT 65.380 217.010 65.700 217.070 ;
        RECT 46.980 216.870 50.505 217.010 ;
        RECT 46.980 216.810 47.300 216.870 ;
        RECT 50.215 216.825 50.505 216.870 ;
        RECT 55.350 216.870 65.700 217.010 ;
        RECT 23.520 216.530 35.340 216.670 ;
        RECT 11.175 216.390 11.465 216.485 ;
        RECT 4.680 216.330 4.970 216.375 ;
        RECT 6.515 216.330 6.805 216.375 ;
        RECT 10.095 216.330 10.385 216.375 ;
        RECT 4.680 216.190 10.385 216.330 ;
        RECT 4.680 216.145 4.970 216.190 ;
        RECT 6.515 216.145 6.805 216.190 ;
        RECT 10.095 216.145 10.385 216.190 ;
        RECT 11.100 216.170 11.465 216.390 ;
        RECT 16.710 216.375 16.850 216.530 ;
        RECT 23.520 216.470 23.840 216.530 ;
        RECT 35.020 216.470 35.340 216.530 ;
        RECT 37.895 216.670 38.185 216.715 ;
        RECT 41.135 216.670 41.785 216.715 ;
        RECT 37.895 216.530 41.785 216.670 ;
        RECT 37.895 216.485 38.485 216.530 ;
        RECT 41.135 216.485 41.785 216.530 ;
        RECT 43.775 216.485 44.065 216.715 ;
        RECT 45.230 216.670 45.370 216.810 ;
        RECT 47.915 216.670 48.205 216.715 ;
        RECT 45.230 216.530 48.205 216.670 ;
        RECT 47.915 216.485 48.205 216.530 ;
        RECT 48.375 216.670 48.665 216.715 ;
        RECT 55.350 216.670 55.490 216.870 ;
        RECT 65.380 216.810 65.700 216.870 ;
        RECT 65.840 217.010 66.160 217.070 ;
        RECT 68.600 217.055 68.920 217.070 ;
        RECT 68.600 217.010 68.985 217.055 ;
        RECT 65.840 216.870 68.985 217.010 ;
        RECT 65.840 216.810 66.160 216.870 ;
        RECT 68.600 216.825 68.985 216.870 ;
        RECT 69.535 217.010 69.825 217.055 ;
        RECT 71.820 217.010 72.140 217.070 ;
        RECT 69.535 216.870 72.140 217.010 ;
        RECT 69.535 216.825 69.825 216.870 ;
        RECT 68.600 216.810 68.920 216.825 ;
        RECT 71.820 216.810 72.140 216.870 ;
        RECT 78.720 216.810 79.040 217.070 ;
        RECT 79.270 216.870 89.990 217.010 ;
        RECT 61.240 216.670 61.560 216.730 ;
        RECT 67.695 216.670 67.985 216.715 ;
        RECT 73.660 216.670 73.980 216.730 ;
        RECT 79.270 216.670 79.410 216.870 ;
        RECT 89.850 216.730 89.990 216.870 ;
        RECT 92.520 216.810 92.840 217.070 ;
        RECT 95.280 216.810 95.600 217.070 ;
        RECT 96.200 217.055 96.520 217.070 ;
        RECT 96.135 216.825 96.520 217.055 ;
        RECT 102.640 217.010 102.960 217.070 ;
        RECT 96.200 216.810 96.520 216.825 ;
        RECT 96.750 216.870 102.960 217.010 ;
        RECT 48.375 216.530 55.490 216.670 ;
        RECT 55.810 216.530 57.330 216.670 ;
        RECT 48.375 216.485 48.665 216.530 ;
        RECT 11.100 216.130 11.420 216.170 ;
        RECT 15.255 216.145 15.545 216.375 ;
        RECT 16.635 216.145 16.925 216.375 ;
        RECT 19.010 216.190 26.050 216.330 ;
        RECT 4.215 215.990 4.505 216.035 ;
        RECT 5.595 215.990 5.885 216.035 ;
        RECT 6.040 215.990 6.360 216.050 ;
        RECT 4.215 215.850 4.890 215.990 ;
        RECT 4.215 215.805 4.505 215.850 ;
        RECT 4.750 215.370 4.890 215.850 ;
        RECT 5.595 215.850 6.360 215.990 ;
        RECT 15.330 215.990 15.470 216.145 ;
        RECT 19.010 216.050 19.150 216.190 ;
        RECT 15.330 215.850 18.230 215.990 ;
        RECT 5.595 215.805 5.885 215.850 ;
        RECT 6.040 215.790 6.360 215.850 ;
        RECT 18.090 215.695 18.230 215.850 ;
        RECT 18.920 215.790 19.240 216.050 ;
        RECT 20.850 216.035 20.990 216.190 ;
        RECT 25.910 216.035 26.050 216.190 ;
        RECT 27.200 216.130 27.520 216.390 ;
        RECT 29.040 216.130 29.360 216.390 ;
        RECT 31.815 216.145 32.105 216.375 ;
        RECT 34.560 216.330 34.880 216.390 ;
        RECT 38.195 216.330 38.485 216.485 ;
        RECT 34.560 216.190 38.485 216.330 ;
        RECT 20.775 215.805 21.065 216.035 ;
        RECT 25.835 215.990 26.125 216.035 ;
        RECT 30.895 215.990 31.185 216.035 ;
        RECT 31.340 215.990 31.660 216.050 ;
        RECT 25.835 215.850 31.660 215.990 ;
        RECT 25.835 215.805 26.125 215.850 ;
        RECT 30.895 215.805 31.185 215.850 ;
        RECT 31.340 215.790 31.660 215.850 ;
        RECT 5.085 215.650 5.375 215.695 ;
        RECT 6.975 215.650 7.265 215.695 ;
        RECT 10.095 215.650 10.385 215.695 ;
        RECT 5.085 215.510 10.385 215.650 ;
        RECT 5.085 215.465 5.375 215.510 ;
        RECT 6.975 215.465 7.265 215.510 ;
        RECT 10.095 215.465 10.385 215.510 ;
        RECT 18.015 215.465 18.305 215.695 ;
        RECT 4.660 215.110 4.980 215.370 ;
        RECT 16.160 215.110 16.480 215.370 ;
        RECT 28.120 215.110 28.440 215.370 ;
        RECT 29.975 215.310 30.265 215.355 ;
        RECT 30.420 215.310 30.740 215.370 ;
        RECT 29.975 215.170 30.740 215.310 ;
        RECT 31.890 215.310 32.030 216.145 ;
        RECT 34.560 216.130 34.880 216.190 ;
        RECT 38.195 216.170 38.485 216.190 ;
        RECT 39.275 216.330 39.565 216.375 ;
        RECT 42.855 216.330 43.145 216.375 ;
        RECT 44.690 216.330 44.980 216.375 ;
        RECT 39.275 216.190 44.980 216.330 ;
        RECT 39.275 216.145 39.565 216.190 ;
        RECT 42.855 216.145 43.145 216.190 ;
        RECT 44.690 216.145 44.980 216.190 ;
        RECT 51.580 216.330 51.900 216.390 ;
        RECT 52.055 216.330 52.345 216.375 ;
        RECT 51.580 216.190 52.345 216.330 ;
        RECT 51.580 216.130 51.900 216.190 ;
        RECT 52.055 216.145 52.345 216.190 ;
        RECT 52.515 216.330 52.805 216.375 ;
        RECT 52.960 216.330 53.280 216.390 ;
        RECT 52.515 216.190 53.280 216.330 ;
        RECT 52.515 216.145 52.805 216.190 ;
        RECT 52.960 216.130 53.280 216.190 ;
        RECT 53.880 216.330 54.200 216.390 ;
        RECT 55.810 216.330 55.950 216.530 ;
        RECT 53.880 216.190 55.950 216.330 ;
        RECT 56.180 216.330 56.500 216.390 ;
        RECT 56.655 216.330 56.945 216.375 ;
        RECT 56.180 216.190 56.945 216.330 ;
        RECT 57.190 216.330 57.330 216.530 ;
        RECT 61.240 216.530 73.980 216.670 ;
        RECT 61.240 216.470 61.560 216.530 ;
        RECT 67.695 216.485 67.985 216.530 ;
        RECT 73.660 216.470 73.980 216.530 ;
        RECT 78.120 216.530 79.410 216.670 ;
        RECT 80.100 216.670 80.420 216.730 ;
        RECT 81.955 216.670 82.245 216.715 ;
        RECT 80.100 216.530 83.090 216.670 ;
        RECT 78.120 216.390 78.260 216.530 ;
        RECT 80.100 216.470 80.420 216.530 ;
        RECT 81.955 216.485 82.245 216.530 ;
        RECT 61.700 216.330 62.020 216.390 ;
        RECT 62.175 216.330 62.465 216.375 ;
        RECT 57.190 216.190 62.465 216.330 ;
        RECT 53.880 216.130 54.200 216.190 ;
        RECT 56.180 216.130 56.500 216.190 ;
        RECT 56.655 216.145 56.945 216.190 ;
        RECT 61.700 216.130 62.020 216.190 ;
        RECT 62.175 216.145 62.465 216.190 ;
        RECT 62.635 216.330 62.925 216.375 ;
        RECT 64.000 216.330 64.320 216.390 ;
        RECT 62.635 216.190 64.320 216.330 ;
        RECT 62.635 216.145 62.925 216.190 ;
        RECT 64.000 216.130 64.320 216.190 ;
        RECT 66.300 216.130 66.620 216.390 ;
        RECT 69.520 216.130 69.840 216.390 ;
        RECT 70.440 216.330 70.760 216.390 ;
        RECT 70.915 216.330 71.205 216.375 ;
        RECT 70.440 216.190 71.205 216.330 ;
        RECT 70.440 216.130 70.760 216.190 ;
        RECT 70.915 216.145 71.205 216.190 ;
        RECT 73.200 216.330 73.520 216.390 ;
        RECT 75.515 216.330 75.805 216.375 ;
        RECT 73.200 216.190 75.805 216.330 ;
        RECT 73.200 216.130 73.520 216.190 ;
        RECT 75.515 216.145 75.805 216.190 ;
        RECT 75.960 216.330 76.280 216.390 ;
        RECT 75.960 216.190 76.475 216.330 ;
        RECT 75.960 216.130 76.280 216.190 ;
        RECT 76.880 216.130 77.200 216.390 ;
        RECT 78.120 216.375 78.580 216.390 ;
        RECT 77.355 216.145 77.645 216.375 ;
        RECT 78.045 216.145 78.580 216.375 ;
        RECT 36.400 215.990 36.720 216.050 ;
        RECT 36.400 215.850 44.910 215.990 ;
        RECT 36.400 215.790 36.720 215.850 ;
        RECT 39.275 215.650 39.565 215.695 ;
        RECT 42.395 215.650 42.685 215.695 ;
        RECT 44.285 215.650 44.575 215.695 ;
        RECT 39.275 215.510 44.575 215.650 ;
        RECT 44.770 215.650 44.910 215.850 ;
        RECT 45.140 215.790 45.460 216.050 ;
        RECT 48.360 215.990 48.680 216.050 ;
        RECT 49.295 215.990 49.585 216.035 ;
        RECT 49.740 215.990 50.060 216.050 ;
        RECT 53.435 215.990 53.725 216.035 ;
        RECT 48.360 215.850 55.030 215.990 ;
        RECT 48.360 215.790 48.680 215.850 ;
        RECT 49.295 215.805 49.585 215.850 ;
        RECT 49.740 215.790 50.060 215.850 ;
        RECT 53.435 215.805 53.725 215.850 ;
        RECT 46.075 215.650 46.365 215.695 ;
        RECT 44.770 215.510 46.365 215.650 ;
        RECT 39.275 215.465 39.565 215.510 ;
        RECT 42.395 215.465 42.685 215.510 ;
        RECT 44.285 215.465 44.575 215.510 ;
        RECT 46.075 215.465 46.365 215.510 ;
        RECT 48.820 215.650 49.140 215.710 ;
        RECT 54.340 215.650 54.660 215.710 ;
        RECT 48.820 215.510 54.660 215.650 ;
        RECT 54.890 215.650 55.030 215.850 ;
        RECT 57.100 215.790 57.420 216.050 ;
        RECT 57.560 215.990 57.880 216.050 ;
        RECT 63.095 215.990 63.385 216.035 ;
        RECT 57.560 215.850 63.385 215.990 ;
        RECT 57.560 215.790 57.880 215.850 ;
        RECT 63.095 215.805 63.385 215.850 ;
        RECT 65.380 215.990 65.700 216.050 ;
        RECT 69.060 215.990 69.380 216.050 ;
        RECT 65.380 215.850 69.380 215.990 ;
        RECT 69.610 215.990 69.750 216.130 ;
        RECT 72.295 215.990 72.585 216.035 ;
        RECT 69.610 215.850 72.585 215.990 ;
        RECT 65.380 215.790 65.700 215.850 ;
        RECT 69.060 215.790 69.380 215.850 ;
        RECT 72.295 215.805 72.585 215.850 ;
        RECT 77.430 215.990 77.570 216.145 ;
        RECT 78.260 216.130 78.580 216.145 ;
        RECT 79.180 216.330 79.500 216.390 ;
        RECT 80.575 216.330 80.865 216.375 ;
        RECT 79.180 216.190 80.865 216.330 ;
        RECT 79.180 216.130 79.500 216.190 ;
        RECT 80.575 216.145 80.865 216.190 ;
        RECT 81.480 216.130 81.800 216.390 ;
        RECT 82.400 216.130 82.720 216.390 ;
        RECT 82.950 216.330 83.090 216.530 ;
        RECT 83.320 216.470 83.640 216.730 ;
        RECT 89.760 216.670 90.080 216.730 ;
        RECT 96.750 216.670 96.890 216.870 ;
        RECT 102.640 216.810 102.960 216.870 ;
        RECT 107.715 217.010 108.005 217.055 ;
        RECT 111.840 217.010 112.160 217.070 ;
        RECT 120.580 217.010 120.900 217.070 ;
        RECT 121.515 217.010 121.805 217.055 ;
        RECT 134.380 217.010 134.700 217.070 ;
        RECT 107.715 216.870 111.610 217.010 ;
        RECT 107.715 216.825 108.005 216.870 ;
        RECT 89.760 216.530 96.890 216.670 ;
        RECT 97.120 216.670 97.440 216.730 ;
        RECT 107.240 216.670 107.560 216.730 ;
        RECT 111.470 216.670 111.610 216.870 ;
        RECT 111.840 216.870 120.365 217.010 ;
        RECT 111.840 216.810 112.160 216.870 ;
        RECT 112.300 216.670 112.620 216.730 ;
        RECT 119.200 216.670 119.520 216.730 ;
        RECT 97.120 216.530 104.250 216.670 ;
        RECT 89.760 216.470 90.080 216.530 ;
        RECT 97.120 216.470 97.440 216.530 ;
        RECT 91.140 216.330 91.460 216.390 ;
        RECT 82.950 216.190 91.460 216.330 ;
        RECT 91.140 216.130 91.460 216.190 ;
        RECT 91.600 216.130 91.920 216.390 ;
        RECT 93.605 216.330 93.895 216.375 ;
        RECT 93.530 216.145 93.895 216.330 ;
        RECT 100.815 216.145 101.105 216.375 ;
        RECT 81.940 215.990 82.260 216.050 ;
        RECT 91.690 215.990 91.830 216.130 ;
        RECT 77.430 215.850 91.830 215.990 ;
        RECT 57.650 215.650 57.790 215.790 ;
        RECT 54.890 215.510 57.790 215.650 ;
        RECT 59.860 215.650 60.180 215.710 ;
        RECT 77.430 215.650 77.570 215.850 ;
        RECT 81.940 215.790 82.260 215.850 ;
        RECT 59.860 215.510 77.570 215.650 ;
        RECT 48.820 215.450 49.140 215.510 ;
        RECT 54.340 215.450 54.660 215.510 ;
        RECT 59.860 215.450 60.180 215.510 ;
        RECT 53.880 215.310 54.200 215.370 ;
        RECT 31.890 215.170 54.200 215.310 ;
        RECT 29.975 215.125 30.265 215.170 ;
        RECT 30.420 215.110 30.740 215.170 ;
        RECT 53.880 215.110 54.200 215.170 ;
        RECT 54.800 215.110 55.120 215.370 ;
        RECT 58.020 215.310 58.340 215.370 ;
        RECT 60.335 215.310 60.625 215.355 ;
        RECT 58.020 215.170 60.625 215.310 ;
        RECT 58.020 215.110 58.340 215.170 ;
        RECT 60.335 215.125 60.625 215.170 ;
        RECT 61.930 215.310 62.250 215.370 ;
        RECT 64.935 215.310 65.225 215.355 ;
        RECT 61.930 215.170 65.225 215.310 ;
        RECT 61.930 215.110 62.250 215.170 ;
        RECT 64.935 215.125 65.225 215.170 ;
        RECT 68.600 215.110 68.920 215.370 ;
        RECT 86.540 215.310 86.860 215.370 ;
        RECT 93.530 215.310 93.670 216.145 ;
        RECT 94.360 215.790 94.680 216.050 ;
        RECT 94.835 215.990 95.125 216.035 ;
        RECT 95.280 215.990 95.600 216.050 ;
        RECT 94.835 215.850 95.600 215.990 ;
        RECT 94.835 215.805 95.125 215.850 ;
        RECT 95.280 215.790 95.600 215.850 ;
        RECT 96.660 215.650 96.980 215.710 ;
        RECT 100.890 215.650 101.030 216.145 ;
        RECT 101.260 216.130 101.580 216.390 ;
        RECT 101.735 216.280 102.025 216.375 ;
        RECT 103.560 216.330 103.880 216.390 ;
        RECT 103.190 216.280 103.880 216.330 ;
        RECT 101.735 216.190 103.880 216.280 ;
        RECT 104.110 216.330 104.250 216.530 ;
        RECT 107.240 216.530 109.770 216.670 ;
        RECT 111.470 216.530 112.620 216.670 ;
        RECT 107.240 216.470 107.560 216.530 ;
        RECT 108.175 216.330 108.465 216.375 ;
        RECT 109.080 216.330 109.400 216.390 ;
        RECT 104.110 216.190 109.400 216.330 ;
        RECT 109.630 216.330 109.770 216.530 ;
        RECT 112.300 216.470 112.620 216.530 ;
        RECT 112.850 216.530 119.520 216.670 ;
        RECT 120.225 216.670 120.365 216.870 ;
        RECT 120.580 216.870 121.805 217.010 ;
        RECT 120.580 216.810 120.900 216.870 ;
        RECT 121.515 216.825 121.805 216.870 ;
        RECT 125.730 216.870 134.150 217.010 ;
        RECT 125.730 216.670 125.870 216.870 ;
        RECT 120.225 216.530 125.870 216.670 ;
        RECT 126.190 216.530 133.690 216.670 ;
        RECT 112.850 216.375 112.990 216.530 ;
        RECT 119.200 216.470 119.520 216.530 ;
        RECT 112.775 216.330 113.065 216.375 ;
        RECT 109.630 216.190 113.065 216.330 ;
        RECT 101.735 216.145 103.330 216.190 ;
        RECT 101.810 216.140 103.330 216.145 ;
        RECT 103.560 216.130 103.880 216.190 ;
        RECT 108.175 216.145 108.465 216.190 ;
        RECT 109.080 216.130 109.400 216.190 ;
        RECT 112.775 216.145 113.065 216.190 ;
        RECT 113.695 216.145 113.985 216.375 ;
        RECT 103.650 215.990 103.790 216.130 ;
        RECT 111.840 215.990 112.160 216.050 ;
        RECT 103.650 215.850 112.160 215.990 ;
        RECT 113.770 215.990 113.910 216.145 ;
        RECT 114.140 216.130 114.460 216.390 ;
        RECT 114.600 216.130 114.920 216.390 ;
        RECT 116.440 216.130 116.760 216.390 ;
        RECT 116.900 216.330 117.220 216.390 ;
        RECT 117.375 216.330 117.665 216.375 ;
        RECT 116.900 216.190 117.665 216.330 ;
        RECT 116.900 216.130 117.220 216.190 ;
        RECT 117.375 216.145 117.665 216.190 ;
        RECT 117.820 216.130 118.140 216.390 ;
        RECT 122.420 216.130 122.740 216.390 ;
        RECT 122.895 216.330 123.185 216.375 ;
        RECT 124.735 216.330 125.025 216.375 ;
        RECT 122.895 216.190 125.025 216.330 ;
        RECT 122.895 216.145 123.185 216.190 ;
        RECT 124.735 216.145 125.025 216.190 ;
        RECT 125.640 216.130 125.960 216.390 ;
        RECT 118.280 215.990 118.600 216.050 ;
        RECT 123.355 215.990 123.645 216.035 ;
        RECT 113.770 215.850 118.600 215.990 ;
        RECT 111.840 215.790 112.160 215.850 ;
        RECT 118.280 215.790 118.600 215.850 ;
        RECT 118.830 215.850 123.645 215.990 ;
        RECT 109.095 215.650 109.385 215.695 ;
        RECT 96.660 215.510 109.385 215.650 ;
        RECT 96.660 215.450 96.980 215.510 ;
        RECT 109.095 215.465 109.385 215.510 ;
        RECT 109.540 215.650 109.860 215.710 ;
        RECT 118.830 215.695 118.970 215.850 ;
        RECT 123.355 215.805 123.645 215.850 ;
        RECT 123.815 215.990 124.105 216.035 ;
        RECT 126.190 215.990 126.330 216.530 ;
        RECT 133.550 216.390 133.690 216.530 ;
        RECT 126.560 216.130 126.880 216.390 ;
        RECT 127.020 216.130 127.340 216.390 ;
        RECT 127.480 216.130 127.800 216.390 ;
        RECT 128.400 216.130 128.720 216.390 ;
        RECT 128.860 216.130 129.180 216.390 ;
        RECT 132.555 216.145 132.845 216.375 ;
        RECT 123.815 215.850 126.330 215.990 ;
        RECT 123.815 215.805 124.105 215.850 ;
        RECT 109.540 215.510 118.510 215.650 ;
        RECT 109.540 215.450 109.860 215.510 ;
        RECT 86.540 215.170 93.670 215.310 ;
        RECT 93.900 215.310 94.220 215.370 ;
        RECT 96.215 215.310 96.505 215.355 ;
        RECT 93.900 215.170 96.505 215.310 ;
        RECT 86.540 215.110 86.860 215.170 ;
        RECT 93.900 215.110 94.220 215.170 ;
        RECT 96.215 215.125 96.505 215.170 ;
        RECT 106.320 215.110 106.640 215.370 ;
        RECT 115.995 215.310 116.285 215.355 ;
        RECT 116.455 215.310 116.745 215.355 ;
        RECT 115.995 215.170 116.745 215.310 ;
        RECT 118.370 215.310 118.510 215.510 ;
        RECT 118.755 215.465 119.045 215.695 ;
        RECT 119.200 215.650 119.520 215.710 ;
        RECT 126.650 215.650 126.790 216.130 ;
        RECT 119.200 215.510 126.790 215.650 ;
        RECT 127.110 215.650 127.250 216.130 ;
        RECT 132.630 215.990 132.770 216.145 ;
        RECT 133.460 216.130 133.780 216.390 ;
        RECT 134.010 216.330 134.150 216.870 ;
        RECT 134.380 216.870 138.290 217.010 ;
        RECT 134.380 216.810 134.700 216.870 ;
        RECT 135.300 216.670 135.620 216.730 ;
        RECT 136.680 216.670 137.000 216.730 ;
        RECT 138.150 216.715 138.290 216.870 ;
        RECT 140.375 216.825 140.665 217.055 ;
        RECT 145.880 217.010 146.200 217.070 ;
        RECT 150.495 217.010 150.785 217.055 ;
        RECT 145.880 216.870 150.785 217.010 ;
        RECT 135.300 216.530 137.000 216.670 ;
        RECT 135.300 216.470 135.620 216.530 ;
        RECT 136.680 216.470 137.000 216.530 ;
        RECT 138.075 216.485 138.365 216.715 ;
        RECT 138.535 216.670 138.825 216.715 ;
        RECT 140.450 216.670 140.590 216.825 ;
        RECT 145.880 216.810 146.200 216.870 ;
        RECT 150.495 216.825 150.785 216.870 ;
        RECT 154.160 216.810 154.480 217.070 ;
        RECT 145.420 216.670 145.740 216.730 ;
        RECT 138.535 216.530 140.590 216.670 ;
        RECT 141.830 216.530 145.740 216.670 ;
        RECT 138.535 216.485 138.825 216.530 ;
        RECT 137.385 216.330 137.675 216.375 ;
        RECT 138.980 216.330 139.300 216.390 ;
        RECT 134.010 216.190 139.300 216.330 ;
        RECT 137.385 216.145 137.675 216.190 ;
        RECT 138.980 216.130 139.300 216.190 ;
        RECT 139.440 216.130 139.760 216.390 ;
        RECT 139.915 216.330 140.205 216.375 ;
        RECT 141.830 216.330 141.970 216.530 ;
        RECT 145.420 216.470 145.740 216.530 ;
        RECT 139.915 216.190 141.970 216.330 ;
        RECT 139.915 216.145 140.205 216.190 ;
        RECT 142.215 216.145 142.505 216.375 ;
        RECT 142.660 216.330 142.980 216.390 ;
        RECT 151.415 216.330 151.705 216.375 ;
        RECT 142.660 216.190 151.705 216.330 ;
        RECT 128.030 215.850 132.770 215.990 ;
        RECT 133.015 215.990 133.305 216.035 ;
        RECT 139.990 215.990 140.130 216.145 ;
        RECT 133.015 215.850 140.130 215.990 ;
        RECT 128.030 215.710 128.170 215.850 ;
        RECT 133.015 215.805 133.305 215.850 ;
        RECT 141.740 215.790 142.060 216.050 ;
        RECT 142.290 215.990 142.430 216.145 ;
        RECT 142.660 216.130 142.980 216.190 ;
        RECT 151.415 216.145 151.705 216.190 ;
        RECT 153.715 216.330 154.005 216.375 ;
        RECT 154.620 216.330 154.940 216.390 ;
        RECT 153.715 216.190 154.940 216.330 ;
        RECT 153.715 216.145 154.005 216.190 ;
        RECT 154.620 216.130 154.940 216.190 ;
        RECT 152.780 215.990 153.100 216.050 ;
        RECT 142.290 215.850 153.100 215.990 ;
        RECT 127.495 215.650 127.785 215.695 ;
        RECT 127.110 215.510 127.785 215.650 ;
        RECT 119.200 215.450 119.520 215.510 ;
        RECT 127.495 215.465 127.785 215.510 ;
        RECT 127.940 215.450 128.260 215.710 ;
        RECT 142.290 215.650 142.430 215.850 ;
        RECT 152.780 215.790 153.100 215.850 ;
        RECT 136.310 215.510 142.430 215.650 ;
        RECT 136.310 215.310 136.450 215.510 ;
        RECT 118.370 215.170 136.450 215.310 ;
        RECT 115.995 215.125 116.285 215.170 ;
        RECT 116.455 215.125 116.745 215.170 ;
        RECT 136.680 215.110 137.000 215.370 ;
        RECT 138.980 215.310 139.300 215.370 ;
        RECT 140.360 215.310 140.680 215.370 ;
        RECT 141.295 215.310 141.585 215.355 ;
        RECT 138.980 215.170 141.585 215.310 ;
        RECT 138.980 215.110 139.300 215.170 ;
        RECT 140.360 215.110 140.680 215.170 ;
        RECT 141.295 215.125 141.585 215.170 ;
        RECT 152.320 215.110 152.640 215.370 ;
        RECT 2.750 214.490 158.230 214.970 ;
        RECT 13.400 214.290 13.720 214.350 ;
        RECT 14.335 214.290 14.625 214.335 ;
        RECT 23.060 214.290 23.380 214.350 ;
        RECT 13.400 214.150 14.625 214.290 ;
        RECT 13.400 214.090 13.720 214.150 ;
        RECT 14.335 214.105 14.625 214.150 ;
        RECT 15.330 214.150 23.380 214.290 ;
        RECT 8.430 213.810 15.010 213.950 ;
        RECT 4.675 213.270 4.965 213.315 ;
        RECT 4.675 213.130 6.270 213.270 ;
        RECT 4.675 213.085 4.965 213.130 ;
        RECT 5.580 212.390 5.900 212.650 ;
        RECT 6.130 212.635 6.270 213.130 ;
        RECT 7.880 213.070 8.200 213.330 ;
        RECT 8.430 213.315 8.570 213.810 ;
        RECT 9.275 213.425 9.565 213.655 ;
        RECT 12.480 213.610 12.800 213.670 ;
        RECT 12.955 213.610 13.245 213.655 ;
        RECT 12.480 213.470 13.245 213.610 ;
        RECT 8.355 213.085 8.645 213.315 ;
        RECT 9.350 213.270 9.490 213.425 ;
        RECT 12.480 213.410 12.800 213.470 ;
        RECT 12.955 213.425 13.245 213.470 ;
        RECT 14.320 213.270 14.640 213.330 ;
        RECT 9.350 213.130 14.640 213.270 ;
        RECT 14.320 213.070 14.640 213.130 ;
        RECT 12.035 212.930 12.325 212.975 ;
        RECT 13.860 212.930 14.180 212.990 ;
        RECT 12.035 212.790 14.180 212.930 ;
        RECT 12.035 212.745 12.325 212.790 ;
        RECT 13.860 212.730 14.180 212.790 ;
        RECT 6.055 212.405 6.345 212.635 ;
        RECT 10.180 212.390 10.500 212.650 ;
        RECT 12.495 212.590 12.785 212.635 ;
        RECT 12.940 212.590 13.260 212.650 ;
        RECT 12.495 212.450 13.260 212.590 ;
        RECT 14.870 212.590 15.010 213.810 ;
        RECT 15.330 213.315 15.470 214.150 ;
        RECT 23.060 214.090 23.380 214.150 ;
        RECT 26.370 214.150 39.850 214.290 ;
        RECT 17.045 213.950 17.335 213.995 ;
        RECT 18.935 213.950 19.225 213.995 ;
        RECT 22.055 213.950 22.345 213.995 ;
        RECT 17.045 213.810 22.345 213.950 ;
        RECT 17.045 213.765 17.335 213.810 ;
        RECT 18.935 213.765 19.225 213.810 ;
        RECT 22.055 213.765 22.345 213.810 ;
        RECT 22.600 213.950 22.920 214.010 ;
        RECT 26.370 213.950 26.510 214.150 ;
        RECT 22.600 213.810 26.510 213.950 ;
        RECT 31.915 213.950 32.205 213.995 ;
        RECT 35.035 213.950 35.325 213.995 ;
        RECT 36.925 213.950 37.215 213.995 ;
        RECT 31.915 213.810 37.215 213.950 ;
        RECT 22.600 213.750 22.920 213.810 ;
        RECT 31.915 213.765 32.205 213.810 ;
        RECT 35.035 213.765 35.325 213.810 ;
        RECT 36.925 213.765 37.215 213.810 ;
        RECT 16.175 213.610 16.465 213.655 ;
        RECT 18.000 213.610 18.320 213.670 ;
        RECT 16.175 213.470 18.320 213.610 ;
        RECT 16.175 213.425 16.465 213.470 ;
        RECT 18.000 213.410 18.320 213.470 ;
        RECT 20.760 213.610 21.080 213.670 ;
        RECT 26.295 213.610 26.585 213.655 ;
        RECT 20.760 213.470 26.585 213.610 ;
        RECT 20.760 213.410 21.080 213.470 ;
        RECT 26.295 213.425 26.585 213.470 ;
        RECT 35.940 213.610 36.260 213.670 ;
        RECT 36.415 213.610 36.705 213.655 ;
        RECT 35.940 213.470 36.705 213.610 ;
        RECT 35.940 213.410 36.260 213.470 ;
        RECT 36.415 213.425 36.705 213.470 ;
        RECT 39.160 213.410 39.480 213.670 ;
        RECT 39.710 213.610 39.850 214.150 ;
        RECT 43.300 214.090 43.620 214.350 ;
        RECT 52.500 214.090 52.820 214.350 ;
        RECT 55.275 214.290 55.565 214.335 ;
        RECT 58.940 214.290 59.260 214.350 ;
        RECT 69.980 214.290 70.300 214.350 ;
        RECT 55.275 214.150 59.260 214.290 ;
        RECT 55.275 214.105 55.565 214.150 ;
        RECT 58.940 214.090 59.260 214.150 ;
        RECT 59.490 214.150 70.300 214.290 ;
        RECT 40.080 213.950 40.400 214.010 ;
        RECT 44.695 213.950 44.985 213.995 ;
        RECT 59.490 213.950 59.630 214.150 ;
        RECT 69.980 214.090 70.300 214.150 ;
        RECT 70.455 214.290 70.745 214.335 ;
        RECT 76.420 214.290 76.740 214.350 ;
        RECT 70.455 214.150 76.740 214.290 ;
        RECT 70.455 214.105 70.745 214.150 ;
        RECT 76.420 214.090 76.740 214.150 ;
        RECT 77.815 214.290 78.105 214.335 ;
        RECT 80.100 214.290 80.420 214.350 ;
        RECT 77.815 214.150 80.420 214.290 ;
        RECT 77.815 214.105 78.105 214.150 ;
        RECT 80.100 214.090 80.420 214.150 ;
        RECT 81.480 214.090 81.800 214.350 ;
        RECT 89.315 214.290 89.605 214.335 ;
        RECT 89.760 214.290 90.080 214.350 ;
        RECT 89.315 214.150 90.080 214.290 ;
        RECT 89.315 214.105 89.605 214.150 ;
        RECT 89.760 214.090 90.080 214.150 ;
        RECT 91.140 214.290 91.460 214.350 ;
        RECT 103.560 214.290 103.880 214.350 ;
        RECT 109.540 214.290 109.860 214.350 ;
        RECT 91.140 214.150 103.330 214.290 ;
        RECT 91.140 214.090 91.460 214.150 ;
        RECT 40.080 213.810 44.985 213.950 ;
        RECT 40.080 213.750 40.400 213.810 ;
        RECT 44.695 213.765 44.985 213.810 ;
        RECT 54.430 213.810 59.630 213.950 ;
        RECT 60.750 213.950 61.040 213.995 ;
        RECT 63.530 213.950 63.820 213.995 ;
        RECT 65.390 213.950 65.680 213.995 ;
        RECT 60.750 213.810 65.680 213.950 ;
        RECT 47.915 213.610 48.205 213.655 ;
        RECT 49.740 213.610 50.060 213.670 ;
        RECT 39.710 213.470 47.670 213.610 ;
        RECT 15.255 213.085 15.545 213.315 ;
        RECT 16.640 213.270 16.930 213.315 ;
        RECT 18.475 213.270 18.765 213.315 ;
        RECT 22.055 213.270 22.345 213.315 ;
        RECT 16.640 213.130 22.345 213.270 ;
        RECT 16.640 213.085 16.930 213.130 ;
        RECT 18.475 213.085 18.765 213.130 ;
        RECT 22.055 213.085 22.345 213.130 ;
        RECT 16.160 212.930 16.480 212.990 ;
        RECT 23.135 212.975 23.425 213.290 ;
        RECT 17.555 212.930 17.845 212.975 ;
        RECT 16.160 212.790 17.845 212.930 ;
        RECT 16.160 212.730 16.480 212.790 ;
        RECT 17.555 212.745 17.845 212.790 ;
        RECT 19.835 212.930 20.485 212.975 ;
        RECT 23.135 212.930 23.725 212.975 ;
        RECT 24.900 212.930 25.220 212.990 ;
        RECT 30.835 212.975 31.125 213.290 ;
        RECT 31.915 213.270 32.205 213.315 ;
        RECT 35.495 213.270 35.785 213.315 ;
        RECT 37.330 213.270 37.620 213.315 ;
        RECT 31.915 213.130 37.620 213.270 ;
        RECT 31.915 213.085 32.205 213.130 ;
        RECT 35.495 213.085 35.785 213.130 ;
        RECT 37.330 213.085 37.620 213.130 ;
        RECT 37.795 213.270 38.085 213.315 ;
        RECT 43.775 213.270 44.065 213.315 ;
        RECT 46.980 213.270 47.300 213.330 ;
        RECT 37.795 213.130 40.310 213.270 ;
        RECT 37.795 213.085 38.085 213.130 ;
        RECT 19.835 212.790 25.220 212.930 ;
        RECT 19.835 212.745 20.485 212.790 ;
        RECT 23.435 212.745 23.725 212.790 ;
        RECT 24.900 212.730 25.220 212.790 ;
        RECT 27.675 212.745 27.965 212.975 ;
        RECT 30.535 212.930 31.125 212.975 ;
        RECT 33.775 212.930 34.425 212.975 ;
        RECT 30.535 212.790 34.790 212.930 ;
        RECT 30.535 212.745 30.825 212.790 ;
        RECT 33.775 212.745 34.425 212.790 ;
        RECT 20.760 212.590 21.080 212.650 ;
        RECT 22.600 212.590 22.920 212.650 ;
        RECT 14.870 212.450 22.920 212.590 ;
        RECT 27.750 212.590 27.890 212.745 ;
        RECT 34.650 212.650 34.790 212.790 ;
        RECT 32.260 212.590 32.580 212.650 ;
        RECT 27.750 212.450 32.580 212.590 ;
        RECT 12.495 212.405 12.785 212.450 ;
        RECT 12.940 212.390 13.260 212.450 ;
        RECT 20.760 212.390 21.080 212.450 ;
        RECT 22.600 212.390 22.920 212.450 ;
        RECT 32.260 212.390 32.580 212.450 ;
        RECT 34.560 212.390 34.880 212.650 ;
        RECT 39.160 212.590 39.480 212.650 ;
        RECT 40.170 212.590 40.310 213.130 ;
        RECT 43.775 213.130 47.300 213.270 ;
        RECT 43.775 213.085 44.065 213.130 ;
        RECT 46.980 213.070 47.300 213.130 ;
        RECT 40.555 212.930 40.845 212.975 ;
        RECT 44.220 212.930 44.540 212.990 ;
        RECT 40.555 212.790 44.540 212.930 ;
        RECT 40.555 212.745 40.845 212.790 ;
        RECT 44.220 212.730 44.540 212.790 ;
        RECT 45.140 212.730 45.460 212.990 ;
        RECT 46.535 212.930 46.825 212.975 ;
        RECT 47.530 212.930 47.670 213.470 ;
        RECT 47.915 213.470 50.060 213.610 ;
        RECT 47.915 213.425 48.205 213.470 ;
        RECT 49.740 213.410 50.060 213.470 ;
        RECT 50.215 213.610 50.505 213.655 ;
        RECT 53.880 213.610 54.200 213.670 ;
        RECT 50.215 213.470 54.200 213.610 ;
        RECT 50.215 213.425 50.505 213.470 ;
        RECT 53.880 213.410 54.200 213.470 ;
        RECT 54.430 213.270 54.570 213.810 ;
        RECT 60.750 213.765 61.040 213.810 ;
        RECT 63.530 213.765 63.820 213.810 ;
        RECT 65.390 213.765 65.680 213.810 ;
        RECT 69.060 213.950 69.380 214.010 ;
        RECT 82.860 213.950 83.180 214.010 ;
        RECT 69.060 213.810 83.180 213.950 ;
        RECT 69.060 213.750 69.380 213.810 ;
        RECT 82.860 213.750 83.180 213.810 ;
        RECT 84.255 213.950 84.545 213.995 ;
        RECT 84.255 213.810 86.310 213.950 ;
        RECT 84.255 213.765 84.545 213.810 ;
        RECT 56.885 213.610 57.175 213.655 ;
        RECT 64.920 213.610 65.240 213.670 ;
        RECT 78.720 213.610 79.040 213.670 ;
        RECT 56.885 213.470 67.910 213.610 ;
        RECT 56.885 213.425 57.175 213.470 ;
        RECT 64.920 213.410 65.240 213.470 ;
        RECT 46.535 212.790 47.670 212.930 ;
        RECT 49.830 213.130 54.570 213.270 ;
        RECT 55.735 213.270 56.025 213.315 ;
        RECT 58.020 213.270 58.340 213.330 ;
        RECT 55.735 213.130 58.340 213.270 ;
        RECT 46.535 212.745 46.825 212.790 ;
        RECT 42.840 212.590 43.160 212.650 ;
        RECT 45.230 212.590 45.370 212.730 ;
        RECT 39.160 212.450 45.370 212.590 ;
        RECT 46.995 212.590 47.285 212.635 ;
        RECT 49.830 212.590 49.970 213.130 ;
        RECT 55.735 213.085 56.025 213.130 ;
        RECT 58.020 213.070 58.340 213.130 ;
        RECT 60.750 213.270 61.040 213.315 ;
        RECT 64.015 213.270 64.305 213.315 ;
        RECT 64.460 213.270 64.780 213.330 ;
        RECT 60.750 213.130 63.285 213.270 ;
        RECT 60.750 213.085 61.040 213.130 ;
        RECT 58.890 212.930 59.180 212.975 ;
        RECT 61.240 212.930 61.560 212.990 ;
        RECT 63.070 212.975 63.285 213.130 ;
        RECT 64.015 213.130 64.780 213.270 ;
        RECT 64.015 213.085 64.305 213.130 ;
        RECT 64.460 213.070 64.780 213.130 ;
        RECT 65.840 213.070 66.160 213.330 ;
        RECT 67.770 213.315 67.910 213.470 ;
        RECT 72.370 213.470 79.040 213.610 ;
        RECT 67.695 213.085 67.985 213.315 ;
        RECT 70.900 213.270 71.220 213.330 ;
        RECT 71.375 213.270 71.665 213.315 ;
        RECT 70.900 213.130 71.665 213.270 ;
        RECT 70.900 213.070 71.220 213.130 ;
        RECT 71.375 213.085 71.665 213.130 ;
        RECT 71.820 213.070 72.140 213.330 ;
        RECT 62.150 212.930 62.440 212.975 ;
        RECT 58.890 212.790 62.440 212.930 ;
        RECT 58.890 212.745 59.180 212.790 ;
        RECT 61.240 212.730 61.560 212.790 ;
        RECT 62.150 212.745 62.440 212.790 ;
        RECT 63.070 212.930 63.360 212.975 ;
        RECT 64.930 212.930 65.220 212.975 ;
        RECT 63.070 212.790 65.220 212.930 ;
        RECT 63.070 212.745 63.360 212.790 ;
        RECT 64.930 212.745 65.220 212.790 ;
        RECT 68.155 212.930 68.445 212.975 ;
        RECT 72.370 212.930 72.510 213.470 ;
        RECT 78.720 213.410 79.040 213.470 ;
        RECT 73.660 213.070 73.980 213.330 ;
        RECT 74.120 213.070 74.440 213.330 ;
        RECT 75.040 213.070 75.360 213.330 ;
        RECT 75.500 213.270 75.820 213.330 ;
        RECT 77.355 213.270 77.645 213.315 ;
        RECT 77.800 213.270 78.120 213.330 ;
        RECT 75.500 213.130 78.120 213.270 ;
        RECT 75.500 213.070 75.820 213.130 ;
        RECT 77.355 213.085 77.645 213.130 ;
        RECT 77.800 213.070 78.120 213.130 ;
        RECT 78.260 213.070 78.580 213.330 ;
        RECT 79.640 213.070 79.960 213.330 ;
        RECT 81.955 213.270 82.245 213.315 ;
        RECT 82.400 213.270 82.720 213.330 ;
        RECT 82.950 213.315 83.090 213.750 ;
        RECT 86.170 213.655 86.310 213.810 ;
        RECT 88.395 213.765 88.685 213.995 ;
        RECT 92.060 213.950 92.380 214.010 ;
        RECT 89.620 213.810 92.380 213.950 ;
        RECT 83.870 213.470 85.390 213.610 ;
        RECT 83.870 213.315 84.010 213.470 ;
        RECT 85.250 213.330 85.390 213.470 ;
        RECT 86.095 213.425 86.385 213.655 ;
        RECT 87.475 213.610 87.765 213.655 ;
        RECT 88.470 213.610 88.610 213.765 ;
        RECT 87.475 213.470 88.610 213.610 ;
        RECT 87.475 213.425 87.765 213.470 ;
        RECT 81.955 213.130 82.720 213.270 ;
        RECT 81.955 213.085 82.245 213.130 ;
        RECT 82.400 213.070 82.720 213.130 ;
        RECT 82.875 213.085 83.165 213.315 ;
        RECT 83.795 213.085 84.085 213.315 ;
        RECT 84.700 213.070 85.020 213.330 ;
        RECT 85.160 213.070 85.480 213.330 ;
        RECT 86.540 213.070 86.860 213.330 ;
        RECT 87.015 213.270 87.305 213.315 ;
        RECT 87.920 213.270 88.240 213.330 ;
        RECT 89.620 213.270 89.760 213.810 ;
        RECT 92.060 213.750 92.380 213.810 ;
        RECT 92.980 213.950 93.300 214.010 ;
        RECT 98.960 213.950 99.280 214.010 ;
        RECT 92.980 213.810 99.280 213.950 ;
        RECT 92.980 213.750 93.300 213.810 ;
        RECT 98.960 213.750 99.280 213.810 ;
        RECT 101.260 213.750 101.580 214.010 ;
        RECT 101.735 213.950 102.025 213.995 ;
        RECT 103.190 213.950 103.330 214.150 ;
        RECT 103.560 214.150 109.860 214.290 ;
        RECT 103.560 214.090 103.880 214.150 ;
        RECT 109.540 214.090 109.860 214.150 ;
        RECT 112.760 214.090 113.080 214.350 ;
        RECT 113.235 214.290 113.525 214.335 ;
        RECT 116.440 214.290 116.760 214.350 ;
        RECT 117.820 214.290 118.140 214.350 ;
        RECT 113.235 214.150 116.760 214.290 ;
        RECT 113.235 214.105 113.525 214.150 ;
        RECT 116.440 214.090 116.760 214.150 ;
        RECT 117.450 214.150 118.140 214.290 ;
        RECT 112.850 213.950 112.990 214.090 ;
        RECT 117.450 213.950 117.590 214.150 ;
        RECT 117.820 214.090 118.140 214.150 ;
        RECT 123.340 214.090 123.660 214.350 ;
        RECT 123.815 214.290 124.105 214.335 ;
        RECT 125.640 214.290 125.960 214.350 ;
        RECT 145.420 214.290 145.740 214.350 ;
        RECT 146.815 214.290 147.105 214.335 ;
        RECT 123.815 214.150 125.960 214.290 ;
        RECT 123.815 214.105 124.105 214.150 ;
        RECT 125.640 214.090 125.960 214.150 ;
        RECT 131.020 214.150 145.190 214.290 ;
        RECT 127.480 213.950 127.800 214.010 ;
        RECT 131.020 213.950 131.160 214.150 ;
        RECT 101.735 213.810 102.870 213.950 ;
        RECT 103.190 213.810 108.390 213.950 ;
        RECT 112.850 213.810 117.590 213.950 ;
        RECT 117.910 213.810 131.160 213.950 ;
        RECT 101.735 213.765 102.025 213.810 ;
        RECT 92.520 213.610 92.840 213.670 ;
        RECT 95.740 213.610 96.060 213.670 ;
        RECT 101.350 213.610 101.490 213.750 ;
        RECT 92.520 213.470 96.060 213.610 ;
        RECT 92.520 213.410 92.840 213.470 ;
        RECT 95.740 213.410 96.060 213.470 ;
        RECT 100.890 213.470 101.490 213.610 ;
        RECT 102.730 213.610 102.870 213.810 ;
        RECT 102.730 213.470 106.550 213.610 ;
        RECT 98.500 213.270 98.820 213.330 ;
        RECT 100.890 213.315 101.030 213.470 ;
        RECT 106.410 213.330 106.550 213.470 ;
        RECT 87.015 213.130 89.760 213.270 ;
        RECT 90.310 213.130 98.820 213.270 ;
        RECT 87.015 213.085 87.305 213.130 ;
        RECT 87.920 213.070 88.240 213.130 ;
        RECT 76.880 212.930 77.200 212.990 ;
        RECT 89.300 212.975 89.620 212.990 ;
        RECT 90.310 212.975 90.450 213.130 ;
        RECT 98.500 213.070 98.820 213.130 ;
        RECT 100.815 213.085 101.105 213.315 ;
        RECT 101.260 213.070 101.580 213.330 ;
        RECT 102.195 213.085 102.485 213.315 ;
        RECT 103.560 213.270 103.880 213.330 ;
        RECT 105.875 213.270 106.165 213.315 ;
        RECT 103.560 213.130 106.165 213.270 ;
        RECT 68.155 212.790 72.510 212.930 ;
        RECT 72.830 212.790 77.200 212.930 ;
        RECT 68.155 212.745 68.445 212.790 ;
        RECT 46.995 212.450 49.970 212.590 ;
        RECT 39.160 212.390 39.480 212.450 ;
        RECT 42.840 212.390 43.160 212.450 ;
        RECT 46.995 212.405 47.285 212.450 ;
        RECT 50.660 212.390 50.980 212.650 ;
        RECT 52.960 212.590 53.280 212.650 ;
        RECT 58.020 212.590 58.340 212.650 ;
        RECT 72.830 212.635 72.970 212.790 ;
        RECT 76.880 212.730 77.200 212.790 ;
        RECT 80.190 212.790 87.690 212.930 ;
        RECT 52.960 212.450 58.340 212.590 ;
        RECT 52.960 212.390 53.280 212.450 ;
        RECT 58.020 212.390 58.340 212.450 ;
        RECT 72.755 212.405 73.045 212.635 ;
        RECT 73.215 212.590 73.505 212.635 ;
        RECT 74.135 212.590 74.425 212.635 ;
        RECT 73.215 212.450 74.425 212.590 ;
        RECT 73.215 212.405 73.505 212.450 ;
        RECT 74.135 212.405 74.425 212.450 ;
        RECT 74.580 212.590 74.900 212.650 ;
        RECT 80.190 212.635 80.330 212.790 ;
        RECT 87.550 212.650 87.690 212.790 ;
        RECT 89.235 212.745 89.620 212.975 ;
        RECT 90.235 212.745 90.525 212.975 ;
        RECT 102.270 212.930 102.410 213.085 ;
        RECT 103.560 213.070 103.880 213.130 ;
        RECT 105.875 213.085 106.165 213.130 ;
        RECT 106.320 213.070 106.640 213.330 ;
        RECT 106.795 213.270 107.085 213.315 ;
        RECT 106.795 213.130 107.470 213.270 ;
        RECT 106.795 213.085 107.085 213.130 ;
        RECT 90.770 212.790 102.410 212.930 ;
        RECT 89.300 212.730 89.620 212.745 ;
        RECT 80.115 212.590 80.405 212.635 ;
        RECT 74.580 212.450 80.405 212.590 ;
        RECT 74.580 212.390 74.900 212.450 ;
        RECT 80.115 212.405 80.405 212.450 ;
        RECT 80.575 212.590 80.865 212.635 ;
        RECT 82.415 212.590 82.705 212.635 ;
        RECT 82.860 212.590 83.180 212.650 ;
        RECT 80.575 212.450 83.180 212.590 ;
        RECT 80.575 212.405 80.865 212.450 ;
        RECT 82.415 212.405 82.705 212.450 ;
        RECT 82.860 212.390 83.180 212.450 ;
        RECT 84.700 212.590 85.020 212.650 ;
        RECT 85.175 212.590 85.465 212.635 ;
        RECT 84.700 212.450 85.465 212.590 ;
        RECT 84.700 212.390 85.020 212.450 ;
        RECT 85.175 212.405 85.465 212.450 ;
        RECT 87.460 212.590 87.780 212.650 ;
        RECT 90.770 212.590 90.910 212.790 ;
        RECT 104.480 212.730 104.800 212.990 ;
        RECT 107.330 212.650 107.470 213.130 ;
        RECT 107.700 213.070 108.020 213.330 ;
        RECT 108.250 213.270 108.390 213.810 ;
        RECT 117.910 213.670 118.050 213.810 ;
        RECT 127.480 213.750 127.800 213.810 ;
        RECT 110.920 213.610 111.240 213.670 ;
        RECT 112.775 213.610 113.065 213.655 ;
        RECT 110.920 213.470 113.065 213.610 ;
        RECT 110.920 213.410 111.240 213.470 ;
        RECT 112.775 213.425 113.065 213.470 ;
        RECT 117.820 213.410 118.140 213.670 ;
        RECT 118.280 213.610 118.600 213.670 ;
        RECT 118.280 213.470 122.190 213.610 ;
        RECT 118.280 213.410 118.600 213.470 ;
        RECT 112.315 213.270 112.605 213.315 ;
        RECT 121.500 213.270 121.820 213.330 ;
        RECT 108.250 213.130 111.150 213.270 ;
        RECT 111.010 212.975 111.150 213.130 ;
        RECT 112.315 213.130 121.820 213.270 ;
        RECT 112.315 213.085 112.605 213.130 ;
        RECT 121.500 213.070 121.820 213.130 ;
        RECT 110.935 212.930 111.225 212.975 ;
        RECT 116.900 212.930 117.220 212.990 ;
        RECT 110.935 212.790 117.220 212.930 ;
        RECT 110.935 212.745 111.225 212.790 ;
        RECT 116.900 212.730 117.220 212.790 ;
        RECT 118.740 212.730 119.060 212.990 ;
        RECT 87.460 212.450 90.910 212.590 ;
        RECT 91.600 212.590 91.920 212.650 ;
        RECT 96.660 212.590 96.980 212.650 ;
        RECT 91.600 212.450 96.980 212.590 ;
        RECT 87.460 212.390 87.780 212.450 ;
        RECT 91.600 212.390 91.920 212.450 ;
        RECT 96.660 212.390 96.980 212.450 ;
        RECT 99.880 212.390 100.200 212.650 ;
        RECT 101.260 212.590 101.580 212.650 ;
        RECT 102.640 212.590 102.960 212.650 ;
        RECT 101.260 212.450 102.960 212.590 ;
        RECT 101.260 212.390 101.580 212.450 ;
        RECT 102.640 212.390 102.960 212.450 ;
        RECT 107.240 212.390 107.560 212.650 ;
        RECT 111.395 212.590 111.685 212.635 ;
        RECT 112.300 212.590 112.620 212.650 ;
        RECT 113.220 212.590 113.540 212.650 ;
        RECT 118.830 212.590 118.970 212.730 ;
        RECT 111.395 212.450 118.970 212.590 ;
        RECT 122.050 212.590 122.190 213.470 ;
        RECT 122.880 213.410 123.200 213.670 ;
        RECT 124.275 213.610 124.565 213.655 ;
        RECT 127.940 213.610 128.260 213.670 ;
        RECT 124.275 213.470 128.260 213.610 ;
        RECT 124.275 213.425 124.565 213.470 ;
        RECT 122.970 213.270 123.110 213.410 ;
        RECT 124.810 213.330 124.950 213.470 ;
        RECT 127.940 213.410 128.260 213.470 ;
        RECT 138.075 213.610 138.365 213.655 ;
        RECT 142.200 213.610 142.520 213.670 ;
        RECT 138.075 213.470 142.520 213.610 ;
        RECT 145.050 213.610 145.190 214.150 ;
        RECT 145.420 214.150 147.105 214.290 ;
        RECT 145.420 214.090 145.740 214.150 ;
        RECT 146.815 214.105 147.105 214.150 ;
        RECT 147.260 214.090 147.580 214.350 ;
        RECT 152.320 214.290 152.640 214.350 ;
        RECT 155.555 214.290 155.845 214.335 ;
        RECT 152.320 214.150 155.845 214.290 ;
        RECT 152.320 214.090 152.640 214.150 ;
        RECT 155.555 214.105 155.845 214.150 ;
        RECT 152.780 213.750 153.100 214.010 ;
        RECT 150.940 213.610 151.260 213.670 ;
        RECT 154.160 213.610 154.480 213.670 ;
        RECT 145.050 213.470 145.650 213.610 ;
        RECT 138.075 213.425 138.365 213.470 ;
        RECT 142.200 213.410 142.520 213.470 ;
        RECT 122.970 213.205 123.115 213.270 ;
        RECT 122.900 212.975 123.190 213.205 ;
        RECT 124.720 213.070 125.040 213.330 ;
        RECT 135.300 213.270 135.620 213.330 ;
        RECT 135.765 213.270 136.055 213.315 ;
        RECT 135.300 213.130 136.055 213.270 ;
        RECT 135.300 213.070 135.620 213.130 ;
        RECT 135.765 213.085 136.055 213.130 ;
        RECT 137.385 213.085 137.675 213.315 ;
        RECT 143.120 213.270 143.440 213.330 ;
        RECT 145.510 213.270 145.650 213.470 ;
        RECT 150.940 213.470 156.230 213.610 ;
        RECT 150.940 213.410 151.260 213.470 ;
        RECT 154.160 213.410 154.480 213.470 ;
        RECT 147.275 213.270 147.565 213.315 ;
        RECT 149.560 213.270 149.880 213.330 ;
        RECT 152.795 213.270 153.085 213.315 ;
        RECT 143.120 213.140 143.810 213.270 ;
        RECT 144.975 213.140 145.265 213.185 ;
        RECT 143.120 213.130 145.265 213.140 ;
        RECT 145.510 213.130 147.030 213.270 ;
        RECT 124.260 212.930 124.580 212.990 ;
        RECT 137.460 212.930 137.600 213.085 ;
        RECT 143.120 213.070 143.440 213.130 ;
        RECT 143.670 213.000 145.265 213.130 ;
        RECT 144.975 212.955 145.265 213.000 ;
        RECT 145.880 212.975 146.200 212.990 ;
        RECT 124.260 212.790 137.600 212.930 ;
        RECT 124.260 212.730 124.580 212.790 ;
        RECT 145.880 212.745 146.315 212.975 ;
        RECT 146.890 212.930 147.030 213.130 ;
        RECT 147.275 213.130 149.880 213.270 ;
        RECT 147.275 213.085 147.565 213.130 ;
        RECT 149.560 213.070 149.880 213.130 ;
        RECT 151.490 213.130 153.085 213.270 ;
        RECT 151.490 212.990 151.630 213.130 ;
        RECT 152.795 213.085 153.085 213.130 ;
        RECT 153.700 213.070 154.020 213.330 ;
        RECT 155.080 213.070 155.400 213.330 ;
        RECT 156.090 213.315 156.230 213.470 ;
        RECT 156.015 213.085 156.305 213.315 ;
        RECT 147.720 212.930 148.040 212.990 ;
        RECT 148.655 212.930 148.945 212.975 ;
        RECT 146.890 212.790 148.945 212.930 ;
        RECT 145.880 212.730 146.200 212.745 ;
        RECT 147.720 212.730 148.040 212.790 ;
        RECT 148.655 212.745 148.945 212.790 ;
        RECT 151.400 212.730 151.720 212.990 ;
        RECT 126.560 212.590 126.880 212.650 ;
        RECT 122.050 212.450 126.880 212.590 ;
        RECT 111.395 212.405 111.685 212.450 ;
        RECT 112.300 212.390 112.620 212.450 ;
        RECT 113.220 212.390 113.540 212.450 ;
        RECT 126.560 212.390 126.880 212.450 ;
        RECT 128.400 212.590 128.720 212.650 ;
        RECT 133.920 212.590 134.240 212.650 ;
        RECT 128.400 212.450 134.240 212.590 ;
        RECT 128.400 212.390 128.720 212.450 ;
        RECT 133.920 212.390 134.240 212.450 ;
        RECT 134.840 212.390 135.160 212.650 ;
        RECT 135.760 212.390 136.080 212.650 ;
        RECT 141.740 212.590 142.060 212.650 ;
        RECT 145.435 212.590 145.725 212.635 ;
        RECT 149.115 212.590 149.405 212.635 ;
        RECT 150.480 212.590 150.800 212.650 ;
        RECT 141.740 212.450 150.800 212.590 ;
        RECT 141.740 212.390 142.060 212.450 ;
        RECT 145.435 212.405 145.725 212.450 ;
        RECT 149.115 212.405 149.405 212.450 ;
        RECT 150.480 212.390 150.800 212.450 ;
        RECT 2.750 211.770 159.030 212.250 ;
        RECT 5.580 211.370 5.900 211.630 ;
        RECT 19.840 211.570 20.160 211.630 ;
        RECT 45.140 211.570 45.460 211.630 ;
        RECT 19.840 211.430 37.550 211.570 ;
        RECT 19.840 211.370 20.160 211.430 ;
        RECT 5.670 211.230 5.810 211.370 ;
        RECT 6.055 211.230 6.345 211.275 ;
        RECT 5.670 211.090 6.345 211.230 ;
        RECT 6.055 211.045 6.345 211.090 ;
        RECT 8.335 211.230 8.985 211.275 ;
        RECT 11.935 211.230 12.225 211.275 ;
        RECT 8.335 211.090 12.225 211.230 ;
        RECT 8.335 211.045 8.985 211.090 ;
        RECT 11.635 211.045 12.225 211.090 ;
        RECT 14.795 211.230 15.085 211.275 ;
        RECT 16.620 211.230 16.940 211.290 ;
        RECT 24.900 211.275 25.220 211.290 ;
        RECT 14.795 211.090 16.940 211.230 ;
        RECT 14.795 211.045 15.085 211.090 ;
        RECT 5.140 210.890 5.430 210.935 ;
        RECT 6.975 210.890 7.265 210.935 ;
        RECT 10.555 210.890 10.845 210.935 ;
        RECT 5.140 210.750 10.845 210.890 ;
        RECT 5.140 210.705 5.430 210.750 ;
        RECT 6.975 210.705 7.265 210.750 ;
        RECT 10.555 210.705 10.845 210.750 ;
        RECT 11.100 210.890 11.420 210.950 ;
        RECT 11.635 210.890 11.925 211.045 ;
        RECT 16.620 211.030 16.940 211.090 ;
        RECT 18.940 211.230 19.230 211.275 ;
        RECT 20.800 211.230 21.090 211.275 ;
        RECT 18.940 211.090 21.090 211.230 ;
        RECT 18.940 211.045 19.230 211.090 ;
        RECT 20.800 211.045 21.090 211.090 ;
        RECT 21.720 211.230 22.010 211.275 ;
        RECT 24.900 211.230 25.270 211.275 ;
        RECT 25.450 211.230 25.590 211.430 ;
        RECT 37.410 211.290 37.550 211.430 ;
        RECT 45.140 211.430 48.360 211.570 ;
        RECT 45.140 211.370 45.460 211.430 ;
        RECT 21.720 211.090 25.590 211.230 ;
        RECT 28.120 211.230 28.440 211.290 ;
        RECT 30.895 211.230 31.185 211.275 ;
        RECT 28.120 211.090 31.185 211.230 ;
        RECT 21.720 211.045 22.010 211.090 ;
        RECT 24.900 211.045 25.270 211.090 ;
        RECT 13.400 210.890 13.720 210.950 ;
        RECT 11.100 210.750 13.720 210.890 ;
        RECT 11.100 210.690 11.420 210.750 ;
        RECT 11.635 210.730 11.925 210.750 ;
        RECT 13.400 210.690 13.720 210.750 ;
        RECT 18.000 210.890 18.320 210.950 ;
        RECT 20.875 210.890 21.090 211.045 ;
        RECT 24.900 211.030 25.220 211.045 ;
        RECT 28.120 211.030 28.440 211.090 ;
        RECT 30.895 211.045 31.185 211.090 ;
        RECT 33.175 211.230 33.825 211.275 ;
        RECT 34.560 211.230 34.880 211.290 ;
        RECT 36.775 211.230 37.065 211.275 ;
        RECT 33.175 211.090 37.065 211.230 ;
        RECT 33.175 211.045 33.825 211.090 ;
        RECT 34.560 211.030 34.880 211.090 ;
        RECT 36.475 211.045 37.065 211.090 ;
        RECT 23.120 210.890 23.410 210.935 ;
        RECT 18.000 210.750 20.530 210.890 ;
        RECT 20.875 210.750 23.410 210.890 ;
        RECT 18.000 210.690 18.320 210.750 ;
        RECT 4.675 210.365 4.965 210.595 ;
        RECT 15.240 210.550 15.560 210.610 ;
        RECT 19.855 210.550 20.145 210.595 ;
        RECT 15.240 210.410 20.145 210.550 ;
        RECT 20.390 210.550 20.530 210.750 ;
        RECT 23.120 210.705 23.410 210.750 ;
        RECT 27.660 210.890 27.980 210.950 ;
        RECT 29.515 210.890 29.805 210.935 ;
        RECT 27.660 210.750 29.805 210.890 ;
        RECT 27.660 210.690 27.980 210.750 ;
        RECT 29.515 210.705 29.805 210.750 ;
        RECT 29.980 210.890 30.270 210.935 ;
        RECT 31.815 210.890 32.105 210.935 ;
        RECT 35.395 210.890 35.685 210.935 ;
        RECT 29.980 210.750 35.685 210.890 ;
        RECT 29.980 210.705 30.270 210.750 ;
        RECT 31.815 210.705 32.105 210.750 ;
        RECT 35.395 210.705 35.685 210.750 ;
        RECT 36.475 210.730 36.765 211.045 ;
        RECT 37.320 211.030 37.640 211.290 ;
        RECT 43.755 211.230 44.405 211.275 ;
        RECT 47.355 211.230 47.645 211.275 ;
        RECT 43.755 211.090 47.645 211.230 ;
        RECT 43.755 211.045 44.405 211.090 ;
        RECT 47.055 211.045 47.645 211.090 ;
        RECT 39.160 210.890 39.480 210.950 ;
        RECT 40.095 210.890 40.385 210.935 ;
        RECT 39.160 210.750 40.385 210.890 ;
        RECT 39.160 210.690 39.480 210.750 ;
        RECT 40.095 210.705 40.385 210.750 ;
        RECT 40.560 210.890 40.850 210.935 ;
        RECT 42.395 210.890 42.685 210.935 ;
        RECT 45.975 210.890 46.265 210.935 ;
        RECT 40.560 210.750 46.265 210.890 ;
        RECT 40.560 210.705 40.850 210.750 ;
        RECT 42.395 210.705 42.685 210.750 ;
        RECT 45.975 210.705 46.265 210.750 ;
        RECT 47.055 210.730 47.345 211.045 ;
        RECT 30.880 210.550 31.200 210.610 ;
        RECT 20.390 210.410 31.200 210.550 ;
        RECT 4.750 209.930 4.890 210.365 ;
        RECT 15.240 210.350 15.560 210.410 ;
        RECT 19.855 210.365 20.145 210.410 ;
        RECT 30.880 210.350 31.200 210.410 ;
        RECT 33.180 210.550 33.500 210.610 ;
        RECT 39.635 210.550 39.925 210.595 ;
        RECT 33.180 210.410 39.925 210.550 ;
        RECT 33.180 210.350 33.500 210.410 ;
        RECT 39.635 210.365 39.925 210.410 ;
        RECT 41.475 210.550 41.765 210.595 ;
        RECT 44.680 210.550 45.000 210.610 ;
        RECT 41.475 210.410 45.000 210.550 ;
        RECT 41.475 210.365 41.765 210.410 ;
        RECT 44.680 210.350 45.000 210.410 ;
        RECT 5.545 210.210 5.835 210.255 ;
        RECT 7.435 210.210 7.725 210.255 ;
        RECT 10.555 210.210 10.845 210.255 ;
        RECT 18.000 210.210 18.320 210.270 ;
        RECT 5.545 210.070 10.845 210.210 ;
        RECT 5.545 210.025 5.835 210.070 ;
        RECT 7.435 210.025 7.725 210.070 ;
        RECT 10.555 210.025 10.845 210.070 ;
        RECT 12.110 210.070 18.320 210.210 ;
        RECT 4.660 209.870 4.980 209.930 ;
        RECT 12.110 209.870 12.250 210.070 ;
        RECT 18.000 210.010 18.320 210.070 ;
        RECT 18.480 210.210 18.770 210.255 ;
        RECT 20.340 210.210 20.630 210.255 ;
        RECT 23.120 210.210 23.410 210.255 ;
        RECT 18.480 210.070 23.410 210.210 ;
        RECT 18.480 210.025 18.770 210.070 ;
        RECT 20.340 210.025 20.630 210.070 ;
        RECT 23.120 210.025 23.410 210.070 ;
        RECT 30.385 210.210 30.675 210.255 ;
        RECT 32.275 210.210 32.565 210.255 ;
        RECT 35.395 210.210 35.685 210.255 ;
        RECT 30.385 210.070 35.685 210.210 ;
        RECT 30.385 210.025 30.675 210.070 ;
        RECT 32.275 210.025 32.565 210.070 ;
        RECT 35.395 210.025 35.685 210.070 ;
        RECT 40.965 210.210 41.255 210.255 ;
        RECT 42.855 210.210 43.145 210.255 ;
        RECT 45.975 210.210 46.265 210.255 ;
        RECT 40.965 210.070 46.265 210.210 ;
        RECT 47.070 210.210 47.210 210.730 ;
        RECT 48.220 210.550 48.360 211.430 ;
        RECT 52.040 211.370 52.360 211.630 ;
        RECT 61.240 211.570 61.560 211.630 ;
        RECT 52.590 211.430 61.560 211.570 ;
        RECT 50.200 210.890 50.520 210.950 ;
        RECT 51.135 210.890 51.425 210.935 ;
        RECT 52.590 210.890 52.730 211.430 ;
        RECT 61.240 211.370 61.560 211.430 ;
        RECT 62.635 211.570 62.925 211.615 ;
        RECT 65.840 211.570 66.160 211.630 ;
        RECT 62.635 211.430 66.160 211.570 ;
        RECT 62.635 211.385 62.925 211.430 ;
        RECT 65.840 211.370 66.160 211.430 ;
        RECT 82.400 211.570 82.720 211.630 ;
        RECT 88.380 211.570 88.700 211.630 ;
        RECT 82.400 211.430 88.700 211.570 ;
        RECT 82.400 211.370 82.720 211.430 ;
        RECT 88.380 211.370 88.700 211.430 ;
        RECT 89.775 211.570 90.065 211.615 ;
        RECT 92.520 211.570 92.840 211.630 ;
        RECT 89.775 211.430 92.840 211.570 ;
        RECT 89.775 211.385 90.065 211.430 ;
        RECT 92.520 211.370 92.840 211.430 ;
        RECT 94.360 211.570 94.680 211.630 ;
        RECT 108.160 211.570 108.480 211.630 ;
        RECT 94.360 211.430 108.480 211.570 ;
        RECT 94.360 211.370 94.680 211.430 ;
        RECT 108.160 211.370 108.480 211.430 ;
        RECT 116.440 211.570 116.760 211.630 ;
        RECT 124.720 211.570 125.040 211.630 ;
        RECT 125.655 211.570 125.945 211.615 ;
        RECT 116.440 211.430 125.945 211.570 ;
        RECT 116.440 211.370 116.760 211.430 ;
        RECT 124.720 211.370 125.040 211.430 ;
        RECT 125.655 211.385 125.945 211.430 ;
        RECT 133.920 211.570 134.240 211.630 ;
        RECT 135.315 211.570 135.605 211.615 ;
        RECT 135.760 211.570 136.080 211.630 ;
        RECT 133.920 211.430 135.070 211.570 ;
        RECT 133.920 211.370 134.240 211.430 ;
        RECT 64.000 211.230 64.320 211.290 ;
        RECT 64.920 211.230 65.240 211.290 ;
        RECT 50.200 210.750 52.730 210.890 ;
        RECT 53.050 211.090 62.390 211.230 ;
        RECT 50.200 210.690 50.520 210.750 ;
        RECT 51.135 210.705 51.425 210.750 ;
        RECT 53.050 210.550 53.190 211.090 ;
        RECT 53.435 210.890 53.725 210.935 ;
        RECT 54.800 210.890 55.120 210.950 ;
        RECT 53.435 210.750 55.120 210.890 ;
        RECT 53.435 210.705 53.725 210.750 ;
        RECT 54.800 210.690 55.120 210.750 ;
        RECT 55.720 210.890 56.040 210.950 ;
        RECT 56.655 210.890 56.945 210.935 ;
        RECT 55.720 210.750 56.945 210.890 ;
        RECT 55.720 210.690 56.040 210.750 ;
        RECT 56.655 210.705 56.945 210.750 ;
        RECT 58.020 210.890 58.340 210.950 ;
        RECT 59.415 210.890 59.705 210.935 ;
        RECT 59.860 210.890 60.180 210.950 ;
        RECT 58.020 210.750 60.180 210.890 ;
        RECT 58.020 210.690 58.340 210.750 ;
        RECT 59.415 210.705 59.705 210.750 ;
        RECT 59.860 210.690 60.180 210.750 ;
        RECT 61.240 210.690 61.560 210.950 ;
        RECT 62.250 210.935 62.390 211.090 ;
        RECT 64.000 211.090 65.240 211.230 ;
        RECT 64.000 211.030 64.320 211.090 ;
        RECT 64.920 211.030 65.240 211.090 ;
        RECT 65.380 211.230 65.700 211.290 ;
        RECT 74.120 211.230 74.440 211.290 ;
        RECT 86.540 211.230 86.860 211.290 ;
        RECT 92.060 211.230 92.380 211.290 ;
        RECT 95.740 211.230 96.060 211.290 ;
        RECT 107.700 211.230 108.020 211.290 ;
        RECT 65.380 211.090 90.450 211.230 ;
        RECT 65.380 211.030 65.700 211.090 ;
        RECT 74.120 211.030 74.440 211.090 ;
        RECT 86.540 211.030 86.860 211.090 ;
        RECT 62.175 210.705 62.465 210.935 ;
        RECT 77.800 210.890 78.120 210.950 ;
        RECT 85.160 210.890 85.480 210.950 ;
        RECT 77.800 210.750 85.480 210.890 ;
        RECT 77.800 210.690 78.120 210.750 ;
        RECT 85.160 210.690 85.480 210.750 ;
        RECT 87.460 210.890 87.780 210.950 ;
        RECT 87.935 210.890 88.225 210.935 ;
        RECT 89.760 210.890 90.080 210.950 ;
        RECT 87.460 210.750 90.080 210.890 ;
        RECT 90.310 210.890 90.450 211.090 ;
        RECT 92.060 211.090 94.130 211.230 ;
        RECT 92.060 211.030 92.380 211.090 ;
        RECT 93.990 210.935 94.130 211.090 ;
        RECT 95.740 211.090 108.020 211.230 ;
        RECT 95.740 211.030 96.060 211.090 ;
        RECT 107.700 211.030 108.020 211.090 ;
        RECT 111.380 211.230 111.700 211.290 ;
        RECT 114.615 211.230 114.905 211.275 ;
        RECT 111.380 211.090 114.905 211.230 ;
        RECT 111.380 211.030 111.700 211.090 ;
        RECT 114.615 211.045 114.905 211.090 ;
        RECT 115.075 211.230 115.365 211.275 ;
        RECT 120.595 211.230 120.885 211.275 ;
        RECT 115.075 211.090 115.875 211.230 ;
        RECT 115.075 211.045 115.365 211.090 ;
        RECT 91.315 210.890 91.605 210.935 ;
        RECT 92.995 210.890 93.285 210.935 ;
        RECT 90.310 210.750 91.605 210.890 ;
        RECT 87.460 210.690 87.780 210.750 ;
        RECT 87.935 210.705 88.225 210.750 ;
        RECT 89.760 210.690 90.080 210.750 ;
        RECT 91.315 210.705 91.605 210.750 ;
        RECT 92.150 210.750 93.285 210.890 ;
        RECT 48.220 210.410 53.190 210.550 ;
        RECT 57.100 210.350 57.420 210.610 ;
        RECT 57.560 210.350 57.880 210.610 ;
        RECT 58.940 210.550 59.260 210.610 ;
        RECT 62.620 210.550 62.940 210.610 ;
        RECT 58.940 210.410 62.940 210.550 ;
        RECT 58.940 210.350 59.260 210.410 ;
        RECT 62.620 210.350 62.940 210.410 ;
        RECT 63.080 210.550 63.400 210.610 ;
        RECT 82.400 210.550 82.720 210.610 ;
        RECT 63.080 210.410 82.720 210.550 ;
        RECT 63.080 210.350 63.400 210.410 ;
        RECT 82.400 210.350 82.720 210.410 ;
        RECT 88.395 210.550 88.685 210.595 ;
        RECT 89.300 210.550 89.620 210.610 ;
        RECT 88.395 210.410 89.620 210.550 ;
        RECT 88.395 210.365 88.685 210.410 ;
        RECT 89.300 210.350 89.620 210.410 ;
        RECT 90.235 210.550 90.525 210.595 ;
        RECT 90.680 210.550 91.000 210.610 ;
        RECT 90.235 210.410 91.000 210.550 ;
        RECT 90.235 210.365 90.525 210.410 ;
        RECT 90.680 210.350 91.000 210.410 ;
        RECT 47.440 210.210 47.760 210.270 ;
        RECT 47.070 210.070 47.760 210.210 ;
        RECT 40.965 210.025 41.255 210.070 ;
        RECT 42.855 210.025 43.145 210.070 ;
        RECT 45.975 210.025 46.265 210.070 ;
        RECT 47.440 210.010 47.760 210.070 ;
        RECT 48.835 210.210 49.125 210.255 ;
        RECT 51.120 210.210 51.440 210.270 ;
        RECT 72.740 210.210 73.060 210.270 ;
        RECT 48.835 210.070 50.890 210.210 ;
        RECT 48.835 210.025 49.125 210.070 ;
        RECT 4.660 209.730 12.250 209.870 ;
        RECT 13.400 209.870 13.720 209.930 ;
        RECT 19.840 209.870 20.160 209.930 ;
        RECT 13.400 209.730 20.160 209.870 ;
        RECT 4.660 209.670 4.980 209.730 ;
        RECT 13.400 209.670 13.720 209.730 ;
        RECT 19.840 209.670 20.160 209.730 ;
        RECT 26.740 209.915 27.060 209.930 ;
        RECT 26.740 209.685 27.275 209.915 ;
        RECT 34.560 209.870 34.880 209.930 ;
        RECT 50.215 209.870 50.505 209.915 ;
        RECT 34.560 209.730 50.505 209.870 ;
        RECT 50.750 209.870 50.890 210.070 ;
        RECT 51.120 210.070 73.060 210.210 ;
        RECT 51.120 210.010 51.440 210.070 ;
        RECT 72.740 210.010 73.060 210.070 ;
        RECT 87.460 210.210 87.780 210.270 ;
        RECT 92.150 210.210 92.290 210.750 ;
        RECT 92.995 210.705 93.285 210.750 ;
        RECT 93.915 210.705 94.205 210.935 ;
        RECT 92.535 210.365 92.825 210.595 ;
        RECT 93.070 210.550 93.210 210.705 ;
        RECT 94.360 210.690 94.680 210.950 ;
        RECT 94.835 210.890 95.125 210.935 ;
        RECT 96.660 210.890 96.980 210.950 ;
        RECT 94.835 210.750 96.980 210.890 ;
        RECT 94.835 210.705 95.125 210.750 ;
        RECT 96.660 210.690 96.980 210.750 ;
        RECT 97.120 210.690 97.440 210.950 ;
        RECT 97.580 210.890 97.900 210.950 ;
        RECT 98.055 210.890 98.345 210.935 ;
        RECT 97.580 210.750 98.345 210.890 ;
        RECT 97.580 210.690 97.900 210.750 ;
        RECT 98.055 210.705 98.345 210.750 ;
        RECT 99.435 210.890 99.725 210.935 ;
        RECT 99.435 210.750 100.110 210.890 ;
        RECT 99.435 210.705 99.725 210.750 ;
        RECT 97.210 210.550 97.350 210.690 ;
        RECT 93.070 210.410 97.350 210.550 ;
        RECT 98.130 210.550 98.270 210.705 ;
        RECT 99.970 210.550 100.110 210.750 ;
        RECT 100.340 210.690 100.660 210.950 ;
        RECT 103.560 210.890 103.880 210.950 ;
        RECT 105.860 210.890 106.180 210.950 ;
        RECT 103.560 210.750 106.180 210.890 ;
        RECT 103.560 210.690 103.880 210.750 ;
        RECT 105.860 210.690 106.180 210.750 ;
        RECT 107.240 210.890 107.560 210.950 ;
        RECT 109.540 210.890 109.860 210.950 ;
        RECT 107.240 210.750 111.610 210.890 ;
        RECT 107.240 210.690 107.560 210.750 ;
        RECT 109.540 210.690 109.860 210.750 ;
        RECT 104.480 210.550 104.800 210.610 ;
        RECT 110.460 210.550 110.780 210.610 ;
        RECT 98.130 210.410 99.650 210.550 ;
        RECT 99.970 210.410 104.800 210.550 ;
        RECT 87.460 210.070 92.290 210.210 ;
        RECT 92.610 210.210 92.750 210.365 ;
        RECT 98.515 210.210 98.805 210.255 ;
        RECT 92.610 210.070 98.805 210.210 ;
        RECT 87.460 210.010 87.780 210.070 ;
        RECT 98.515 210.025 98.805 210.070 ;
        RECT 98.960 210.010 99.280 210.270 ;
        RECT 99.510 210.210 99.650 210.410 ;
        RECT 104.480 210.350 104.800 210.410 ;
        RECT 105.030 210.410 110.780 210.550 ;
        RECT 105.030 210.210 105.170 210.410 ;
        RECT 110.460 210.350 110.780 210.410 ;
        RECT 110.920 210.350 111.240 210.610 ;
        RECT 111.470 210.595 111.610 210.750 ;
        RECT 111.840 210.690 112.160 210.950 ;
        RECT 115.735 210.890 115.875 211.090 ;
        RECT 116.530 211.090 120.885 211.230 ;
        RECT 116.530 210.890 116.670 211.090 ;
        RECT 120.595 211.045 120.885 211.090 ;
        RECT 121.960 211.230 122.280 211.290 ;
        RECT 122.435 211.230 122.725 211.275 ;
        RECT 123.340 211.230 123.660 211.290 ;
        RECT 133.460 211.230 133.780 211.290 ;
        RECT 121.960 211.090 123.660 211.230 ;
        RECT 121.960 211.030 122.280 211.090 ;
        RECT 122.435 211.045 122.725 211.090 ;
        RECT 123.340 211.030 123.660 211.090 ;
        RECT 125.730 211.090 128.170 211.230 ;
        RECT 115.735 210.750 116.670 210.890 ;
        RECT 116.900 210.690 117.220 210.950 ;
        RECT 117.360 210.890 117.680 210.950 ;
        RECT 118.295 210.890 118.585 210.935 ;
        RECT 117.360 210.750 118.585 210.890 ;
        RECT 117.360 210.690 117.680 210.750 ;
        RECT 118.295 210.705 118.585 210.750 ;
        RECT 119.215 210.890 119.505 210.935 ;
        RECT 119.660 210.890 119.980 210.950 ;
        RECT 119.215 210.750 119.980 210.890 ;
        RECT 119.215 210.705 119.505 210.750 ;
        RECT 119.660 210.690 119.980 210.750 ;
        RECT 121.500 210.690 121.820 210.950 ;
        RECT 122.895 210.705 123.185 210.935 ;
        RECT 111.395 210.365 111.685 210.595 ;
        RECT 112.775 210.550 113.065 210.595 ;
        RECT 113.235 210.550 113.525 210.595 ;
        RECT 112.775 210.410 113.525 210.550 ;
        RECT 112.775 210.365 113.065 210.410 ;
        RECT 113.235 210.365 113.525 210.410 ;
        RECT 99.510 210.070 105.170 210.210 ;
        RECT 107.240 210.210 107.560 210.270 ;
        RECT 111.010 210.210 111.150 210.350 ;
        RECT 107.240 210.070 111.150 210.210 ;
        RECT 111.470 210.210 111.610 210.365 ;
        RECT 115.060 210.350 115.380 210.610 ;
        RECT 115.660 210.365 115.950 210.595 ;
        RECT 122.970 210.550 123.110 210.705 ;
        RECT 123.800 210.690 124.120 210.950 ;
        RECT 124.735 210.880 125.025 210.935 ;
        RECT 125.730 210.890 125.870 211.090 ;
        RECT 128.030 210.950 128.170 211.090 ;
        RECT 132.630 211.090 134.610 211.230 ;
        RECT 132.630 210.950 132.770 211.090 ;
        RECT 133.460 211.030 133.780 211.090 ;
        RECT 125.270 210.880 125.870 210.890 ;
        RECT 124.735 210.750 125.870 210.880 ;
        RECT 124.735 210.740 125.410 210.750 ;
        RECT 124.735 210.705 125.025 210.740 ;
        RECT 126.115 210.705 126.405 210.935 ;
        RECT 124.275 210.550 124.565 210.595 ;
        RECT 122.970 210.410 124.565 210.550 ;
        RECT 124.275 210.365 124.565 210.410 ;
        RECT 125.640 210.550 125.960 210.610 ;
        RECT 126.190 210.550 126.330 210.705 ;
        RECT 126.560 210.690 126.880 210.950 ;
        RECT 127.940 210.690 128.260 210.950 ;
        RECT 131.620 210.890 131.940 210.950 ;
        RECT 132.095 210.890 132.385 210.935 ;
        RECT 131.620 210.750 132.385 210.890 ;
        RECT 131.620 210.690 131.940 210.750 ;
        RECT 132.095 210.705 132.385 210.750 ;
        RECT 132.540 210.690 132.860 210.950 ;
        RECT 133.000 210.690 133.320 210.950 ;
        RECT 134.470 210.935 134.610 211.090 ;
        RECT 134.395 210.705 134.685 210.935 ;
        RECT 125.640 210.410 126.330 210.550 ;
        RECT 115.150 210.210 115.290 210.350 ;
        RECT 111.470 210.070 115.290 210.210 ;
        RECT 107.240 210.010 107.560 210.070 ;
        RECT 52.960 209.870 53.280 209.930 ;
        RECT 50.750 209.730 53.280 209.870 ;
        RECT 26.740 209.670 27.060 209.685 ;
        RECT 34.560 209.670 34.880 209.730 ;
        RECT 50.215 209.685 50.505 209.730 ;
        RECT 52.960 209.670 53.280 209.730 ;
        RECT 54.800 209.670 55.120 209.930 ;
        RECT 55.260 209.870 55.580 209.930 ;
        RECT 70.900 209.870 71.220 209.930 ;
        RECT 81.940 209.870 82.260 209.930 ;
        RECT 55.260 209.730 82.260 209.870 ;
        RECT 55.260 209.670 55.580 209.730 ;
        RECT 70.900 209.670 71.220 209.730 ;
        RECT 81.940 209.670 82.260 209.730 ;
        RECT 87.000 209.870 87.320 209.930 ;
        RECT 87.935 209.870 88.225 209.915 ;
        RECT 87.000 209.730 88.225 209.870 ;
        RECT 87.000 209.670 87.320 209.730 ;
        RECT 87.935 209.685 88.225 209.730 ;
        RECT 89.300 209.870 89.620 209.930 ;
        RECT 90.695 209.870 90.985 209.915 ;
        RECT 89.300 209.730 90.985 209.870 ;
        RECT 89.300 209.670 89.620 209.730 ;
        RECT 90.695 209.685 90.985 209.730 ;
        RECT 92.520 209.870 92.840 209.930 ;
        RECT 96.215 209.870 96.505 209.915 ;
        RECT 92.520 209.730 96.505 209.870 ;
        RECT 92.520 209.670 92.840 209.730 ;
        RECT 96.215 209.685 96.505 209.730 ;
        RECT 96.675 209.870 96.965 209.915 ;
        RECT 104.020 209.870 104.340 209.930 ;
        RECT 96.675 209.730 104.340 209.870 ;
        RECT 96.675 209.685 96.965 209.730 ;
        RECT 104.020 209.670 104.340 209.730 ;
        RECT 104.480 209.870 104.800 209.930 ;
        RECT 115.735 209.870 115.875 210.365 ;
        RECT 125.640 210.350 125.960 210.410 ;
        RECT 133.920 210.350 134.240 210.610 ;
        RECT 134.930 210.550 135.070 211.430 ;
        RECT 135.315 211.430 136.080 211.570 ;
        RECT 135.315 211.385 135.605 211.430 ;
        RECT 135.760 211.370 136.080 211.430 ;
        RECT 145.880 211.370 146.200 211.630 ;
        RECT 147.260 211.370 147.580 211.630 ;
        RECT 153.700 211.570 154.020 211.630 ;
        RECT 147.810 211.430 154.020 211.570 ;
        RECT 145.970 211.230 146.110 211.370 ;
        RECT 139.530 211.090 146.110 211.230 ;
        RECT 137.140 210.890 137.460 210.950 ;
        RECT 139.530 210.935 139.670 211.090 ;
        RECT 139.455 210.890 139.745 210.935 ;
        RECT 137.140 210.750 139.745 210.890 ;
        RECT 137.140 210.690 137.460 210.750 ;
        RECT 139.455 210.705 139.745 210.750 ;
        RECT 140.360 210.690 140.680 210.950 ;
        RECT 140.835 210.890 141.125 210.935 ;
        RECT 147.350 210.890 147.490 211.370 ;
        RECT 140.835 210.750 147.490 210.890 ;
        RECT 140.835 210.705 141.125 210.750 ;
        RECT 147.810 210.550 147.950 211.430 ;
        RECT 153.700 211.370 154.020 211.430 ;
        RECT 148.640 211.230 148.960 211.290 ;
        RECT 153.255 211.230 153.545 211.275 ;
        RECT 155.080 211.230 155.400 211.290 ;
        RECT 148.640 211.090 155.400 211.230 ;
        RECT 148.640 211.030 148.960 211.090 ;
        RECT 153.255 211.045 153.545 211.090 ;
        RECT 155.080 211.030 155.400 211.090 ;
        RECT 151.875 210.705 152.165 210.935 ;
        RECT 134.930 210.410 147.950 210.550 ;
        RECT 151.950 210.550 152.090 210.705 ;
        RECT 152.320 210.690 152.640 210.950 ;
        RECT 153.700 210.690 154.020 210.950 ;
        RECT 153.790 210.550 153.930 210.690 ;
        RECT 151.950 210.410 153.930 210.550 ;
        RECT 116.455 210.210 116.745 210.255 ;
        RECT 133.475 210.210 133.765 210.255 ;
        RECT 116.455 210.070 133.765 210.210 ;
        RECT 116.455 210.025 116.745 210.070 ;
        RECT 133.475 210.025 133.765 210.070 ;
        RECT 139.915 210.210 140.205 210.255 ;
        RECT 140.360 210.210 140.680 210.270 ;
        RECT 142.660 210.210 142.980 210.270 ;
        RECT 139.915 210.070 142.980 210.210 ;
        RECT 139.915 210.025 140.205 210.070 ;
        RECT 140.360 210.010 140.680 210.070 ;
        RECT 142.660 210.010 142.980 210.070 ;
        RECT 104.480 209.730 115.875 209.870 ;
        RECT 104.480 209.670 104.800 209.730 ;
        RECT 117.820 209.670 118.140 209.930 ;
        RECT 118.740 209.870 119.060 209.930 ;
        RECT 120.135 209.870 120.425 209.915 ;
        RECT 118.740 209.730 120.425 209.870 ;
        RECT 118.740 209.670 119.060 209.730 ;
        RECT 120.135 209.685 120.425 209.730 ;
        RECT 130.240 209.870 130.560 209.930 ;
        RECT 138.535 209.870 138.825 209.915 ;
        RECT 130.240 209.730 138.825 209.870 ;
        RECT 130.240 209.670 130.560 209.730 ;
        RECT 138.535 209.685 138.825 209.730 ;
        RECT 2.750 209.050 158.230 209.530 ;
        RECT 4.660 208.650 4.980 208.910 ;
        RECT 15.240 208.650 15.560 208.910 ;
        RECT 17.095 208.665 17.385 208.895 ;
        RECT 45.140 208.850 45.460 208.910 ;
        RECT 50.200 208.850 50.520 208.910 ;
        RECT 30.050 208.710 43.070 208.850 ;
        RECT 4.215 208.170 4.505 208.215 ;
        RECT 4.750 208.170 4.890 208.650 ;
        RECT 5.085 208.510 5.375 208.555 ;
        RECT 6.975 208.510 7.265 208.555 ;
        RECT 10.095 208.510 10.385 208.555 ;
        RECT 5.085 208.370 10.385 208.510 ;
        RECT 5.085 208.325 5.375 208.370 ;
        RECT 6.975 208.325 7.265 208.370 ;
        RECT 10.095 208.325 10.385 208.370 ;
        RECT 4.215 208.030 4.890 208.170 ;
        RECT 17.170 208.170 17.310 208.665 ;
        RECT 20.775 208.170 21.065 208.215 ;
        RECT 17.170 208.030 21.065 208.170 ;
        RECT 4.215 207.985 4.505 208.030 ;
        RECT 20.775 207.985 21.065 208.030 ;
        RECT 4.680 207.830 4.970 207.875 ;
        RECT 6.515 207.830 6.805 207.875 ;
        RECT 10.095 207.830 10.385 207.875 ;
        RECT 4.680 207.690 10.385 207.830 ;
        RECT 4.680 207.645 4.970 207.690 ;
        RECT 6.515 207.645 6.805 207.690 ;
        RECT 10.095 207.645 10.385 207.690 ;
        RECT 11.175 207.830 11.465 207.850 ;
        RECT 13.400 207.830 13.720 207.890 ;
        RECT 11.175 207.690 13.720 207.830 ;
        RECT 5.580 207.290 5.900 207.550 ;
        RECT 11.175 207.535 11.465 207.690 ;
        RECT 13.400 207.630 13.720 207.690 ;
        RECT 14.335 207.830 14.625 207.875 ;
        RECT 20.850 207.830 20.990 207.985 ;
        RECT 21.680 207.970 22.000 208.230 ;
        RECT 23.060 208.170 23.380 208.230 ;
        RECT 23.535 208.170 23.825 208.215 ;
        RECT 27.675 208.170 27.965 208.215 ;
        RECT 30.050 208.170 30.190 208.710 ;
        RECT 30.435 208.325 30.725 208.555 ;
        RECT 23.060 208.030 30.190 208.170 ;
        RECT 23.060 207.970 23.380 208.030 ;
        RECT 23.535 207.985 23.825 208.030 ;
        RECT 27.675 207.985 27.965 208.030 ;
        RECT 26.740 207.830 27.060 207.890 ;
        RECT 29.960 207.830 30.280 207.890 ;
        RECT 14.335 207.690 18.230 207.830 ;
        RECT 20.850 207.690 30.280 207.830 ;
        RECT 30.510 207.830 30.650 208.325 ;
        RECT 39.620 208.310 39.940 208.570 ;
        RECT 42.930 208.510 43.070 208.710 ;
        RECT 45.140 208.710 50.520 208.850 ;
        RECT 45.140 208.650 45.460 208.710 ;
        RECT 50.200 208.650 50.520 208.710 ;
        RECT 50.675 208.850 50.965 208.895 ;
        RECT 51.120 208.850 51.440 208.910 ;
        RECT 50.675 208.710 51.440 208.850 ;
        RECT 50.675 208.665 50.965 208.710 ;
        RECT 51.120 208.650 51.440 208.710 ;
        RECT 53.420 208.650 53.740 208.910 ;
        RECT 57.100 208.850 57.420 208.910 ;
        RECT 64.000 208.850 64.320 208.910 ;
        RECT 68.140 208.850 68.460 208.910 ;
        RECT 57.100 208.710 64.320 208.850 ;
        RECT 57.100 208.650 57.420 208.710 ;
        RECT 64.000 208.650 64.320 208.710 ;
        RECT 65.470 208.710 68.460 208.850 ;
        RECT 47.915 208.510 48.205 208.555 ;
        RECT 65.470 208.510 65.610 208.710 ;
        RECT 68.140 208.650 68.460 208.710 ;
        RECT 71.375 208.665 71.665 208.895 ;
        RECT 71.820 208.850 72.140 208.910 ;
        RECT 72.755 208.850 73.045 208.895 ;
        RECT 71.820 208.710 73.045 208.850 ;
        RECT 42.930 208.370 43.990 208.510 ;
        RECT 31.340 208.170 31.660 208.230 ;
        RECT 42.930 208.215 43.070 208.370 ;
        RECT 34.115 208.170 34.405 208.215 ;
        RECT 31.340 208.030 34.405 208.170 ;
        RECT 31.340 207.970 31.660 208.030 ;
        RECT 34.115 207.985 34.405 208.030 ;
        RECT 42.855 207.985 43.145 208.215 ;
        RECT 43.850 208.170 43.990 208.370 ;
        RECT 47.915 208.370 65.610 208.510 ;
        RECT 65.855 208.510 66.145 208.555 ;
        RECT 71.450 208.510 71.590 208.665 ;
        RECT 71.820 208.650 72.140 208.710 ;
        RECT 72.755 208.665 73.045 208.710 ;
        RECT 73.215 208.850 73.505 208.895 ;
        RECT 73.660 208.850 73.980 208.910 ;
        RECT 73.215 208.710 73.980 208.850 ;
        RECT 73.215 208.665 73.505 208.710 ;
        RECT 73.660 208.650 73.980 208.710 ;
        RECT 76.420 208.650 76.740 208.910 ;
        RECT 76.880 208.850 77.200 208.910 ;
        RECT 81.035 208.850 81.325 208.895 ;
        RECT 76.880 208.710 81.325 208.850 ;
        RECT 76.880 208.650 77.200 208.710 ;
        RECT 81.035 208.665 81.325 208.710 ;
        RECT 82.400 208.850 82.720 208.910 ;
        RECT 94.360 208.850 94.680 208.910 ;
        RECT 94.835 208.850 95.125 208.895 ;
        RECT 82.400 208.710 89.530 208.850 ;
        RECT 82.400 208.650 82.720 208.710 ;
        RECT 72.280 208.510 72.600 208.570 ;
        RECT 87.460 208.510 87.780 208.570 ;
        RECT 65.855 208.370 72.600 208.510 ;
        RECT 47.915 208.325 48.205 208.370 ;
        RECT 65.855 208.325 66.145 208.370 ;
        RECT 49.740 208.170 50.060 208.230 ;
        RECT 63.080 208.170 63.400 208.230 ;
        RECT 65.930 208.170 66.070 208.325 ;
        RECT 72.280 208.310 72.600 208.370 ;
        RECT 73.750 208.370 87.780 208.510 ;
        RECT 89.390 208.510 89.530 208.710 ;
        RECT 94.360 208.710 95.125 208.850 ;
        RECT 94.360 208.650 94.680 208.710 ;
        RECT 94.835 208.665 95.125 208.710 ;
        RECT 95.280 208.850 95.600 208.910 ;
        RECT 95.755 208.850 96.045 208.895 ;
        RECT 95.280 208.710 96.045 208.850 ;
        RECT 95.280 208.650 95.600 208.710 ;
        RECT 95.755 208.665 96.045 208.710 ;
        RECT 96.675 208.850 96.965 208.895 ;
        RECT 104.480 208.850 104.800 208.910 ;
        RECT 111.380 208.850 111.700 208.910 ;
        RECT 96.675 208.710 104.800 208.850 ;
        RECT 96.675 208.665 96.965 208.710 ;
        RECT 104.480 208.650 104.800 208.710 ;
        RECT 109.630 208.710 111.700 208.850 ;
        RECT 92.980 208.510 93.300 208.570 ;
        RECT 89.390 208.370 93.300 208.510 ;
        RECT 73.750 208.170 73.890 208.370 ;
        RECT 87.460 208.310 87.780 208.370 ;
        RECT 92.980 208.310 93.300 208.370 ;
        RECT 97.120 208.510 97.440 208.570 ;
        RECT 98.040 208.510 98.360 208.570 ;
        RECT 109.630 208.510 109.770 208.710 ;
        RECT 111.380 208.650 111.700 208.710 ;
        RECT 116.900 208.850 117.220 208.910 ;
        RECT 121.975 208.850 122.265 208.895 ;
        RECT 116.900 208.710 122.265 208.850 ;
        RECT 116.900 208.650 117.220 208.710 ;
        RECT 121.975 208.665 122.265 208.710 ;
        RECT 124.260 208.650 124.580 208.910 ;
        RECT 130.715 208.665 131.005 208.895 ;
        RECT 133.000 208.850 133.320 208.910 ;
        RECT 133.475 208.850 133.765 208.895 ;
        RECT 133.000 208.710 133.765 208.850 ;
        RECT 97.120 208.370 97.810 208.510 ;
        RECT 97.120 208.310 97.440 208.370 ;
        RECT 43.850 208.030 50.060 208.170 ;
        RECT 49.740 207.970 50.060 208.030 ;
        RECT 59.030 208.030 63.400 208.170 ;
        RECT 36.860 207.830 37.180 207.890 ;
        RECT 30.510 207.690 37.180 207.830 ;
        RECT 14.335 207.645 14.625 207.690 ;
        RECT 7.875 207.490 8.525 207.535 ;
        RECT 11.175 207.490 11.765 207.535 ;
        RECT 7.875 207.350 11.765 207.490 ;
        RECT 7.875 207.305 8.525 207.350 ;
        RECT 11.475 207.305 11.765 207.350 ;
        RECT 16.160 207.290 16.480 207.550 ;
        RECT 18.090 207.490 18.230 207.690 ;
        RECT 26.740 207.630 27.060 207.690 ;
        RECT 29.960 207.630 30.280 207.690 ;
        RECT 36.860 207.630 37.180 207.690 ;
        RECT 40.080 207.830 40.400 207.890 ;
        RECT 40.555 207.830 40.845 207.875 ;
        RECT 40.080 207.690 40.845 207.830 ;
        RECT 40.080 207.630 40.400 207.690 ;
        RECT 40.555 207.645 40.845 207.690 ;
        RECT 43.775 207.830 44.065 207.875 ;
        RECT 52.960 207.830 53.280 207.890 ;
        RECT 43.775 207.690 53.280 207.830 ;
        RECT 43.775 207.645 44.065 207.690 ;
        RECT 52.960 207.630 53.280 207.690 ;
        RECT 53.895 207.830 54.185 207.875 ;
        RECT 54.800 207.830 55.120 207.890 ;
        RECT 53.895 207.690 55.120 207.830 ;
        RECT 53.895 207.645 54.185 207.690 ;
        RECT 54.800 207.630 55.120 207.690 ;
        RECT 57.100 207.630 57.420 207.890 ;
        RECT 57.575 207.830 57.865 207.875 ;
        RECT 59.030 207.830 59.170 208.030 ;
        RECT 63.080 207.970 63.400 208.030 ;
        RECT 63.630 208.030 66.070 208.170 ;
        RECT 71.450 208.030 73.890 208.170 ;
        RECT 74.135 208.170 74.425 208.215 ;
        RECT 81.940 208.170 82.260 208.230 ;
        RECT 74.135 208.030 82.260 208.170 ;
        RECT 57.575 207.690 59.170 207.830 ;
        RECT 57.575 207.645 57.865 207.690 ;
        RECT 59.400 207.630 59.720 207.890 ;
        RECT 63.630 207.875 63.770 208.030 ;
        RECT 62.175 207.645 62.465 207.875 ;
        RECT 63.555 207.830 63.845 207.875 ;
        RECT 63.445 207.690 63.845 207.830 ;
        RECT 63.555 207.645 63.845 207.690 ;
        RECT 27.200 207.490 27.520 207.550 ;
        RECT 18.090 207.350 18.690 207.490 ;
        RECT 12.940 206.950 13.260 207.210 ;
        RECT 16.620 207.150 16.940 207.210 ;
        RECT 17.175 207.150 17.465 207.195 ;
        RECT 16.620 207.010 17.465 207.150 ;
        RECT 16.620 206.950 16.940 207.010 ;
        RECT 17.175 206.965 17.465 207.010 ;
        RECT 18.000 206.950 18.320 207.210 ;
        RECT 18.550 207.195 18.690 207.350 ;
        RECT 24.530 207.350 26.970 207.490 ;
        RECT 24.530 207.210 24.670 207.350 ;
        RECT 26.830 207.210 26.970 207.350 ;
        RECT 27.200 207.350 31.570 207.490 ;
        RECT 27.200 207.290 27.520 207.350 ;
        RECT 18.475 206.965 18.765 207.195 ;
        RECT 20.300 206.950 20.620 207.210 ;
        RECT 23.980 206.950 24.300 207.210 ;
        RECT 24.440 206.950 24.760 207.210 ;
        RECT 26.280 206.950 26.600 207.210 ;
        RECT 26.740 206.950 27.060 207.210 ;
        RECT 28.120 206.950 28.440 207.210 ;
        RECT 28.595 207.150 28.885 207.195 ;
        RECT 29.960 207.150 30.280 207.210 ;
        RECT 31.430 207.195 31.570 207.350 ;
        RECT 33.180 207.290 33.500 207.550 ;
        RECT 37.795 207.490 38.085 207.535 ;
        RECT 39.620 207.490 39.940 207.550 ;
        RECT 45.140 207.490 45.460 207.550 ;
        RECT 46.535 207.490 46.825 207.535 ;
        RECT 37.795 207.350 45.460 207.490 ;
        RECT 37.795 207.305 38.085 207.350 ;
        RECT 39.620 207.290 39.940 207.350 ;
        RECT 45.140 207.290 45.460 207.350 ;
        RECT 45.690 207.350 46.825 207.490 ;
        RECT 28.595 207.010 30.280 207.150 ;
        RECT 28.595 206.965 28.885 207.010 ;
        RECT 29.960 206.950 30.280 207.010 ;
        RECT 31.355 206.965 31.645 207.195 ;
        RECT 32.720 207.150 33.040 207.210 ;
        RECT 33.655 207.150 33.945 207.195 ;
        RECT 32.720 207.010 33.945 207.150 ;
        RECT 32.720 206.950 33.040 207.010 ;
        RECT 33.655 206.965 33.945 207.010 ;
        RECT 37.320 206.950 37.640 207.210 ;
        RECT 43.300 206.950 43.620 207.210 ;
        RECT 45.690 207.195 45.830 207.350 ;
        RECT 46.535 207.305 46.825 207.350 ;
        RECT 49.280 207.290 49.600 207.550 ;
        RECT 58.020 207.290 58.340 207.550 ;
        RECT 58.725 207.490 59.015 207.535 ;
        RECT 61.255 207.490 61.545 207.535 ;
        RECT 58.725 207.350 61.545 207.490 ;
        RECT 58.725 207.305 59.015 207.350 ;
        RECT 61.255 207.305 61.545 207.350 ;
        RECT 45.615 206.965 45.905 207.195 ;
        RECT 56.180 206.950 56.500 207.210 ;
        RECT 62.250 207.150 62.390 207.645 ;
        RECT 64.920 207.630 65.240 207.890 ;
        RECT 65.855 207.830 66.145 207.875 ;
        RECT 68.140 207.830 68.460 207.890 ;
        RECT 65.855 207.690 68.460 207.830 ;
        RECT 65.855 207.645 66.145 207.690 ;
        RECT 68.140 207.630 68.460 207.690 ;
        RECT 69.520 207.630 69.840 207.890 ;
        RECT 69.995 207.830 70.285 207.875 ;
        RECT 71.450 207.830 71.590 208.030 ;
        RECT 74.135 207.985 74.425 208.030 ;
        RECT 81.940 207.970 82.260 208.030 ;
        RECT 85.620 208.170 85.940 208.230 ;
        RECT 92.060 208.170 92.380 208.230 ;
        RECT 97.670 208.170 97.810 208.370 ;
        RECT 98.040 208.370 109.770 208.510 ;
        RECT 98.040 208.310 98.360 208.370 ;
        RECT 103.560 208.170 103.880 208.230 ;
        RECT 85.620 208.030 97.350 208.170 ;
        RECT 97.670 208.030 101.030 208.170 ;
        RECT 85.620 207.970 85.940 208.030 ;
        RECT 69.995 207.690 71.590 207.830 ;
        RECT 69.995 207.645 70.285 207.690 ;
        RECT 71.820 207.630 72.140 207.890 ;
        RECT 73.200 207.830 73.520 207.890 ;
        RECT 74.595 207.830 74.885 207.875 ;
        RECT 73.200 207.690 74.885 207.830 ;
        RECT 73.200 207.630 73.520 207.690 ;
        RECT 74.595 207.645 74.885 207.690 ;
        RECT 75.055 207.645 75.345 207.875 ;
        RECT 75.515 207.830 75.805 207.875 ;
        RECT 76.420 207.830 76.740 207.890 ;
        RECT 75.515 207.690 76.740 207.830 ;
        RECT 75.515 207.645 75.805 207.690 ;
        RECT 63.095 207.490 63.385 207.535 ;
        RECT 68.600 207.490 68.920 207.550 ;
        RECT 63.095 207.350 68.920 207.490 ;
        RECT 63.095 207.305 63.385 207.350 ;
        RECT 68.600 207.290 68.920 207.350 ;
        RECT 69.060 207.150 69.380 207.210 ;
        RECT 62.250 207.010 69.380 207.150 ;
        RECT 73.290 207.150 73.430 207.630 ;
        RECT 73.660 207.490 73.980 207.550 ;
        RECT 75.130 207.490 75.270 207.645 ;
        RECT 76.420 207.630 76.740 207.690 ;
        RECT 77.340 207.630 77.660 207.890 ;
        RECT 77.800 207.630 78.120 207.890 ;
        RECT 78.275 207.645 78.565 207.875 ;
        RECT 78.735 207.645 79.025 207.875 ;
        RECT 82.415 207.645 82.705 207.875 ;
        RECT 73.660 207.350 75.270 207.490 ;
        RECT 75.960 207.490 76.280 207.550 ;
        RECT 78.350 207.490 78.490 207.645 ;
        RECT 75.960 207.350 78.490 207.490 ;
        RECT 78.810 207.490 78.950 207.645 ;
        RECT 81.940 207.490 82.260 207.550 ;
        RECT 78.810 207.350 82.260 207.490 ;
        RECT 73.660 207.290 73.980 207.350 ;
        RECT 75.960 207.290 76.280 207.350 ;
        RECT 81.940 207.290 82.260 207.350 ;
        RECT 82.490 207.150 82.630 207.645 ;
        RECT 82.860 207.630 83.180 207.890 ;
        RECT 83.335 207.830 83.625 207.875 ;
        RECT 84.240 207.830 84.560 207.890 ;
        RECT 83.335 207.690 84.560 207.830 ;
        RECT 83.335 207.645 83.625 207.690 ;
        RECT 84.240 207.630 84.560 207.690 ;
        RECT 84.700 207.630 85.020 207.890 ;
        RECT 85.175 207.645 85.465 207.875 ;
        RECT 82.860 207.150 83.180 207.210 ;
        RECT 73.290 207.010 83.180 207.150 ;
        RECT 85.250 207.150 85.390 207.645 ;
        RECT 86.080 207.630 86.400 207.890 ;
        RECT 86.630 207.875 86.770 208.030 ;
        RECT 92.060 207.970 92.380 208.030 ;
        RECT 86.555 207.645 86.845 207.875 ;
        RECT 87.015 207.830 87.305 207.875 ;
        RECT 87.460 207.830 87.780 207.890 ;
        RECT 87.015 207.690 87.780 207.830 ;
        RECT 87.015 207.645 87.305 207.690 ;
        RECT 87.460 207.630 87.780 207.690 ;
        RECT 88.380 207.830 88.700 207.890 ;
        RECT 94.820 207.830 95.140 207.890 ;
        RECT 88.380 207.690 95.140 207.830 ;
        RECT 88.380 207.630 88.700 207.690 ;
        RECT 94.820 207.630 95.140 207.690 ;
        RECT 95.280 207.830 95.600 207.890 ;
        RECT 97.210 207.875 97.350 208.030 ;
        RECT 96.215 207.830 96.505 207.875 ;
        RECT 95.280 207.690 96.505 207.830 ;
        RECT 95.280 207.630 95.600 207.690 ;
        RECT 96.215 207.645 96.505 207.690 ;
        RECT 97.135 207.830 97.425 207.875 ;
        RECT 97.135 207.690 98.730 207.830 ;
        RECT 97.135 207.645 97.425 207.690 ;
        RECT 98.590 207.550 98.730 207.690 ;
        RECT 88.840 207.490 89.160 207.550 ;
        RECT 87.550 207.350 89.160 207.490 ;
        RECT 87.550 207.150 87.690 207.350 ;
        RECT 88.840 207.290 89.160 207.350 ;
        RECT 92.980 207.490 93.300 207.550 ;
        RECT 93.915 207.490 94.205 207.535 ;
        RECT 92.980 207.350 94.205 207.490 ;
        RECT 92.980 207.290 93.300 207.350 ;
        RECT 93.915 207.305 94.205 207.350 ;
        RECT 94.450 207.350 98.275 207.490 ;
        RECT 85.250 207.010 87.690 207.150 ;
        RECT 87.935 207.150 88.225 207.195 ;
        RECT 88.380 207.150 88.700 207.210 ;
        RECT 87.935 207.010 88.700 207.150 ;
        RECT 69.060 206.950 69.380 207.010 ;
        RECT 82.860 206.950 83.180 207.010 ;
        RECT 87.935 206.965 88.225 207.010 ;
        RECT 88.380 206.950 88.700 207.010 ;
        RECT 89.300 207.150 89.620 207.210 ;
        RECT 94.450 207.150 94.590 207.350 ;
        RECT 89.300 207.010 94.590 207.150 ;
        RECT 94.965 207.150 95.255 207.195 ;
        RECT 97.120 207.150 97.440 207.210 ;
        RECT 94.965 207.010 97.440 207.150 ;
        RECT 98.135 207.150 98.275 207.350 ;
        RECT 98.500 207.290 98.820 207.550 ;
        RECT 100.890 207.210 101.030 208.030 ;
        RECT 101.350 208.030 103.880 208.170 ;
        RECT 101.350 207.875 101.490 208.030 ;
        RECT 103.560 207.970 103.880 208.030 ;
        RECT 107.255 207.985 107.545 208.215 ;
        RECT 101.275 207.645 101.565 207.875 ;
        RECT 101.720 207.630 102.040 207.890 ;
        RECT 102.180 207.630 102.500 207.890 ;
        RECT 102.655 207.830 102.945 207.875 ;
        RECT 103.100 207.830 103.420 207.890 ;
        RECT 102.655 207.690 103.420 207.830 ;
        RECT 102.655 207.645 102.945 207.690 ;
        RECT 103.100 207.630 103.420 207.690 ;
        RECT 103.580 207.550 103.870 207.765 ;
        RECT 104.020 207.630 104.340 207.890 ;
        RECT 104.940 207.630 105.260 207.890 ;
        RECT 105.875 207.830 106.165 207.875 ;
        RECT 107.330 207.830 107.470 207.985 ;
        RECT 108.160 207.970 108.480 208.230 ;
        RECT 109.630 208.215 109.770 208.370 ;
        RECT 110.460 208.510 110.780 208.570 ;
        RECT 123.800 208.510 124.120 208.570 ;
        RECT 125.640 208.510 125.960 208.570 ;
        RECT 110.460 208.370 125.960 208.510 ;
        RECT 110.460 208.310 110.780 208.370 ;
        RECT 123.800 208.310 124.120 208.370 ;
        RECT 125.640 208.310 125.960 208.370 ;
        RECT 130.790 208.510 130.930 208.665 ;
        RECT 133.000 208.650 133.320 208.710 ;
        RECT 133.475 208.665 133.765 208.710 ;
        RECT 147.260 208.650 147.580 208.910 ;
        RECT 149.560 208.650 149.880 208.910 ;
        RECT 154.175 208.665 154.465 208.895 ;
        RECT 137.140 208.510 137.460 208.570 ;
        RECT 130.790 208.370 137.460 208.510 ;
        RECT 109.555 207.985 109.845 208.215 ;
        RECT 110.920 208.170 111.240 208.230 ;
        RECT 111.395 208.170 111.685 208.215 ;
        RECT 110.920 208.030 111.685 208.170 ;
        RECT 110.920 207.970 111.240 208.030 ;
        RECT 111.395 207.985 111.685 208.030 ;
        RECT 111.855 208.170 112.145 208.215 ;
        RECT 113.220 208.170 113.540 208.230 ;
        RECT 111.855 208.030 113.540 208.170 ;
        RECT 111.855 207.985 112.145 208.030 ;
        RECT 113.220 207.970 113.540 208.030 ;
        RECT 115.520 207.970 115.840 208.230 ;
        RECT 119.660 208.170 119.980 208.230 ;
        RECT 121.040 208.170 121.360 208.230 ;
        RECT 130.790 208.170 130.930 208.370 ;
        RECT 137.140 208.310 137.460 208.370 ;
        RECT 144.975 208.510 145.265 208.555 ;
        RECT 145.420 208.510 145.740 208.570 ;
        RECT 144.975 208.370 145.740 208.510 ;
        RECT 147.350 208.510 147.490 208.650 ;
        RECT 151.400 208.510 151.720 208.570 ;
        RECT 154.250 208.510 154.390 208.665 ;
        RECT 147.350 208.370 154.390 208.510 ;
        RECT 144.975 208.325 145.265 208.370 ;
        RECT 145.420 208.310 145.740 208.370 ;
        RECT 151.400 208.310 151.720 208.370 ;
        RECT 119.660 208.030 130.930 208.170 ;
        RECT 136.680 208.170 137.000 208.230 ;
        RECT 154.160 208.170 154.480 208.230 ;
        RECT 155.080 208.170 155.400 208.230 ;
        RECT 136.680 208.030 153.010 208.170 ;
        RECT 119.660 207.970 119.980 208.030 ;
        RECT 121.040 207.970 121.360 208.030 ;
        RECT 136.680 207.970 137.000 208.030 ;
        RECT 105.875 207.690 107.470 207.830 ;
        RECT 105.875 207.645 106.165 207.690 ;
        RECT 103.560 207.290 103.880 207.550 ;
        RECT 105.415 207.490 105.705 207.535 ;
        RECT 108.250 207.490 108.390 207.970 ;
        RECT 108.620 207.630 108.940 207.890 ;
        RECT 109.080 207.830 109.400 207.890 ;
        RECT 112.315 207.830 112.605 207.875 ;
        RECT 109.080 207.690 112.605 207.830 ;
        RECT 109.080 207.630 109.400 207.690 ;
        RECT 112.315 207.645 112.605 207.690 ;
        RECT 110.920 207.490 111.240 207.550 ;
        RECT 105.415 207.350 107.930 207.490 ;
        RECT 108.250 207.350 111.240 207.490 ;
        RECT 112.390 207.490 112.530 207.645 ;
        RECT 112.760 207.630 113.080 207.890 ;
        RECT 115.075 207.830 115.365 207.875 ;
        RECT 115.980 207.830 116.300 207.890 ;
        RECT 115.075 207.690 116.300 207.830 ;
        RECT 115.075 207.645 115.365 207.690 ;
        RECT 115.980 207.630 116.300 207.690 ;
        RECT 117.375 207.830 117.665 207.875 ;
        RECT 118.280 207.830 118.600 207.890 ;
        RECT 117.375 207.690 118.600 207.830 ;
        RECT 117.375 207.645 117.665 207.690 ;
        RECT 118.280 207.630 118.600 207.690 ;
        RECT 119.200 207.630 119.520 207.890 ;
        RECT 120.135 207.645 120.425 207.875 ;
        RECT 122.895 207.645 123.185 207.875 ;
        RECT 113.220 207.490 113.540 207.550 ;
        RECT 115.520 207.490 115.840 207.550 ;
        RECT 120.210 207.490 120.350 207.645 ;
        RECT 112.390 207.350 113.540 207.490 ;
        RECT 105.415 207.305 105.705 207.350 ;
        RECT 98.960 207.150 99.280 207.210 ;
        RECT 98.135 207.010 99.280 207.150 ;
        RECT 89.300 206.950 89.620 207.010 ;
        RECT 94.965 206.965 95.255 207.010 ;
        RECT 97.120 206.950 97.440 207.010 ;
        RECT 98.960 206.950 99.280 207.010 ;
        RECT 100.340 206.950 100.660 207.210 ;
        RECT 100.800 206.950 101.120 207.210 ;
        RECT 101.720 207.150 102.040 207.210 ;
        RECT 106.795 207.150 107.085 207.195 ;
        RECT 101.720 207.010 107.085 207.150 ;
        RECT 107.790 207.150 107.930 207.350 ;
        RECT 110.920 207.290 111.240 207.350 ;
        RECT 113.220 207.290 113.540 207.350 ;
        RECT 113.770 207.350 114.830 207.490 ;
        RECT 110.475 207.150 110.765 207.195 ;
        RECT 107.790 207.010 110.765 207.150 ;
        RECT 101.720 206.950 102.040 207.010 ;
        RECT 106.795 206.965 107.085 207.010 ;
        RECT 110.475 206.965 110.765 207.010 ;
        RECT 111.840 207.150 112.160 207.210 ;
        RECT 113.770 207.150 113.910 207.350 ;
        RECT 111.840 207.010 113.910 207.150 ;
        RECT 111.840 206.950 112.160 207.010 ;
        RECT 114.140 206.950 114.460 207.210 ;
        RECT 114.690 207.150 114.830 207.350 ;
        RECT 115.520 207.350 120.350 207.490 ;
        RECT 122.970 207.490 123.110 207.645 ;
        RECT 123.340 207.630 123.660 207.890 ;
        RECT 124.735 207.830 125.025 207.875 ;
        RECT 129.320 207.830 129.640 207.890 ;
        RECT 124.735 207.690 129.640 207.830 ;
        RECT 124.735 207.645 125.025 207.690 ;
        RECT 129.320 207.630 129.640 207.690 ;
        RECT 130.240 207.630 130.560 207.890 ;
        RECT 131.635 207.645 131.925 207.875 ;
        RECT 130.330 207.490 130.470 207.630 ;
        RECT 122.970 207.350 130.470 207.490 ;
        RECT 115.520 207.290 115.840 207.350 ;
        RECT 130.700 207.290 131.020 207.550 ;
        RECT 115.995 207.150 116.285 207.195 ;
        RECT 116.440 207.150 116.760 207.210 ;
        RECT 114.690 207.010 116.760 207.150 ;
        RECT 115.995 206.965 116.285 207.010 ;
        RECT 116.440 206.950 116.760 207.010 ;
        RECT 116.915 207.150 117.205 207.195 ;
        RECT 119.215 207.150 119.505 207.195 ;
        RECT 116.915 207.010 119.505 207.150 ;
        RECT 116.915 206.965 117.205 207.010 ;
        RECT 119.215 206.965 119.505 207.010 ;
        RECT 120.580 207.150 120.900 207.210 ;
        RECT 131.710 207.150 131.850 207.645 ;
        RECT 132.080 207.630 132.400 207.890 ;
        RECT 134.380 207.630 134.700 207.890 ;
        RECT 135.760 207.630 136.080 207.890 ;
        RECT 144.960 207.630 145.280 207.890 ;
        RECT 145.880 207.630 146.200 207.890 ;
        RECT 146.340 207.630 146.660 207.890 ;
        RECT 146.800 207.630 147.120 207.890 ;
        RECT 147.275 207.645 147.565 207.875 ;
        RECT 135.315 207.490 135.605 207.535 ;
        RECT 133.090 207.350 135.605 207.490 ;
        RECT 145.050 207.490 145.190 207.630 ;
        RECT 147.350 207.490 147.490 207.645 ;
        RECT 148.180 207.630 148.500 207.890 ;
        RECT 149.100 207.830 149.420 207.890 ;
        RECT 150.495 207.830 150.785 207.875 ;
        RECT 149.100 207.690 150.785 207.830 ;
        RECT 149.100 207.630 149.420 207.690 ;
        RECT 150.495 207.645 150.785 207.690 ;
        RECT 150.940 207.830 151.260 207.890 ;
        RECT 151.840 207.830 152.130 207.875 ;
        RECT 150.940 207.690 152.130 207.830 ;
        RECT 150.940 207.630 151.260 207.690 ;
        RECT 151.840 207.645 152.130 207.690 ;
        RECT 152.380 207.645 152.670 207.875 ;
        RECT 145.050 207.350 147.490 207.490 ;
        RECT 133.090 207.195 133.230 207.350 ;
        RECT 135.315 207.305 135.605 207.350 ;
        RECT 120.580 207.010 131.850 207.150 ;
        RECT 120.580 206.950 120.900 207.010 ;
        RECT 133.015 206.965 133.305 207.195 ;
        RECT 133.460 207.150 133.780 207.210 ;
        RECT 152.410 207.150 152.550 207.645 ;
        RECT 152.870 207.490 153.010 208.030 ;
        RECT 154.160 208.030 155.400 208.170 ;
        RECT 154.160 207.970 154.480 208.030 ;
        RECT 155.080 207.970 155.400 208.030 ;
        RECT 153.240 207.830 153.560 207.890 ;
        RECT 153.240 207.690 155.310 207.830 ;
        RECT 153.240 207.630 153.560 207.690 ;
        RECT 155.170 207.535 155.310 207.690 ;
        RECT 154.015 207.490 154.305 207.535 ;
        RECT 152.870 207.350 154.305 207.490 ;
        RECT 154.015 207.305 154.305 207.350 ;
        RECT 155.095 207.305 155.385 207.535 ;
        RECT 133.460 207.010 152.550 207.150 ;
        RECT 133.460 206.950 133.780 207.010 ;
        RECT 153.240 206.950 153.560 207.210 ;
        RECT 2.750 206.330 159.030 206.810 ;
        RECT 5.580 206.130 5.900 206.190 ;
        RECT 6.055 206.130 6.345 206.175 ;
        RECT 5.580 205.990 6.345 206.130 ;
        RECT 5.580 205.930 5.900 205.990 ;
        RECT 6.055 205.945 6.345 205.990 ;
        RECT 7.435 205.945 7.725 206.175 ;
        RECT 10.180 206.130 10.500 206.190 ;
        RECT 7.970 205.990 10.500 206.130 ;
        RECT 7.510 205.790 7.650 205.945 ;
        RECT 4.750 205.650 7.650 205.790 ;
        RECT 4.750 205.495 4.890 205.650 ;
        RECT 4.675 205.265 4.965 205.495 ;
        RECT 6.975 205.450 7.265 205.495 ;
        RECT 7.970 205.450 8.110 205.990 ;
        RECT 10.180 205.930 10.500 205.990 ;
        RECT 10.640 205.930 10.960 206.190 ;
        RECT 13.860 206.130 14.180 206.190 ;
        RECT 15.715 206.130 16.005 206.175 ;
        RECT 13.860 205.990 16.005 206.130 ;
        RECT 13.860 205.930 14.180 205.990 ;
        RECT 15.715 205.945 16.005 205.990 ;
        RECT 16.160 205.930 16.480 206.190 ;
        RECT 19.855 206.130 20.145 206.175 ;
        RECT 20.300 206.130 20.620 206.190 ;
        RECT 19.855 205.990 20.620 206.130 ;
        RECT 19.855 205.945 20.145 205.990 ;
        RECT 20.300 205.930 20.620 205.990 ;
        RECT 21.695 206.130 21.985 206.175 ;
        RECT 23.520 206.130 23.840 206.190 ;
        RECT 21.695 205.990 23.840 206.130 ;
        RECT 21.695 205.945 21.985 205.990 ;
        RECT 23.520 205.930 23.840 205.990 ;
        RECT 23.980 205.930 24.300 206.190 ;
        RECT 26.280 205.930 26.600 206.190 ;
        RECT 31.340 206.130 31.660 206.190 ;
        RECT 41.920 206.130 42.240 206.190 ;
        RECT 31.340 205.990 42.240 206.130 ;
        RECT 31.340 205.930 31.660 205.990 ;
        RECT 41.920 205.930 42.240 205.990 ;
        RECT 42.395 206.130 42.685 206.175 ;
        RECT 43.300 206.130 43.620 206.190 ;
        RECT 48.820 206.130 49.140 206.190 ;
        RECT 42.395 205.990 43.620 206.130 ;
        RECT 42.395 205.945 42.685 205.990 ;
        RECT 43.300 205.930 43.620 205.990 ;
        RECT 45.230 205.990 49.140 206.130 ;
        RECT 9.275 205.790 9.565 205.835 ;
        RECT 10.730 205.790 10.870 205.930 ;
        RECT 9.275 205.650 10.870 205.790 ;
        RECT 12.940 205.790 13.260 205.850 ;
        RECT 16.250 205.790 16.390 205.930 ;
        RECT 12.940 205.650 16.390 205.790 ;
        RECT 18.015 205.790 18.305 205.835 ;
        RECT 18.460 205.790 18.780 205.850 ;
        RECT 25.835 205.790 26.125 205.835 ;
        RECT 18.015 205.650 26.125 205.790 ;
        RECT 26.370 205.790 26.510 205.930 ;
        RECT 30.895 205.790 31.185 205.835 ;
        RECT 26.370 205.650 31.185 205.790 ;
        RECT 9.275 205.605 9.565 205.650 ;
        RECT 12.940 205.590 13.260 205.650 ;
        RECT 18.015 205.605 18.305 205.650 ;
        RECT 18.460 205.590 18.780 205.650 ;
        RECT 25.835 205.605 26.125 205.650 ;
        RECT 30.895 205.605 31.185 205.650 ;
        RECT 34.675 205.790 34.965 205.835 ;
        RECT 37.915 205.790 38.565 205.835 ;
        RECT 34.675 205.650 38.565 205.790 ;
        RECT 34.675 205.605 35.265 205.650 ;
        RECT 37.915 205.605 38.565 205.650 ;
        RECT 39.160 205.790 39.480 205.850 ;
        RECT 44.695 205.790 44.985 205.835 ;
        RECT 39.160 205.650 44.985 205.790 ;
        RECT 6.975 205.310 8.110 205.450 ;
        RECT 13.415 205.450 13.705 205.495 ;
        RECT 17.080 205.450 17.400 205.510 ;
        RECT 13.415 205.310 17.400 205.450 ;
        RECT 6.975 205.265 7.265 205.310 ;
        RECT 13.415 205.265 13.705 205.310 ;
        RECT 17.080 205.250 17.400 205.310 ;
        RECT 17.540 205.250 17.860 205.510 ;
        RECT 22.155 205.450 22.445 205.495 ;
        RECT 25.360 205.450 25.680 205.510 ;
        RECT 29.055 205.450 29.345 205.495 ;
        RECT 18.090 205.310 21.450 205.450 ;
        RECT 9.735 204.925 10.025 205.155 ;
        RECT 10.655 204.925 10.945 205.155 ;
        RECT 5.595 204.430 5.885 204.475 ;
        RECT 6.040 204.430 6.360 204.490 ;
        RECT 5.595 204.290 6.360 204.430 ;
        RECT 9.810 204.430 9.950 204.925 ;
        RECT 10.730 204.770 10.870 204.925 ;
        RECT 12.480 204.910 12.800 205.170 ;
        RECT 12.940 204.910 13.260 205.170 ;
        RECT 14.320 204.770 14.640 204.830 ;
        RECT 18.090 204.770 18.230 205.310 ;
        RECT 18.935 205.110 19.225 205.155 ;
        RECT 20.300 205.110 20.620 205.170 ;
        RECT 18.935 204.970 20.620 205.110 ;
        RECT 18.935 204.925 19.225 204.970 ;
        RECT 20.300 204.910 20.620 204.970 ;
        RECT 10.730 204.630 14.640 204.770 ;
        RECT 14.320 204.570 14.640 204.630 ;
        RECT 14.870 204.630 18.230 204.770 ;
        RECT 14.870 204.430 15.010 204.630 ;
        RECT 9.810 204.290 15.010 204.430 ;
        RECT 5.595 204.245 5.885 204.290 ;
        RECT 6.040 204.230 6.360 204.290 ;
        RECT 15.240 204.230 15.560 204.490 ;
        RECT 20.390 204.430 20.530 204.910 ;
        RECT 21.310 204.830 21.450 205.310 ;
        RECT 22.155 205.310 25.680 205.450 ;
        RECT 22.155 205.265 22.445 205.310 ;
        RECT 25.360 205.250 25.680 205.310 ;
        RECT 28.670 205.310 29.345 205.450 ;
        RECT 28.670 205.170 28.810 205.310 ;
        RECT 29.055 205.265 29.345 205.310 ;
        RECT 29.975 205.265 30.265 205.495 ;
        RECT 34.975 205.290 35.265 205.605 ;
        RECT 39.160 205.590 39.480 205.650 ;
        RECT 44.695 205.605 44.985 205.650 ;
        RECT 36.055 205.450 36.345 205.495 ;
        RECT 39.635 205.450 39.925 205.495 ;
        RECT 41.470 205.450 41.760 205.495 ;
        RECT 36.055 205.310 41.760 205.450 ;
        RECT 22.615 204.925 22.905 205.155 ;
        RECT 23.520 205.110 23.840 205.170 ;
        RECT 26.295 205.110 26.585 205.155 ;
        RECT 23.520 204.970 26.585 205.110 ;
        RECT 21.220 204.570 21.540 204.830 ;
        RECT 22.690 204.430 22.830 204.925 ;
        RECT 23.520 204.910 23.840 204.970 ;
        RECT 26.295 204.925 26.585 204.970 ;
        RECT 27.200 204.910 27.520 205.170 ;
        RECT 28.580 204.910 28.900 205.170 ;
        RECT 23.980 204.770 24.300 204.830 ;
        RECT 29.055 204.770 29.345 204.815 ;
        RECT 23.980 204.630 29.345 204.770 ;
        RECT 23.980 204.570 24.300 204.630 ;
        RECT 29.055 204.585 29.345 204.630 ;
        RECT 20.390 204.290 22.830 204.430 ;
        RECT 24.900 204.430 25.220 204.490 ;
        RECT 30.050 204.430 30.190 205.265 ;
        RECT 34.560 205.110 34.880 205.170 ;
        RECT 35.110 205.110 35.250 205.290 ;
        RECT 36.055 205.265 36.345 205.310 ;
        RECT 39.635 205.265 39.925 205.310 ;
        RECT 41.470 205.265 41.760 205.310 ;
        RECT 41.920 205.250 42.240 205.510 ;
        RECT 43.300 205.450 43.620 205.510 ;
        RECT 44.235 205.450 44.525 205.495 ;
        RECT 45.230 205.450 45.370 205.990 ;
        RECT 48.820 205.930 49.140 205.990 ;
        RECT 49.280 206.130 49.600 206.190 ;
        RECT 50.215 206.130 50.505 206.175 ;
        RECT 49.280 205.990 50.505 206.130 ;
        RECT 49.280 205.930 49.600 205.990 ;
        RECT 50.215 205.945 50.505 205.990 ;
        RECT 56.180 206.130 56.500 206.190 ;
        RECT 62.620 206.130 62.940 206.190 ;
        RECT 85.620 206.130 85.940 206.190 ;
        RECT 56.180 205.990 57.790 206.130 ;
        RECT 56.180 205.930 56.500 205.990 ;
        RECT 47.915 205.790 48.205 205.835 ;
        RECT 50.660 205.790 50.980 205.850 ;
        RECT 57.650 205.835 57.790 205.990 ;
        RECT 62.620 205.990 85.940 206.130 ;
        RECT 62.620 205.930 62.940 205.990 ;
        RECT 85.620 205.930 85.940 205.990 ;
        RECT 86.080 206.130 86.400 206.190 ;
        RECT 87.935 206.130 88.225 206.175 ;
        RECT 86.080 205.990 88.225 206.130 ;
        RECT 86.080 205.930 86.400 205.990 ;
        RECT 87.935 205.945 88.225 205.990 ;
        RECT 88.380 205.930 88.700 206.190 ;
        RECT 88.840 205.930 89.160 206.190 ;
        RECT 91.600 206.130 91.920 206.190 ;
        RECT 89.390 205.990 91.920 206.130 ;
        RECT 47.915 205.650 50.980 205.790 ;
        RECT 47.915 205.605 48.205 205.650 ;
        RECT 50.660 205.590 50.980 205.650 ;
        RECT 57.575 205.605 57.865 205.835 ;
        RECT 64.920 205.790 65.240 205.850 ;
        RECT 83.320 205.790 83.640 205.850 ;
        RECT 88.470 205.790 88.610 205.930 ;
        RECT 64.920 205.650 83.640 205.790 ;
        RECT 64.920 205.590 65.240 205.650 ;
        RECT 83.320 205.590 83.640 205.650 ;
        RECT 85.710 205.650 88.610 205.790 ;
        RECT 43.300 205.310 45.370 205.450 ;
        RECT 48.375 205.450 48.665 205.495 ;
        RECT 51.580 205.450 51.900 205.510 ;
        RECT 48.375 205.310 51.900 205.450 ;
        RECT 43.300 205.250 43.620 205.310 ;
        RECT 44.235 205.265 44.525 205.310 ;
        RECT 48.375 205.265 48.665 205.310 ;
        RECT 51.580 205.250 51.900 205.310 ;
        RECT 55.260 205.450 55.580 205.510 ;
        RECT 56.195 205.450 56.485 205.495 ;
        RECT 55.260 205.310 56.485 205.450 ;
        RECT 55.260 205.250 55.580 205.310 ;
        RECT 56.195 205.265 56.485 205.310 ;
        RECT 34.560 204.970 35.250 205.110 ;
        RECT 40.555 205.110 40.845 205.155 ;
        RECT 40.555 204.970 43.450 205.110 ;
        RECT 34.560 204.910 34.880 204.970 ;
        RECT 40.555 204.925 40.845 204.970 ;
        RECT 36.055 204.770 36.345 204.815 ;
        RECT 39.175 204.770 39.465 204.815 ;
        RECT 41.065 204.770 41.355 204.815 ;
        RECT 36.055 204.630 41.355 204.770 ;
        RECT 43.310 204.770 43.450 204.970 ;
        RECT 45.140 204.910 45.460 205.170 ;
        RECT 47.455 205.110 47.745 205.155 ;
        RECT 49.740 205.110 50.060 205.170 ;
        RECT 47.455 204.970 50.060 205.110 ;
        RECT 47.455 204.925 47.745 204.970 ;
        RECT 49.740 204.910 50.060 204.970 ;
        RECT 53.420 204.910 53.740 205.170 ;
        RECT 54.800 204.770 55.120 204.830 ;
        RECT 43.310 204.630 55.120 204.770 ;
        RECT 36.055 204.585 36.345 204.630 ;
        RECT 39.175 204.585 39.465 204.630 ;
        RECT 41.065 204.585 41.355 204.630 ;
        RECT 54.800 204.570 55.120 204.630 ;
        RECT 55.260 204.570 55.580 204.830 ;
        RECT 56.270 204.770 56.410 205.265 ;
        RECT 58.020 205.250 58.340 205.510 ;
        RECT 58.955 205.450 59.245 205.495 ;
        RECT 59.400 205.450 59.720 205.510 ;
        RECT 66.760 205.450 67.080 205.510 ;
        RECT 58.955 205.310 67.080 205.450 ;
        RECT 58.955 205.265 59.245 205.310 ;
        RECT 59.400 205.250 59.720 205.310 ;
        RECT 66.760 205.250 67.080 205.310 ;
        RECT 68.140 205.250 68.460 205.510 ;
        RECT 68.600 205.250 68.920 205.510 ;
        RECT 69.520 205.250 69.840 205.510 ;
        RECT 84.700 205.250 85.020 205.510 ;
        RECT 85.710 205.495 85.850 205.650 ;
        RECT 85.635 205.265 85.925 205.495 ;
        RECT 86.080 205.250 86.400 205.510 ;
        RECT 86.555 205.450 86.845 205.495 ;
        RECT 89.390 205.450 89.530 205.990 ;
        RECT 91.600 205.930 91.920 205.990 ;
        RECT 92.060 206.130 92.380 206.190 ;
        RECT 97.580 206.130 97.900 206.190 ;
        RECT 104.480 206.130 104.800 206.190 ;
        RECT 92.060 205.990 97.900 206.130 ;
        RECT 92.060 205.930 92.380 205.990 ;
        RECT 97.580 205.930 97.900 205.990 ;
        RECT 101.810 205.990 104.800 206.130 ;
        RECT 90.680 205.790 91.000 205.850 ;
        RECT 90.680 205.650 100.110 205.790 ;
        RECT 90.680 205.590 91.000 205.650 ;
        RECT 99.970 205.510 100.110 205.650 ;
        RECT 86.555 205.310 89.530 205.450 ;
        RECT 86.555 205.265 86.845 205.310 ;
        RECT 89.760 205.250 90.080 205.510 ;
        RECT 95.280 205.250 95.600 205.510 ;
        RECT 95.740 205.250 96.060 205.510 ;
        RECT 96.215 205.265 96.505 205.495 ;
        RECT 57.115 205.110 57.405 205.155 ;
        RECT 58.495 205.110 58.785 205.155 ;
        RECT 57.115 204.970 58.785 205.110 ;
        RECT 68.230 205.110 68.370 205.250 ;
        RECT 77.800 205.110 78.120 205.170 ;
        RECT 68.230 204.970 78.120 205.110 ;
        RECT 57.115 204.925 57.405 204.970 ;
        RECT 58.495 204.925 58.785 204.970 ;
        RECT 77.800 204.910 78.120 204.970 ;
        RECT 82.860 205.110 83.180 205.170 ;
        RECT 82.860 204.970 89.070 205.110 ;
        RECT 82.860 204.910 83.180 204.970 ;
        RECT 72.740 204.770 73.060 204.830 ;
        RECT 75.960 204.770 76.280 204.830 ;
        RECT 56.270 204.630 68.830 204.770 ;
        RECT 24.900 204.290 30.190 204.430 ;
        RECT 24.900 204.230 25.220 204.290 ;
        RECT 32.260 204.230 32.580 204.490 ;
        RECT 33.195 204.430 33.485 204.475 ;
        RECT 36.860 204.430 37.180 204.490 ;
        RECT 43.300 204.430 43.620 204.490 ;
        RECT 33.195 204.290 43.620 204.430 ;
        RECT 33.195 204.245 33.485 204.290 ;
        RECT 36.860 204.230 37.180 204.290 ;
        RECT 43.300 204.230 43.620 204.290 ;
        RECT 45.600 204.430 45.920 204.490 ;
        RECT 50.675 204.430 50.965 204.475 ;
        RECT 45.600 204.290 50.965 204.430 ;
        RECT 45.600 204.230 45.920 204.290 ;
        RECT 50.675 204.245 50.965 204.290 ;
        RECT 57.575 204.430 57.865 204.475 ;
        RECT 58.940 204.430 59.260 204.490 ;
        RECT 57.575 204.290 59.260 204.430 ;
        RECT 57.575 204.245 57.865 204.290 ;
        RECT 58.940 204.230 59.260 204.290 ;
        RECT 63.080 204.430 63.400 204.490 ;
        RECT 65.380 204.430 65.700 204.490 ;
        RECT 63.080 204.290 65.700 204.430 ;
        RECT 68.690 204.430 68.830 204.630 ;
        RECT 72.740 204.630 76.280 204.770 ;
        RECT 72.740 204.570 73.060 204.630 ;
        RECT 75.960 204.570 76.280 204.630 ;
        RECT 84.240 204.770 84.560 204.830 ;
        RECT 88.380 204.770 88.700 204.830 ;
        RECT 84.240 204.630 88.700 204.770 ;
        RECT 88.930 204.770 89.070 204.970 ;
        RECT 90.235 204.925 90.525 205.155 ;
        RECT 90.695 204.925 90.985 205.155 ;
        RECT 91.155 205.110 91.445 205.155 ;
        RECT 92.060 205.110 92.380 205.170 ;
        RECT 91.155 204.970 92.380 205.110 ;
        RECT 91.155 204.925 91.445 204.970 ;
        RECT 90.310 204.770 90.450 204.925 ;
        RECT 88.930 204.630 90.450 204.770 ;
        RECT 90.770 204.770 90.910 204.925 ;
        RECT 92.060 204.910 92.380 204.970 ;
        RECT 95.830 204.770 95.970 205.250 ;
        RECT 96.290 205.110 96.430 205.265 ;
        RECT 96.660 205.250 96.980 205.510 ;
        RECT 97.120 205.250 97.440 205.510 ;
        RECT 98.960 205.250 99.280 205.510 ;
        RECT 99.880 205.250 100.200 205.510 ;
        RECT 100.355 205.450 100.645 205.495 ;
        RECT 101.810 205.450 101.950 205.990 ;
        RECT 104.480 205.930 104.800 205.990 ;
        RECT 104.940 206.130 105.260 206.190 ;
        RECT 108.160 206.130 108.480 206.190 ;
        RECT 111.840 206.130 112.160 206.190 ;
        RECT 104.940 205.990 112.160 206.130 ;
        RECT 104.940 205.930 105.260 205.990 ;
        RECT 108.160 205.930 108.480 205.990 ;
        RECT 111.840 205.930 112.160 205.990 ;
        RECT 112.315 206.130 112.605 206.175 ;
        RECT 112.760 206.130 113.080 206.190 ;
        RECT 112.315 205.990 113.080 206.130 ;
        RECT 112.315 205.945 112.605 205.990 ;
        RECT 112.760 205.930 113.080 205.990 ;
        RECT 114.600 205.930 114.920 206.190 ;
        RECT 115.060 206.130 115.380 206.190 ;
        RECT 123.340 206.130 123.660 206.190 ;
        RECT 123.815 206.130 124.105 206.175 ;
        RECT 115.060 205.990 119.430 206.130 ;
        RECT 115.060 205.930 115.380 205.990 ;
        RECT 108.635 205.790 108.925 205.835 ;
        RECT 118.740 205.790 119.060 205.850 ;
        RECT 102.330 205.650 108.925 205.790 ;
        RECT 102.330 205.495 102.470 205.650 ;
        RECT 108.635 205.605 108.925 205.650 ;
        RECT 109.170 205.650 119.060 205.790 ;
        RECT 119.290 205.790 119.430 205.990 ;
        RECT 123.340 205.990 124.105 206.130 ;
        RECT 123.340 205.930 123.660 205.990 ;
        RECT 123.815 205.945 124.105 205.990 ;
        RECT 134.380 205.930 134.700 206.190 ;
        RECT 146.340 206.130 146.660 206.190 ;
        RECT 146.815 206.130 147.105 206.175 ;
        RECT 146.340 205.990 147.105 206.130 ;
        RECT 146.340 205.930 146.660 205.990 ;
        RECT 146.815 205.945 147.105 205.990 ;
        RECT 153.240 205.930 153.560 206.190 ;
        RECT 134.470 205.790 134.610 205.930 ;
        RECT 153.330 205.790 153.470 205.930 ;
        RECT 119.290 205.650 133.230 205.790 ;
        RECT 134.470 205.650 135.070 205.790 ;
        RECT 100.355 205.310 101.950 205.450 ;
        RECT 100.355 205.265 100.645 205.310 ;
        RECT 102.195 205.265 102.485 205.495 ;
        RECT 102.640 205.250 102.960 205.510 ;
        RECT 105.860 205.250 106.180 205.510 ;
        RECT 107.240 205.450 107.560 205.510 ;
        RECT 109.170 205.495 109.310 205.650 ;
        RECT 118.740 205.590 119.060 205.650 ;
        RECT 133.090 205.510 133.230 205.650 ;
        RECT 108.175 205.450 108.465 205.495 ;
        RECT 107.240 205.310 108.465 205.450 ;
        RECT 107.240 205.250 107.560 205.310 ;
        RECT 108.175 205.265 108.465 205.310 ;
        RECT 109.095 205.265 109.385 205.495 ;
        RECT 110.475 205.450 110.765 205.495 ;
        RECT 113.695 205.450 113.985 205.495 ;
        RECT 110.475 205.310 113.985 205.450 ;
        RECT 110.475 205.265 110.765 205.310 ;
        RECT 113.695 205.265 113.985 205.310 ;
        RECT 115.980 205.450 116.300 205.510 ;
        RECT 133.000 205.450 133.320 205.510 ;
        RECT 134.930 205.495 135.070 205.650 ;
        RECT 145.050 205.650 153.470 205.790 ;
        RECT 133.475 205.450 133.765 205.495 ;
        RECT 115.980 205.310 125.870 205.450 ;
        RECT 99.050 205.110 99.190 205.250 ;
        RECT 100.815 205.110 101.105 205.155 ;
        RECT 96.290 204.970 97.350 205.110 ;
        RECT 99.050 204.970 101.105 205.110 ;
        RECT 90.770 204.630 95.970 204.770 ;
        RECT 84.240 204.570 84.560 204.630 ;
        RECT 88.380 204.570 88.700 204.630 ;
        RECT 70.900 204.430 71.220 204.490 ;
        RECT 68.690 204.290 71.220 204.430 ;
        RECT 63.080 204.230 63.400 204.290 ;
        RECT 65.380 204.230 65.700 204.290 ;
        RECT 70.900 204.230 71.220 204.290 ;
        RECT 71.820 204.430 72.140 204.490 ;
        RECT 74.120 204.430 74.440 204.490 ;
        RECT 71.820 204.290 74.440 204.430 ;
        RECT 71.820 204.230 72.140 204.290 ;
        RECT 74.120 204.230 74.440 204.290 ;
        RECT 75.040 204.430 75.360 204.490 ;
        RECT 88.840 204.430 89.160 204.490 ;
        RECT 75.040 204.290 89.160 204.430 ;
        RECT 90.310 204.430 90.450 204.630 ;
        RECT 96.660 204.430 96.980 204.490 ;
        RECT 90.310 204.290 96.980 204.430 ;
        RECT 97.210 204.430 97.350 204.970 ;
        RECT 100.815 204.925 101.105 204.970 ;
        RECT 101.275 205.110 101.565 205.155 ;
        RECT 101.275 204.970 102.470 205.110 ;
        RECT 101.275 204.925 101.565 204.970 ;
        RECT 98.515 204.770 98.805 204.815 ;
        RECT 102.330 204.770 102.470 204.970 ;
        RECT 103.100 204.910 103.420 205.170 ;
        RECT 105.950 205.110 106.090 205.250 ;
        RECT 104.570 204.970 106.090 205.110 ;
        RECT 107.700 205.110 108.020 205.170 ;
        RECT 110.015 205.110 110.305 205.155 ;
        RECT 107.700 204.970 110.305 205.110 ;
        RECT 104.570 204.815 104.710 204.970 ;
        RECT 107.700 204.910 108.020 204.970 ;
        RECT 110.015 204.925 110.305 204.970 ;
        RECT 98.515 204.630 101.950 204.770 ;
        RECT 102.330 204.630 103.330 204.770 ;
        RECT 98.515 204.585 98.805 204.630 ;
        RECT 98.975 204.430 99.265 204.475 ;
        RECT 97.210 204.290 99.265 204.430 ;
        RECT 75.040 204.230 75.360 204.290 ;
        RECT 88.840 204.230 89.160 204.290 ;
        RECT 96.660 204.230 96.980 204.290 ;
        RECT 98.975 204.245 99.265 204.290 ;
        RECT 99.880 204.430 100.200 204.490 ;
        RECT 101.260 204.430 101.580 204.490 ;
        RECT 99.880 204.290 101.580 204.430 ;
        RECT 101.810 204.430 101.950 204.630 ;
        RECT 102.655 204.430 102.945 204.475 ;
        RECT 101.810 204.290 102.945 204.430 ;
        RECT 103.190 204.430 103.330 204.630 ;
        RECT 104.495 204.585 104.785 204.815 ;
        RECT 105.860 204.770 106.180 204.830 ;
        RECT 110.550 204.770 110.690 205.265 ;
        RECT 115.980 205.250 116.300 205.310 ;
        RECT 125.730 205.170 125.870 205.310 ;
        RECT 133.000 205.310 133.765 205.450 ;
        RECT 133.000 205.250 133.320 205.310 ;
        RECT 133.475 205.265 133.765 205.310 ;
        RECT 134.395 205.265 134.685 205.495 ;
        RECT 134.855 205.265 135.145 205.495 ;
        RECT 135.315 205.450 135.605 205.495 ;
        RECT 135.315 205.310 144.270 205.450 ;
        RECT 135.315 205.265 135.605 205.310 ;
        RECT 110.935 204.925 111.225 205.155 ;
        RECT 111.395 204.925 111.685 205.155 ;
        RECT 112.775 205.110 113.065 205.155 ;
        RECT 114.600 205.110 114.920 205.170 ;
        RECT 112.775 204.970 114.920 205.110 ;
        RECT 112.775 204.925 113.065 204.970 ;
        RECT 105.860 204.630 110.690 204.770 ;
        RECT 105.860 204.570 106.180 204.630 ;
        RECT 104.940 204.430 105.260 204.490 ;
        RECT 103.190 204.290 105.260 204.430 ;
        RECT 99.880 204.230 100.200 204.290 ;
        RECT 101.260 204.230 101.580 204.290 ;
        RECT 102.655 204.245 102.945 204.290 ;
        RECT 104.940 204.230 105.260 204.290 ;
        RECT 106.320 204.430 106.640 204.490 ;
        RECT 110.460 204.430 110.780 204.490 ;
        RECT 111.010 204.430 111.150 204.925 ;
        RECT 111.470 204.770 111.610 204.925 ;
        RECT 114.600 204.910 114.920 204.970 ;
        RECT 120.580 204.910 120.900 205.170 ;
        RECT 124.720 204.910 125.040 205.170 ;
        RECT 125.180 204.910 125.500 205.170 ;
        RECT 125.640 204.910 125.960 205.170 ;
        RECT 126.115 204.925 126.405 205.155 ;
        RECT 130.700 205.110 131.020 205.170 ;
        RECT 134.470 205.110 134.610 205.265 ;
        RECT 130.700 204.970 134.610 205.110 ;
        RECT 113.220 204.770 113.540 204.830 ;
        RECT 120.670 204.770 120.810 204.910 ;
        RECT 111.470 204.630 120.810 204.770 ;
        RECT 126.190 204.770 126.330 204.925 ;
        RECT 130.700 204.910 131.020 204.970 ;
        RECT 136.235 204.925 136.525 205.155 ;
        RECT 144.130 205.110 144.270 205.310 ;
        RECT 144.500 205.250 144.820 205.510 ;
        RECT 145.050 205.495 145.190 205.650 ;
        RECT 144.975 205.265 145.265 205.495 ;
        RECT 145.420 205.450 145.740 205.510 ;
        RECT 145.895 205.450 146.185 205.495 ;
        RECT 145.420 205.310 146.185 205.450 ;
        RECT 145.420 205.250 145.740 205.310 ;
        RECT 145.895 205.265 146.185 205.310 ;
        RECT 149.560 205.110 149.880 205.170 ;
        RECT 144.130 204.970 149.880 205.110 ;
        RECT 135.775 204.770 136.065 204.815 ;
        RECT 126.190 204.630 136.065 204.770 ;
        RECT 113.220 204.570 113.540 204.630 ;
        RECT 135.775 204.585 136.065 204.630 ;
        RECT 106.320 204.290 111.150 204.430 ;
        RECT 117.360 204.430 117.680 204.490 ;
        RECT 120.120 204.430 120.440 204.490 ;
        RECT 117.360 204.290 120.440 204.430 ;
        RECT 106.320 204.230 106.640 204.290 ;
        RECT 110.460 204.230 110.780 204.290 ;
        RECT 117.360 204.230 117.680 204.290 ;
        RECT 120.120 204.230 120.440 204.290 ;
        RECT 124.260 204.430 124.580 204.490 ;
        RECT 134.840 204.430 135.160 204.490 ;
        RECT 136.310 204.430 136.450 204.925 ;
        RECT 149.560 204.910 149.880 204.970 ;
        RECT 145.435 204.585 145.725 204.815 ;
        RECT 140.820 204.430 141.140 204.490 ;
        RECT 124.260 204.290 141.140 204.430 ;
        RECT 124.260 204.230 124.580 204.290 ;
        RECT 134.840 204.230 135.160 204.290 ;
        RECT 140.820 204.230 141.140 204.290 ;
        RECT 144.500 204.430 144.820 204.490 ;
        RECT 145.510 204.430 145.650 204.585 ;
        RECT 144.500 204.290 145.650 204.430 ;
        RECT 144.500 204.230 144.820 204.290 ;
        RECT 2.750 203.610 158.230 204.090 ;
        RECT 12.940 203.410 13.260 203.470 ;
        RECT 13.860 203.410 14.180 203.470 ;
        RECT 12.940 203.270 14.180 203.410 ;
        RECT 12.940 203.210 13.260 203.270 ;
        RECT 13.860 203.210 14.180 203.270 ;
        RECT 15.240 203.210 15.560 203.470 ;
        RECT 17.540 203.410 17.860 203.470 ;
        RECT 18.935 203.410 19.225 203.455 ;
        RECT 24.440 203.410 24.760 203.470 ;
        RECT 17.540 203.270 19.225 203.410 ;
        RECT 17.540 203.210 17.860 203.270 ;
        RECT 18.935 203.225 19.225 203.270 ;
        RECT 19.470 203.270 24.760 203.410 ;
        RECT 6.005 203.070 6.295 203.115 ;
        RECT 7.895 203.070 8.185 203.115 ;
        RECT 11.015 203.070 11.305 203.115 ;
        RECT 14.335 203.070 14.625 203.115 ;
        RECT 6.005 202.930 11.305 203.070 ;
        RECT 6.005 202.885 6.295 202.930 ;
        RECT 7.895 202.885 8.185 202.930 ;
        RECT 11.015 202.885 11.305 202.930 ;
        RECT 13.720 202.930 14.625 203.070 ;
        RECT 5.120 202.530 5.440 202.790 ;
        RECT 6.515 202.730 6.805 202.775 ;
        RECT 13.720 202.730 13.860 202.930 ;
        RECT 14.335 202.885 14.625 202.930 ;
        RECT 6.515 202.590 13.860 202.730 ;
        RECT 6.515 202.545 6.805 202.590 ;
        RECT 15.330 202.435 15.470 203.210 ;
        RECT 16.160 203.070 16.480 203.130 ;
        RECT 19.470 203.070 19.610 203.270 ;
        RECT 24.440 203.210 24.760 203.270 ;
        RECT 24.900 203.210 25.220 203.470 ;
        RECT 27.200 203.410 27.520 203.470 ;
        RECT 25.450 203.270 27.520 203.410 ;
        RECT 16.160 202.930 19.610 203.070 ;
        RECT 16.160 202.870 16.480 202.930 ;
        RECT 17.170 202.435 17.310 202.930 ;
        RECT 20.760 202.870 21.080 203.130 ;
        RECT 24.990 203.070 25.130 203.210 ;
        RECT 21.310 202.930 25.130 203.070 ;
        RECT 17.555 202.545 17.845 202.775 ;
        RECT 18.000 202.730 18.320 202.790 ;
        RECT 18.000 202.590 19.610 202.730 ;
        RECT 5.600 202.390 5.890 202.435 ;
        RECT 7.435 202.390 7.725 202.435 ;
        RECT 11.015 202.390 11.305 202.435 ;
        RECT 5.600 202.250 11.305 202.390 ;
        RECT 5.600 202.205 5.890 202.250 ;
        RECT 7.435 202.205 7.725 202.250 ;
        RECT 11.015 202.205 11.305 202.250 ;
        RECT 12.095 202.095 12.385 202.410 ;
        RECT 15.255 202.205 15.545 202.435 ;
        RECT 17.095 202.205 17.385 202.435 ;
        RECT 17.630 202.390 17.770 202.545 ;
        RECT 18.000 202.530 18.320 202.590 ;
        RECT 19.470 202.435 19.610 202.590 ;
        RECT 21.310 202.435 21.450 202.930 ;
        RECT 24.900 202.730 25.220 202.790 ;
        RECT 25.450 202.775 25.590 203.270 ;
        RECT 27.200 203.210 27.520 203.270 ;
        RECT 28.120 203.210 28.440 203.470 ;
        RECT 28.580 203.210 28.900 203.470 ;
        RECT 41.015 203.410 41.305 203.455 ;
        RECT 52.500 203.410 52.820 203.470 ;
        RECT 41.015 203.270 52.820 203.410 ;
        RECT 41.015 203.225 41.305 203.270 ;
        RECT 52.500 203.210 52.820 203.270 ;
        RECT 54.800 203.210 55.120 203.470 ;
        RECT 55.260 203.210 55.580 203.470 ;
        RECT 56.195 203.410 56.485 203.455 ;
        RECT 58.020 203.410 58.340 203.470 ;
        RECT 79.180 203.410 79.500 203.470 ;
        RECT 56.195 203.270 58.340 203.410 ;
        RECT 56.195 203.225 56.485 203.270 ;
        RECT 58.020 203.210 58.340 203.270 ;
        RECT 61.330 203.270 79.500 203.410 ;
        RECT 31.765 203.070 32.055 203.115 ;
        RECT 33.655 203.070 33.945 203.115 ;
        RECT 36.775 203.070 37.065 203.115 ;
        RECT 25.910 202.930 30.190 203.070 ;
        RECT 21.770 202.590 25.220 202.730 ;
        RECT 19.395 202.390 19.685 202.435 ;
        RECT 21.235 202.390 21.525 202.435 ;
        RECT 17.630 202.250 18.230 202.390 ;
        RECT 8.795 202.050 9.445 202.095 ;
        RECT 12.095 202.050 12.685 202.095 ;
        RECT 13.400 202.050 13.720 202.110 ;
        RECT 8.795 201.910 13.720 202.050 ;
        RECT 8.795 201.865 9.445 201.910 ;
        RECT 12.395 201.865 12.685 201.910 ;
        RECT 13.400 201.850 13.720 201.910 ;
        RECT 16.620 202.050 16.940 202.110 ;
        RECT 18.090 202.050 18.230 202.250 ;
        RECT 19.395 202.250 21.525 202.390 ;
        RECT 19.395 202.205 19.685 202.250 ;
        RECT 21.235 202.205 21.525 202.250 ;
        RECT 16.620 201.910 18.230 202.050 ;
        RECT 16.620 201.850 16.940 201.910 ;
        RECT 18.090 201.710 18.230 201.910 ;
        RECT 18.920 202.050 19.240 202.110 ;
        RECT 19.855 202.050 20.145 202.095 ;
        RECT 18.920 201.910 20.145 202.050 ;
        RECT 18.920 201.850 19.240 201.910 ;
        RECT 19.855 201.865 20.145 201.910 ;
        RECT 20.300 202.050 20.620 202.110 ;
        RECT 20.775 202.050 21.065 202.095 ;
        RECT 21.770 202.050 21.910 202.590 ;
        RECT 24.900 202.530 25.220 202.590 ;
        RECT 25.375 202.545 25.665 202.775 ;
        RECT 25.910 202.390 26.050 202.930 ;
        RECT 30.050 202.730 30.190 202.930 ;
        RECT 31.765 202.930 37.065 203.070 ;
        RECT 31.765 202.885 32.055 202.930 ;
        RECT 33.655 202.885 33.945 202.930 ;
        RECT 36.775 202.885 37.065 202.930 ;
        RECT 41.460 203.070 41.780 203.130 ;
        RECT 43.725 203.070 44.015 203.115 ;
        RECT 45.615 203.070 45.905 203.115 ;
        RECT 48.735 203.070 49.025 203.115 ;
        RECT 41.460 202.930 43.530 203.070 ;
        RECT 41.460 202.870 41.780 202.930 ;
        RECT 41.920 202.730 42.240 202.790 ;
        RECT 42.855 202.730 43.145 202.775 ;
        RECT 30.050 202.590 41.230 202.730 ;
        RECT 22.690 202.250 26.050 202.390 ;
        RECT 26.740 202.390 27.060 202.450 ;
        RECT 30.050 202.435 30.190 202.590 ;
        RECT 29.515 202.390 29.805 202.435 ;
        RECT 26.740 202.250 29.805 202.390 ;
        RECT 20.300 201.910 21.910 202.050 ;
        RECT 20.300 201.850 20.620 201.910 ;
        RECT 20.775 201.865 21.065 201.910 ;
        RECT 22.140 201.850 22.460 202.110 ;
        RECT 22.690 201.710 22.830 202.250 ;
        RECT 26.740 202.190 27.060 202.250 ;
        RECT 29.515 202.205 29.805 202.250 ;
        RECT 29.975 202.205 30.265 202.435 ;
        RECT 30.420 202.190 30.740 202.450 ;
        RECT 30.880 202.190 31.200 202.450 ;
        RECT 41.090 202.435 41.230 202.590 ;
        RECT 41.920 202.590 43.145 202.730 ;
        RECT 43.390 202.730 43.530 202.930 ;
        RECT 43.725 202.930 49.025 203.070 ;
        RECT 43.725 202.885 44.015 202.930 ;
        RECT 45.615 202.885 45.905 202.930 ;
        RECT 48.735 202.885 49.025 202.930 ;
        RECT 51.580 202.870 51.900 203.130 ;
        RECT 55.350 203.070 55.490 203.210 ;
        RECT 57.100 203.070 57.420 203.130 ;
        RECT 55.350 202.930 57.420 203.070 ;
        RECT 57.100 202.870 57.420 202.930 ;
        RECT 58.940 202.870 59.260 203.130 ;
        RECT 61.330 202.775 61.470 203.270 ;
        RECT 79.180 203.210 79.500 203.270 ;
        RECT 85.160 203.210 85.480 203.470 ;
        RECT 86.080 203.410 86.400 203.470 ;
        RECT 87.015 203.410 87.305 203.455 ;
        RECT 86.080 203.270 87.305 203.410 ;
        RECT 86.080 203.210 86.400 203.270 ;
        RECT 87.015 203.225 87.305 203.270 ;
        RECT 87.460 203.410 87.780 203.470 ;
        RECT 87.460 203.270 97.350 203.410 ;
        RECT 87.460 203.210 87.780 203.270 ;
        RECT 63.080 203.070 63.400 203.130 ;
        RECT 64.920 203.070 65.240 203.130 ;
        RECT 74.135 203.070 74.425 203.115 ;
        RECT 62.710 202.930 63.400 203.070 ;
        RECT 62.710 202.775 62.850 202.930 ;
        RECT 63.080 202.870 63.400 202.930 ;
        RECT 63.630 202.930 65.240 203.070 ;
        RECT 60.795 202.730 61.085 202.775 ;
        RECT 43.390 202.590 55.950 202.730 ;
        RECT 41.920 202.530 42.240 202.590 ;
        RECT 42.855 202.545 43.145 202.590 ;
        RECT 31.360 202.390 31.650 202.435 ;
        RECT 33.195 202.390 33.485 202.435 ;
        RECT 36.775 202.390 37.065 202.435 ;
        RECT 31.360 202.250 37.065 202.390 ;
        RECT 31.360 202.205 31.650 202.250 ;
        RECT 33.195 202.205 33.485 202.250 ;
        RECT 36.775 202.205 37.065 202.250 ;
        RECT 28.545 202.050 28.835 202.095 ;
        RECT 30.510 202.050 30.650 202.190 ;
        RECT 32.275 202.050 32.565 202.095 ;
        RECT 28.545 201.910 30.190 202.050 ;
        RECT 30.510 201.910 32.565 202.050 ;
        RECT 28.545 201.865 28.835 201.910 ;
        RECT 30.050 201.770 30.190 201.910 ;
        RECT 32.275 201.865 32.565 201.910 ;
        RECT 34.555 202.050 35.205 202.095 ;
        RECT 37.320 202.050 37.640 202.110 ;
        RECT 37.855 202.095 38.145 202.410 ;
        RECT 40.095 202.205 40.385 202.435 ;
        RECT 41.015 202.205 41.305 202.435 ;
        RECT 43.320 202.390 43.610 202.435 ;
        RECT 45.155 202.390 45.445 202.435 ;
        RECT 48.735 202.390 49.025 202.435 ;
        RECT 43.320 202.250 49.025 202.390 ;
        RECT 43.320 202.205 43.610 202.250 ;
        RECT 45.155 202.205 45.445 202.250 ;
        RECT 48.735 202.205 49.025 202.250 ;
        RECT 49.740 202.410 50.060 202.450 ;
        RECT 37.855 202.050 38.445 202.095 ;
        RECT 34.555 201.910 38.445 202.050 ;
        RECT 34.555 201.865 35.205 201.910 ;
        RECT 37.320 201.850 37.640 201.910 ;
        RECT 38.155 201.865 38.445 201.910 ;
        RECT 38.700 202.050 39.020 202.110 ;
        RECT 40.170 202.050 40.310 202.205 ;
        RECT 38.700 201.910 40.310 202.050 ;
        RECT 41.090 202.050 41.230 202.205 ;
        RECT 49.740 202.190 50.105 202.410 ;
        RECT 51.580 202.190 51.900 202.450 ;
        RECT 52.975 202.390 53.265 202.435 ;
        RECT 53.420 202.390 53.740 202.450 ;
        RECT 55.810 202.435 55.950 202.590 ;
        RECT 59.490 202.590 61.085 202.730 ;
        RECT 52.975 202.250 53.740 202.390 ;
        RECT 52.975 202.205 53.265 202.250 ;
        RECT 53.420 202.190 53.740 202.250 ;
        RECT 54.355 202.390 54.645 202.435 ;
        RECT 54.355 202.250 55.030 202.390 ;
        RECT 54.355 202.205 54.645 202.250 ;
        RECT 42.840 202.050 43.160 202.110 ;
        RECT 49.815 202.095 50.105 202.190 ;
        RECT 41.090 201.910 43.160 202.050 ;
        RECT 38.700 201.850 39.020 201.910 ;
        RECT 42.840 201.850 43.160 201.910 ;
        RECT 44.235 201.865 44.525 202.095 ;
        RECT 46.515 202.050 47.165 202.095 ;
        RECT 49.815 202.050 50.405 202.095 ;
        RECT 46.515 201.910 50.405 202.050 ;
        RECT 51.670 202.050 51.810 202.190 ;
        RECT 53.895 202.050 54.185 202.095 ;
        RECT 51.670 201.910 54.185 202.050 ;
        RECT 46.515 201.865 47.165 201.910 ;
        RECT 50.115 201.865 50.405 201.910 ;
        RECT 18.090 201.570 22.830 201.710 ;
        RECT 23.060 201.510 23.380 201.770 ;
        RECT 23.980 201.710 24.300 201.770 ;
        RECT 25.835 201.710 26.125 201.755 ;
        RECT 23.980 201.570 26.125 201.710 ;
        RECT 23.980 201.510 24.300 201.570 ;
        RECT 25.835 201.525 26.125 201.570 ;
        RECT 26.280 201.510 26.600 201.770 ;
        RECT 29.960 201.510 30.280 201.770 ;
        RECT 35.940 201.710 36.260 201.770 ;
        RECT 39.160 201.710 39.480 201.770 ;
        RECT 39.635 201.710 39.925 201.755 ;
        RECT 35.940 201.570 39.925 201.710 ;
        RECT 44.310 201.710 44.450 201.865 ;
        RECT 53.050 201.770 53.190 201.910 ;
        RECT 53.895 201.865 54.185 201.910 ;
        RECT 54.890 201.770 55.030 202.250 ;
        RECT 55.735 202.205 56.025 202.435 ;
        RECT 57.100 202.190 57.420 202.450 ;
        RECT 58.020 202.190 58.340 202.450 ;
        RECT 58.495 202.390 58.785 202.435 ;
        RECT 58.940 202.390 59.260 202.450 ;
        RECT 58.495 202.250 59.260 202.390 ;
        RECT 58.495 202.205 58.785 202.250 ;
        RECT 58.940 202.190 59.260 202.250 ;
        RECT 59.490 202.050 59.630 202.590 ;
        RECT 60.795 202.545 61.085 202.590 ;
        RECT 61.255 202.545 61.545 202.775 ;
        RECT 62.635 202.545 62.925 202.775 ;
        RECT 59.875 202.390 60.165 202.435 ;
        RECT 62.710 202.390 62.850 202.545 ;
        RECT 59.875 202.250 62.850 202.390 ;
        RECT 63.095 202.390 63.385 202.435 ;
        RECT 63.630 202.390 63.770 202.930 ;
        RECT 64.920 202.870 65.240 202.930 ;
        RECT 65.470 202.930 74.425 203.070 ;
        RECT 65.470 202.730 65.610 202.930 ;
        RECT 74.135 202.885 74.425 202.930 ;
        RECT 75.500 202.870 75.820 203.130 ;
        RECT 75.960 203.070 76.280 203.130 ;
        RECT 97.210 203.070 97.350 203.270 ;
        RECT 97.580 203.210 97.900 203.470 ;
        RECT 98.040 203.210 98.360 203.470 ;
        RECT 102.180 203.210 102.500 203.470 ;
        RECT 103.560 203.410 103.880 203.470 ;
        RECT 111.840 203.410 112.160 203.470 ;
        RECT 120.135 203.410 120.425 203.455 ;
        RECT 120.580 203.410 120.900 203.470 ;
        RECT 103.560 203.270 112.160 203.410 ;
        RECT 103.560 203.210 103.880 203.270 ;
        RECT 111.840 203.210 112.160 203.270 ;
        RECT 112.390 203.270 120.900 203.410 ;
        RECT 112.390 203.130 112.530 203.270 ;
        RECT 120.135 203.225 120.425 203.270 ;
        RECT 120.580 203.210 120.900 203.270 ;
        RECT 122.420 203.410 122.740 203.470 ;
        RECT 123.815 203.410 124.105 203.455 ;
        RECT 122.420 203.270 124.105 203.410 ;
        RECT 122.420 203.210 122.740 203.270 ;
        RECT 123.815 203.225 124.105 203.270 ;
        RECT 124.260 203.410 124.580 203.470 ;
        RECT 124.735 203.410 125.025 203.455 ;
        RECT 130.700 203.410 131.020 203.470 ;
        RECT 124.260 203.270 131.020 203.410 ;
        RECT 124.260 203.210 124.580 203.270 ;
        RECT 124.735 203.225 125.025 203.270 ;
        RECT 130.700 203.210 131.020 203.270 ;
        RECT 133.460 203.410 133.780 203.470 ;
        RECT 137.615 203.410 137.905 203.455 ;
        RECT 133.460 203.270 137.905 203.410 ;
        RECT 133.460 203.210 133.780 203.270 ;
        RECT 137.615 203.225 137.905 203.270 ;
        RECT 146.340 203.410 146.660 203.470 ;
        RECT 146.815 203.410 147.105 203.455 ;
        RECT 147.720 203.410 148.040 203.470 ;
        RECT 146.340 203.270 148.040 203.410 ;
        RECT 146.340 203.210 146.660 203.270 ;
        RECT 146.815 203.225 147.105 203.270 ;
        RECT 147.720 203.210 148.040 203.270 ;
        RECT 150.940 203.210 151.260 203.470 ;
        RECT 152.320 203.210 152.640 203.470 ;
        RECT 101.260 203.070 101.580 203.130 ;
        RECT 75.960 202.930 96.350 203.070 ;
        RECT 97.210 202.930 102.410 203.070 ;
        RECT 75.960 202.870 76.280 202.930 ;
        RECT 63.095 202.250 63.770 202.390 ;
        RECT 64.090 202.590 65.610 202.730 ;
        RECT 65.855 202.730 66.145 202.775 ;
        RECT 70.455 202.730 70.745 202.775 ;
        RECT 65.855 202.590 70.745 202.730 ;
        RECT 59.875 202.205 60.165 202.250 ;
        RECT 63.095 202.205 63.385 202.250 ;
        RECT 61.700 202.050 62.020 202.110 ;
        RECT 64.090 202.050 64.230 202.590 ;
        RECT 65.855 202.545 66.145 202.590 ;
        RECT 70.455 202.545 70.745 202.590 ;
        RECT 71.835 202.730 72.125 202.775 ;
        RECT 75.590 202.730 75.730 202.870 ;
        RECT 71.835 202.590 75.730 202.730 ;
        RECT 71.835 202.545 72.125 202.590 ;
        RECT 64.475 202.205 64.765 202.435 ;
        RECT 64.935 202.390 65.225 202.435 ;
        RECT 66.300 202.390 66.620 202.450 ;
        RECT 64.935 202.250 66.620 202.390 ;
        RECT 64.935 202.205 65.225 202.250 ;
        RECT 59.490 201.910 64.230 202.050 ;
        RECT 64.550 202.050 64.690 202.205 ;
        RECT 66.300 202.190 66.620 202.250 ;
        RECT 69.520 202.190 69.840 202.450 ;
        RECT 69.995 202.205 70.285 202.435 ;
        RECT 70.915 202.390 71.205 202.435 ;
        RECT 72.295 202.390 72.585 202.435 ;
        RECT 70.915 202.250 72.585 202.390 ;
        RECT 70.915 202.205 71.205 202.250 ;
        RECT 72.295 202.205 72.585 202.250 ;
        RECT 70.070 202.050 70.210 202.205 ;
        RECT 73.200 202.190 73.520 202.450 ;
        RECT 73.675 202.205 73.965 202.435 ;
        RECT 73.750 202.050 73.890 202.205 ;
        RECT 74.580 202.190 74.900 202.450 ;
        RECT 75.040 202.190 75.360 202.450 ;
        RECT 76.050 202.435 76.190 202.870 ;
        RECT 79.195 202.545 79.485 202.775 ;
        RECT 80.560 202.730 80.880 202.790 ;
        RECT 94.820 202.730 95.140 202.790 ;
        RECT 80.560 202.590 94.590 202.730 ;
        RECT 75.975 202.205 76.265 202.435 ;
        RECT 76.880 202.190 77.200 202.450 ;
        RECT 77.340 202.190 77.660 202.450 ;
        RECT 77.815 202.390 78.105 202.435 ;
        RECT 78.260 202.390 78.580 202.450 ;
        RECT 77.815 202.250 78.580 202.390 ;
        RECT 79.270 202.390 79.410 202.545 ;
        RECT 80.560 202.530 80.880 202.590 ;
        RECT 79.655 202.390 79.945 202.435 ;
        RECT 79.270 202.250 79.945 202.390 ;
        RECT 77.815 202.205 78.105 202.250 ;
        RECT 78.260 202.190 78.580 202.250 ;
        RECT 79.655 202.205 79.945 202.250 ;
        RECT 80.100 202.190 80.420 202.450 ;
        RECT 81.035 202.390 81.325 202.435 ;
        RECT 81.035 202.250 84.010 202.390 ;
        RECT 81.035 202.205 81.325 202.250 ;
        RECT 75.130 202.050 75.270 202.190 ;
        RECT 64.550 201.910 67.450 202.050 ;
        RECT 70.070 201.910 72.510 202.050 ;
        RECT 73.750 201.910 75.270 202.050 ;
        RECT 76.970 202.050 77.110 202.190 ;
        RECT 83.870 202.110 84.010 202.250 ;
        RECT 84.240 202.190 84.560 202.450 ;
        RECT 84.700 202.390 85.020 202.450 ;
        RECT 85.635 202.390 85.925 202.435 ;
        RECT 84.700 202.250 85.925 202.390 ;
        RECT 84.700 202.190 85.020 202.250 ;
        RECT 85.635 202.205 85.925 202.250 ;
        RECT 86.080 202.390 86.400 202.450 ;
        RECT 89.300 202.390 89.620 202.450 ;
        RECT 86.080 202.250 89.620 202.390 ;
        RECT 86.080 202.190 86.400 202.250 ;
        RECT 89.300 202.190 89.620 202.250 ;
        RECT 93.440 202.390 93.760 202.450 ;
        RECT 94.450 202.435 94.590 202.590 ;
        RECT 94.820 202.590 95.970 202.730 ;
        RECT 94.820 202.530 95.140 202.590 ;
        RECT 93.915 202.390 94.205 202.435 ;
        RECT 93.440 202.250 94.205 202.390 ;
        RECT 93.440 202.190 93.760 202.250 ;
        RECT 93.915 202.205 94.205 202.250 ;
        RECT 94.375 202.205 94.665 202.435 ;
        RECT 95.280 202.190 95.600 202.450 ;
        RECT 95.830 202.435 95.970 202.590 ;
        RECT 95.755 202.205 96.045 202.435 ;
        RECT 96.210 202.390 96.350 202.930 ;
        RECT 101.260 202.870 101.580 202.930 ;
        RECT 102.270 202.775 102.410 202.930 ;
        RECT 103.100 202.870 103.420 203.130 ;
        RECT 104.020 202.870 104.340 203.130 ;
        RECT 106.320 203.070 106.640 203.130 ;
        RECT 112.300 203.070 112.620 203.130 ;
        RECT 115.060 203.070 115.380 203.130 ;
        RECT 106.320 202.930 112.620 203.070 ;
        RECT 106.320 202.870 106.640 202.930 ;
        RECT 112.300 202.870 112.620 202.930 ;
        RECT 113.310 202.930 115.380 203.070 ;
        RECT 96.675 202.770 96.965 202.775 ;
        RECT 97.115 202.770 97.405 202.775 ;
        RECT 96.675 202.630 97.405 202.770 ;
        RECT 96.675 202.545 96.965 202.630 ;
        RECT 97.115 202.545 97.405 202.630 ;
        RECT 97.670 202.590 100.110 202.730 ;
        RECT 97.670 202.390 97.810 202.590 ;
        RECT 98.500 202.390 98.820 202.450 ;
        RECT 96.210 202.250 97.810 202.390 ;
        RECT 98.130 202.250 98.820 202.390 ;
        RECT 99.970 202.390 100.110 202.590 ;
        RECT 102.195 202.545 102.485 202.775 ;
        RECT 103.190 202.730 103.330 202.870 ;
        RECT 103.190 202.590 103.790 202.730 ;
        RECT 102.730 202.435 103.330 202.440 ;
        RECT 102.730 202.400 103.405 202.435 ;
        RECT 102.330 202.390 103.405 202.400 ;
        RECT 99.970 202.300 103.405 202.390 ;
        RECT 99.970 202.260 102.870 202.300 ;
        RECT 99.970 202.250 102.470 202.260 ;
        RECT 76.970 201.910 83.090 202.050 ;
        RECT 61.700 201.850 62.020 201.910 ;
        RECT 67.310 201.770 67.450 201.910 ;
        RECT 48.360 201.710 48.680 201.770 ;
        RECT 44.310 201.570 48.680 201.710 ;
        RECT 35.940 201.510 36.260 201.570 ;
        RECT 39.160 201.510 39.480 201.570 ;
        RECT 39.635 201.525 39.925 201.570 ;
        RECT 48.360 201.510 48.680 201.570 ;
        RECT 52.040 201.510 52.360 201.770 ;
        RECT 52.960 201.510 53.280 201.770 ;
        RECT 54.800 201.510 55.120 201.770 ;
        RECT 59.860 201.710 60.180 201.770 ;
        RECT 63.555 201.710 63.845 201.755 ;
        RECT 59.860 201.570 63.845 201.710 ;
        RECT 59.860 201.510 60.180 201.570 ;
        RECT 63.555 201.525 63.845 201.570 ;
        RECT 67.220 201.510 67.540 201.770 ;
        RECT 72.370 201.710 72.510 201.910 ;
        RECT 82.950 201.770 83.090 201.910 ;
        RECT 83.780 201.850 84.100 202.110 ;
        RECT 88.380 202.050 88.700 202.110 ;
        RECT 96.660 202.050 96.980 202.110 ;
        RECT 98.130 202.050 98.270 202.250 ;
        RECT 98.500 202.190 98.820 202.250 ;
        RECT 88.380 201.910 96.350 202.050 ;
        RECT 88.380 201.850 88.700 201.910 ;
        RECT 79.655 201.710 79.945 201.755 ;
        RECT 72.370 201.570 79.945 201.710 ;
        RECT 79.655 201.525 79.945 201.570 ;
        RECT 80.100 201.710 80.420 201.770 ;
        RECT 82.400 201.710 82.720 201.770 ;
        RECT 80.100 201.570 82.720 201.710 ;
        RECT 80.100 201.510 80.420 201.570 ;
        RECT 82.400 201.510 82.720 201.570 ;
        RECT 82.860 201.510 83.180 201.770 ;
        RECT 86.080 201.710 86.400 201.770 ;
        RECT 87.920 201.710 88.240 201.770 ;
        RECT 86.080 201.570 88.240 201.710 ;
        RECT 86.080 201.510 86.400 201.570 ;
        RECT 87.920 201.510 88.240 201.570 ;
        RECT 92.520 201.710 92.840 201.770 ;
        RECT 95.740 201.710 96.060 201.770 ;
        RECT 92.520 201.570 96.060 201.710 ;
        RECT 96.210 201.710 96.350 201.910 ;
        RECT 96.660 201.910 98.270 202.050 ;
        RECT 100.340 202.050 100.660 202.110 ;
        RECT 101.735 202.050 102.025 202.095 ;
        RECT 100.340 201.910 102.025 202.050 ;
        RECT 102.730 202.050 102.870 202.260 ;
        RECT 103.115 202.205 103.405 202.300 ;
        RECT 103.650 202.390 103.790 202.590 ;
        RECT 113.310 202.435 113.450 202.930 ;
        RECT 115.060 202.870 115.380 202.930 ;
        RECT 115.995 203.070 116.285 203.115 ;
        RECT 129.320 203.070 129.640 203.130 ;
        RECT 115.995 202.930 129.640 203.070 ;
        RECT 115.995 202.885 116.285 202.930 ;
        RECT 129.320 202.870 129.640 202.930 ;
        RECT 131.160 203.070 131.480 203.130 ;
        RECT 140.360 203.070 140.680 203.130 ;
        RECT 131.160 202.930 140.680 203.070 ;
        RECT 131.160 202.870 131.480 202.930 ;
        RECT 113.680 202.530 114.000 202.790 ;
        RECT 115.520 202.730 115.840 202.790 ;
        RECT 121.500 202.730 121.820 202.790 ;
        RECT 115.520 202.590 121.820 202.730 ;
        RECT 115.520 202.530 115.840 202.590 ;
        RECT 121.500 202.530 121.820 202.590 ;
        RECT 122.420 202.730 122.740 202.790 ;
        RECT 123.355 202.730 123.645 202.775 ;
        RECT 125.195 202.730 125.485 202.775 ;
        RECT 122.420 202.590 125.485 202.730 ;
        RECT 122.420 202.530 122.740 202.590 ;
        RECT 123.355 202.545 123.645 202.590 ;
        RECT 125.195 202.545 125.485 202.590 ;
        RECT 133.475 202.730 133.765 202.775 ;
        RECT 136.220 202.730 136.540 202.790 ;
        RECT 133.475 202.590 136.540 202.730 ;
        RECT 133.475 202.545 133.765 202.590 ;
        RECT 136.220 202.530 136.540 202.590 ;
        RECT 136.680 202.730 137.000 202.790 ;
        RECT 136.680 202.590 137.600 202.730 ;
        RECT 136.680 202.530 137.000 202.590 ;
        RECT 113.235 202.390 113.525 202.435 ;
        RECT 103.650 202.250 113.525 202.390 ;
        RECT 113.235 202.205 113.525 202.250 ;
        RECT 114.140 202.390 114.460 202.450 ;
        RECT 114.615 202.390 114.905 202.435 ;
        RECT 114.140 202.250 114.905 202.390 ;
        RECT 114.140 202.190 114.460 202.250 ;
        RECT 114.615 202.205 114.905 202.250 ;
        RECT 115.060 202.190 115.380 202.450 ;
        RECT 117.360 202.390 117.680 202.450 ;
        RECT 118.740 202.390 119.060 202.450 ;
        RECT 119.675 202.390 119.965 202.435 ;
        RECT 117.360 202.250 119.965 202.390 ;
        RECT 117.360 202.190 117.680 202.250 ;
        RECT 118.740 202.190 119.060 202.250 ;
        RECT 119.675 202.205 119.965 202.250 ;
        RECT 120.120 202.390 120.440 202.450 ;
        RECT 121.975 202.390 122.265 202.435 ;
        RECT 120.120 202.250 122.265 202.390 ;
        RECT 120.120 202.190 120.440 202.250 ;
        RECT 121.975 202.205 122.265 202.250 ;
        RECT 124.260 202.390 124.580 202.450 ;
        RECT 124.735 202.390 125.025 202.435 ;
        RECT 124.260 202.250 125.025 202.390 ;
        RECT 124.260 202.190 124.580 202.250 ;
        RECT 124.735 202.205 125.025 202.250 ;
        RECT 126.115 202.390 126.405 202.435 ;
        RECT 126.115 202.250 136.910 202.390 ;
        RECT 137.460 202.265 137.600 202.590 ;
        RECT 126.115 202.205 126.405 202.250 ;
        RECT 120.210 202.050 120.350 202.190 ;
        RECT 102.730 201.910 120.350 202.050 ;
        RECT 121.055 202.050 121.345 202.095 ;
        RECT 123.340 202.050 123.660 202.110 ;
        RECT 127.020 202.050 127.340 202.110 ;
        RECT 128.400 202.050 128.720 202.110 ;
        RECT 121.055 201.910 123.660 202.050 ;
        RECT 96.660 201.850 96.980 201.910 ;
        RECT 100.340 201.850 100.660 201.910 ;
        RECT 101.735 201.865 102.025 201.910 ;
        RECT 121.055 201.865 121.345 201.910 ;
        RECT 123.340 201.850 123.660 201.910 ;
        RECT 124.350 201.910 128.720 202.050 ;
        RECT 104.940 201.710 105.260 201.770 ;
        RECT 109.540 201.710 109.860 201.770 ;
        RECT 96.210 201.570 109.860 201.710 ;
        RECT 92.520 201.510 92.840 201.570 ;
        RECT 95.740 201.510 96.060 201.570 ;
        RECT 104.940 201.510 105.260 201.570 ;
        RECT 109.540 201.510 109.860 201.570 ;
        RECT 121.515 201.710 121.805 201.755 ;
        RECT 124.350 201.710 124.490 201.910 ;
        RECT 127.020 201.850 127.340 201.910 ;
        RECT 128.400 201.850 128.720 201.910 ;
        RECT 129.320 202.050 129.640 202.110 ;
        RECT 133.475 202.050 133.765 202.095 ;
        RECT 129.320 201.910 133.765 202.050 ;
        RECT 129.320 201.850 129.640 201.910 ;
        RECT 133.475 201.865 133.765 201.910 ;
        RECT 133.935 202.050 134.225 202.095 ;
        RECT 134.840 202.050 135.160 202.110 ;
        RECT 133.935 201.910 135.160 202.050 ;
        RECT 133.935 201.865 134.225 201.910 ;
        RECT 134.840 201.850 135.160 201.910 ;
        RECT 121.515 201.570 124.490 201.710 ;
        RECT 126.100 201.710 126.420 201.770 ;
        RECT 136.770 201.755 136.910 202.250 ;
        RECT 137.385 202.035 137.675 202.265 ;
        RECT 138.150 202.050 138.290 202.930 ;
        RECT 140.360 202.870 140.680 202.930 ;
        RECT 151.030 202.730 151.170 203.210 ;
        RECT 151.875 202.730 152.165 202.775 ;
        RECT 151.030 202.590 152.165 202.730 ;
        RECT 152.410 202.730 152.550 203.210 ;
        RECT 152.795 202.730 153.085 202.775 ;
        RECT 152.410 202.590 153.085 202.730 ;
        RECT 151.875 202.545 152.165 202.590 ;
        RECT 152.795 202.545 153.085 202.590 ;
        RECT 143.120 202.390 143.440 202.450 ;
        RECT 150.480 202.390 150.800 202.450 ;
        RECT 152.335 202.390 152.625 202.435 ;
        RECT 143.120 202.250 152.625 202.390 ;
        RECT 143.120 202.190 143.440 202.250 ;
        RECT 150.480 202.190 150.800 202.250 ;
        RECT 152.335 202.205 152.625 202.250 ;
        RECT 153.240 202.190 153.560 202.450 ;
        RECT 138.535 202.050 138.825 202.095 ;
        RECT 138.150 201.910 138.825 202.050 ;
        RECT 138.535 201.865 138.825 201.910 ;
        RECT 138.980 202.050 139.300 202.110 ;
        RECT 145.435 202.050 145.725 202.095 ;
        RECT 150.020 202.050 150.340 202.110 ;
        RECT 138.980 201.910 150.340 202.050 ;
        RECT 138.980 201.850 139.300 201.910 ;
        RECT 145.435 201.865 145.725 201.910 ;
        RECT 150.020 201.850 150.340 201.910 ;
        RECT 131.085 201.710 131.375 201.755 ;
        RECT 126.100 201.570 131.375 201.710 ;
        RECT 121.515 201.525 121.805 201.570 ;
        RECT 126.100 201.510 126.420 201.570 ;
        RECT 131.085 201.525 131.375 201.570 ;
        RECT 136.695 201.525 136.985 201.755 ;
        RECT 150.955 201.710 151.245 201.755 ;
        RECT 152.320 201.710 152.640 201.770 ;
        RECT 150.955 201.570 152.640 201.710 ;
        RECT 150.955 201.525 151.245 201.570 ;
        RECT 152.320 201.510 152.640 201.570 ;
        RECT 2.750 200.890 159.030 201.370 ;
        RECT 13.860 200.690 14.180 200.750 ;
        RECT 18.920 200.690 19.240 200.750 ;
        RECT 4.290 200.550 13.630 200.690 ;
        RECT 4.290 200.055 4.430 200.550 ;
        RECT 7.875 200.350 8.525 200.395 ;
        RECT 11.475 200.350 11.765 200.395 ;
        RECT 12.940 200.350 13.260 200.410 ;
        RECT 7.875 200.210 13.260 200.350 ;
        RECT 7.875 200.165 8.525 200.210 ;
        RECT 11.175 200.165 11.765 200.210 ;
        RECT 4.215 199.825 4.505 200.055 ;
        RECT 4.680 200.010 4.970 200.055 ;
        RECT 6.515 200.010 6.805 200.055 ;
        RECT 10.095 200.010 10.385 200.055 ;
        RECT 4.680 199.870 10.385 200.010 ;
        RECT 4.680 199.825 4.970 199.870 ;
        RECT 6.515 199.825 6.805 199.870 ;
        RECT 10.095 199.825 10.385 199.870 ;
        RECT 11.175 199.850 11.465 200.165 ;
        RECT 12.940 200.150 13.260 200.210 ;
        RECT 13.490 200.070 13.630 200.550 ;
        RECT 13.860 200.550 19.240 200.690 ;
        RECT 13.860 200.490 14.180 200.550 ;
        RECT 18.920 200.490 19.240 200.550 ;
        RECT 19.840 200.690 20.160 200.750 ;
        RECT 29.040 200.690 29.360 200.750 ;
        RECT 31.355 200.690 31.645 200.735 ;
        RECT 34.100 200.690 34.420 200.750 ;
        RECT 38.700 200.690 39.020 200.750 ;
        RECT 19.840 200.550 20.530 200.690 ;
        RECT 19.840 200.490 20.160 200.550 ;
        RECT 17.075 200.350 17.725 200.395 ;
        RECT 20.390 200.350 20.530 200.550 ;
        RECT 29.040 200.550 31.645 200.690 ;
        RECT 29.040 200.490 29.360 200.550 ;
        RECT 31.355 200.505 31.645 200.550 ;
        RECT 31.890 200.550 39.020 200.690 ;
        RECT 20.675 200.350 20.965 200.395 ;
        RECT 17.075 200.210 20.965 200.350 ;
        RECT 17.075 200.165 17.725 200.210 ;
        RECT 20.375 200.165 20.965 200.210 ;
        RECT 22.600 200.350 22.920 200.410 ;
        RECT 28.120 200.350 28.440 200.410 ;
        RECT 31.890 200.350 32.030 200.550 ;
        RECT 34.100 200.490 34.420 200.550 ;
        RECT 38.700 200.490 39.020 200.550 ;
        RECT 39.175 200.690 39.465 200.735 ;
        RECT 40.080 200.690 40.400 200.750 ;
        RECT 43.300 200.690 43.620 200.750 ;
        RECT 45.140 200.690 45.460 200.750 ;
        RECT 39.175 200.550 40.400 200.690 ;
        RECT 39.175 200.505 39.465 200.550 ;
        RECT 40.080 200.490 40.400 200.550 ;
        RECT 42.010 200.550 43.620 200.690 ;
        RECT 22.600 200.210 25.590 200.350 ;
        RECT 13.400 199.810 13.720 200.070 ;
        RECT 13.880 200.010 14.170 200.055 ;
        RECT 15.715 200.010 16.005 200.055 ;
        RECT 19.295 200.010 19.585 200.055 ;
        RECT 13.880 199.870 19.585 200.010 ;
        RECT 13.880 199.825 14.170 199.870 ;
        RECT 15.715 199.825 16.005 199.870 ;
        RECT 19.295 199.825 19.585 199.870 ;
        RECT 20.375 199.850 20.665 200.165 ;
        RECT 22.600 200.150 22.920 200.210 ;
        RECT 22.140 200.010 22.460 200.070 ;
        RECT 25.450 200.055 25.590 200.210 ;
        RECT 28.120 200.210 32.030 200.350 ;
        RECT 33.195 200.350 33.485 200.395 ;
        RECT 35.940 200.350 36.260 200.410 ;
        RECT 33.195 200.210 36.260 200.350 ;
        RECT 28.120 200.150 28.440 200.210 ;
        RECT 33.195 200.165 33.485 200.210 ;
        RECT 35.940 200.150 36.260 200.210 ;
        RECT 40.935 200.350 41.225 200.395 ;
        RECT 41.460 200.350 41.780 200.410 ;
        RECT 42.010 200.395 42.150 200.550 ;
        RECT 43.300 200.490 43.620 200.550 ;
        RECT 44.335 200.550 45.460 200.690 ;
        RECT 44.335 200.395 44.475 200.550 ;
        RECT 45.140 200.490 45.460 200.550 ;
        RECT 45.690 200.550 48.590 200.690 ;
        RECT 40.935 200.210 41.780 200.350 ;
        RECT 40.935 200.165 41.225 200.210 ;
        RECT 41.460 200.150 41.780 200.210 ;
        RECT 41.935 200.165 42.225 200.395 ;
        RECT 42.470 200.210 43.530 200.350 ;
        RECT 23.995 200.010 24.285 200.055 ;
        RECT 22.140 199.870 24.285 200.010 ;
        RECT 22.140 199.810 22.460 199.870 ;
        RECT 23.995 199.825 24.285 199.870 ;
        RECT 24.455 199.825 24.745 200.055 ;
        RECT 25.375 199.825 25.665 200.055 ;
        RECT 30.435 199.825 30.725 200.055 ;
        RECT 33.655 200.010 33.945 200.055 ;
        RECT 36.875 200.010 37.165 200.055 ;
        RECT 33.655 199.870 37.165 200.010 ;
        RECT 33.655 199.825 33.945 199.870 ;
        RECT 36.875 199.825 37.165 199.870 ;
        RECT 5.580 199.470 5.900 199.730 ;
        RECT 14.780 199.470 15.100 199.730 ;
        RECT 19.840 199.670 20.160 199.730 ;
        RECT 24.530 199.670 24.670 199.825 ;
        RECT 19.840 199.530 24.670 199.670 ;
        RECT 27.200 199.670 27.520 199.730 ;
        RECT 27.675 199.670 27.965 199.715 ;
        RECT 27.200 199.530 27.965 199.670 ;
        RECT 19.840 199.470 20.160 199.530 ;
        RECT 27.200 199.470 27.520 199.530 ;
        RECT 27.675 199.485 27.965 199.530 ;
        RECT 5.085 199.330 5.375 199.375 ;
        RECT 6.975 199.330 7.265 199.375 ;
        RECT 10.095 199.330 10.385 199.375 ;
        RECT 5.085 199.190 10.385 199.330 ;
        RECT 5.085 199.145 5.375 199.190 ;
        RECT 6.975 199.145 7.265 199.190 ;
        RECT 10.095 199.145 10.385 199.190 ;
        RECT 14.285 199.330 14.575 199.375 ;
        RECT 16.175 199.330 16.465 199.375 ;
        RECT 19.295 199.330 19.585 199.375 ;
        RECT 30.510 199.330 30.650 199.825 ;
        RECT 32.260 199.670 32.580 199.730 ;
        RECT 33.730 199.670 33.870 199.825 ;
        RECT 37.320 199.810 37.640 200.070 ;
        RECT 42.470 200.055 42.610 200.210 ;
        RECT 40.630 199.870 41.690 200.010 ;
        RECT 32.260 199.530 33.870 199.670 ;
        RECT 34.115 199.670 34.405 199.715 ;
        RECT 35.480 199.670 35.800 199.730 ;
        RECT 34.115 199.530 35.800 199.670 ;
        RECT 32.260 199.470 32.580 199.530 ;
        RECT 34.115 199.485 34.405 199.530 ;
        RECT 35.480 199.470 35.800 199.530 ;
        RECT 36.400 199.470 36.720 199.730 ;
        RECT 40.630 199.330 40.770 199.870 ;
        RECT 14.285 199.190 19.585 199.330 ;
        RECT 14.285 199.145 14.575 199.190 ;
        RECT 16.175 199.145 16.465 199.190 ;
        RECT 19.295 199.145 19.585 199.190 ;
        RECT 19.930 199.190 24.670 199.330 ;
        RECT 30.510 199.190 40.770 199.330 ;
        RECT 12.955 198.990 13.245 199.035 ;
        RECT 15.240 198.990 15.560 199.050 ;
        RECT 18.460 198.990 18.780 199.050 ;
        RECT 19.930 198.990 20.070 199.190 ;
        RECT 24.530 199.050 24.670 199.190 ;
        RECT 12.955 198.850 20.070 198.990 ;
        RECT 22.155 198.990 22.445 199.035 ;
        RECT 23.520 198.990 23.840 199.050 ;
        RECT 22.155 198.850 23.840 198.990 ;
        RECT 12.955 198.805 13.245 198.850 ;
        RECT 15.240 198.790 15.560 198.850 ;
        RECT 18.460 198.790 18.780 198.850 ;
        RECT 22.155 198.805 22.445 198.850 ;
        RECT 23.520 198.790 23.840 198.850 ;
        RECT 24.440 198.790 24.760 199.050 ;
        RECT 29.500 198.790 29.820 199.050 ;
        RECT 33.640 198.990 33.960 199.050 ;
        RECT 39.160 198.990 39.480 199.050 ;
        RECT 40.095 198.990 40.385 199.035 ;
        RECT 33.640 198.850 40.385 198.990 ;
        RECT 33.640 198.790 33.960 198.850 ;
        RECT 39.160 198.790 39.480 198.850 ;
        RECT 40.095 198.805 40.385 198.850 ;
        RECT 41.000 198.790 41.320 199.050 ;
        RECT 41.550 198.990 41.690 199.870 ;
        RECT 42.395 199.825 42.685 200.055 ;
        RECT 42.860 199.825 43.150 200.055 ;
        RECT 42.930 199.670 43.070 199.825 ;
        RECT 42.475 199.530 43.070 199.670 ;
        RECT 43.390 199.670 43.530 200.210 ;
        RECT 44.235 200.165 44.525 200.395 ;
        RECT 43.760 199.810 44.080 200.070 ;
        RECT 44.925 200.010 45.215 200.055 ;
        RECT 45.690 200.010 45.830 200.550 ;
        RECT 46.980 200.350 47.300 200.410 ;
        RECT 47.455 200.350 47.745 200.395 ;
        RECT 46.980 200.210 47.745 200.350 ;
        RECT 46.980 200.150 47.300 200.210 ;
        RECT 47.455 200.165 47.745 200.210 ;
        RECT 44.925 199.870 45.830 200.010 ;
        RECT 44.925 199.825 45.215 199.870 ;
        RECT 46.060 199.810 46.380 200.070 ;
        RECT 46.540 199.825 46.830 200.055 ;
        RECT 46.150 199.670 46.290 199.810 ;
        RECT 43.390 199.530 46.290 199.670 ;
        RECT 46.615 199.670 46.755 199.825 ;
        RECT 47.900 199.810 48.220 200.070 ;
        RECT 48.450 200.055 48.590 200.550 ;
        RECT 49.740 200.490 50.060 200.750 ;
        RECT 52.040 200.690 52.360 200.750 ;
        RECT 51.670 200.550 52.360 200.690 ;
        RECT 49.280 200.350 49.600 200.410 ;
        RECT 51.670 200.395 51.810 200.550 ;
        RECT 52.040 200.490 52.360 200.550 ;
        RECT 52.960 200.690 53.280 200.750 ;
        RECT 61.700 200.735 62.020 200.750 ;
        RECT 59.415 200.690 59.705 200.735 ;
        RECT 61.680 200.690 62.020 200.735 ;
        RECT 82.860 200.690 83.180 200.750 ;
        RECT 52.960 200.550 59.705 200.690 ;
        RECT 61.505 200.550 62.020 200.690 ;
        RECT 52.960 200.490 53.280 200.550 ;
        RECT 49.280 200.210 51.350 200.350 ;
        RECT 49.280 200.150 49.600 200.210 ;
        RECT 50.660 200.055 50.980 200.070 ;
        RECT 51.210 200.055 51.350 200.210 ;
        RECT 51.595 200.165 51.885 200.395 ;
        RECT 54.800 200.350 55.120 200.410 ;
        RECT 56.730 200.395 56.870 200.550 ;
        RECT 59.415 200.505 59.705 200.550 ;
        RECT 61.680 200.505 62.020 200.550 ;
        RECT 61.700 200.490 62.020 200.505 ;
        RECT 75.820 200.550 83.180 200.690 ;
        RECT 55.575 200.350 55.865 200.395 ;
        RECT 54.800 200.210 55.865 200.350 ;
        RECT 54.800 200.150 55.120 200.210 ;
        RECT 55.575 200.165 55.865 200.210 ;
        RECT 56.655 200.165 56.945 200.395 ;
        RECT 57.100 200.350 57.420 200.410 ;
        RECT 61.255 200.350 61.545 200.395 ;
        RECT 63.080 200.350 63.400 200.410 ;
        RECT 75.820 200.350 75.960 200.550 ;
        RECT 82.860 200.490 83.180 200.550 ;
        RECT 84.700 200.490 85.020 200.750 ;
        RECT 86.555 200.505 86.845 200.735 ;
        RECT 88.840 200.690 89.160 200.750 ;
        RECT 89.315 200.690 89.605 200.735 ;
        RECT 92.520 200.690 92.840 200.750 ;
        RECT 88.840 200.550 89.605 200.690 ;
        RECT 86.630 200.350 86.770 200.505 ;
        RECT 88.840 200.490 89.160 200.550 ;
        RECT 89.315 200.505 89.605 200.550 ;
        RECT 89.850 200.550 92.840 200.690 ;
        RECT 89.850 200.350 89.990 200.550 ;
        RECT 92.520 200.490 92.840 200.550 ;
        RECT 93.440 200.690 93.760 200.750 ;
        RECT 93.440 200.550 97.810 200.690 ;
        RECT 93.440 200.490 93.760 200.550 ;
        RECT 57.100 200.210 61.010 200.350 ;
        RECT 57.100 200.150 57.420 200.210 ;
        RECT 48.400 199.960 48.690 200.055 ;
        RECT 50.650 200.010 50.980 200.055 ;
        RECT 49.370 199.960 50.980 200.010 ;
        RECT 48.400 199.870 50.980 199.960 ;
        RECT 48.400 199.825 49.510 199.870 ;
        RECT 50.650 199.825 50.980 199.870 ;
        RECT 51.135 199.825 51.425 200.055 ;
        RECT 52.500 200.010 52.820 200.070 ;
        RECT 52.305 199.870 52.820 200.010 ;
        RECT 48.450 199.820 49.510 199.825 ;
        RECT 50.660 199.810 50.980 199.825 ;
        RECT 52.500 199.810 52.820 199.870 ;
        RECT 52.960 199.810 53.280 200.070 ;
        RECT 53.880 200.010 54.200 200.070 ;
        RECT 58.495 200.010 58.785 200.055 ;
        RECT 53.880 199.870 58.785 200.010 ;
        RECT 53.880 199.810 54.200 199.870 ;
        RECT 58.495 199.825 58.785 199.870 ;
        RECT 58.940 199.810 59.260 200.070 ;
        RECT 59.860 200.010 60.180 200.070 ;
        RECT 60.870 200.055 61.010 200.210 ;
        RECT 61.255 200.210 75.960 200.350 ;
        RECT 83.870 200.210 89.990 200.350 ;
        RECT 94.820 200.350 95.140 200.410 ;
        RECT 94.820 200.210 96.430 200.350 ;
        RECT 61.255 200.165 61.545 200.210 ;
        RECT 63.080 200.150 63.400 200.210 ;
        RECT 60.335 200.010 60.625 200.055 ;
        RECT 59.860 199.870 60.625 200.010 ;
        RECT 59.860 199.810 60.180 199.870 ;
        RECT 60.335 199.825 60.625 199.870 ;
        RECT 60.795 199.825 61.085 200.055 ;
        RECT 62.160 200.010 62.480 200.070 ;
        RECT 67.680 200.010 68.000 200.070 ;
        RECT 62.160 199.870 68.000 200.010 ;
        RECT 46.615 199.530 60.550 199.670 ;
        RECT 42.475 199.390 42.615 199.530 ;
        RECT 42.380 199.130 42.700 199.390 ;
        RECT 45.615 199.330 45.905 199.375 ;
        RECT 47.440 199.330 47.760 199.390 ;
        RECT 51.120 199.330 51.440 199.390 ;
        RECT 45.615 199.190 47.760 199.330 ;
        RECT 45.615 199.145 45.905 199.190 ;
        RECT 47.440 199.130 47.760 199.190 ;
        RECT 49.370 199.190 51.440 199.330 ;
        RECT 43.300 198.990 43.620 199.050 ;
        RECT 49.370 199.035 49.510 199.190 ;
        RECT 51.120 199.130 51.440 199.190 ;
        RECT 53.420 199.330 53.740 199.390 ;
        RECT 56.180 199.330 56.500 199.390 ;
        RECT 60.410 199.375 60.550 199.530 ;
        RECT 57.575 199.330 57.865 199.375 ;
        RECT 53.420 199.190 55.950 199.330 ;
        RECT 53.420 199.130 53.740 199.190 ;
        RECT 41.550 198.850 43.620 198.990 ;
        RECT 43.300 198.790 43.620 198.850 ;
        RECT 49.295 198.805 49.585 199.035 ;
        RECT 54.340 198.990 54.660 199.050 ;
        RECT 55.810 199.035 55.950 199.190 ;
        RECT 56.180 199.190 57.865 199.330 ;
        RECT 56.180 199.130 56.500 199.190 ;
        RECT 57.575 199.145 57.865 199.190 ;
        RECT 60.335 199.145 60.625 199.375 ;
        RECT 54.815 198.990 55.105 199.035 ;
        RECT 54.340 198.850 55.105 198.990 ;
        RECT 54.340 198.790 54.660 198.850 ;
        RECT 54.815 198.805 55.105 198.850 ;
        RECT 55.735 198.805 56.025 199.035 ;
        RECT 59.860 198.990 60.180 199.050 ;
        RECT 60.870 198.990 61.010 199.825 ;
        RECT 62.160 199.810 62.480 199.870 ;
        RECT 67.680 199.810 68.000 199.870 ;
        RECT 68.140 200.010 68.460 200.070 ;
        RECT 83.320 200.010 83.640 200.070 ;
        RECT 83.870 200.010 84.010 200.210 ;
        RECT 94.820 200.150 95.140 200.210 ;
        RECT 68.140 199.870 84.010 200.010 ;
        RECT 68.140 199.810 68.460 199.870 ;
        RECT 83.320 199.810 83.640 199.870 ;
        RECT 86.095 199.825 86.385 200.055 ;
        RECT 86.540 200.010 86.860 200.070 ;
        RECT 87.015 200.010 87.305 200.055 ;
        RECT 86.540 199.870 87.305 200.010 ;
        RECT 64.000 199.670 64.320 199.730 ;
        RECT 66.760 199.670 67.080 199.730 ;
        RECT 81.020 199.670 81.340 199.730 ;
        RECT 64.000 199.530 81.340 199.670 ;
        RECT 86.170 199.670 86.310 199.825 ;
        RECT 86.540 199.810 86.860 199.870 ;
        RECT 87.015 199.825 87.305 199.870 ;
        RECT 87.460 200.010 87.780 200.070 ;
        RECT 87.935 200.010 88.225 200.055 ;
        RECT 87.460 199.870 88.225 200.010 ;
        RECT 87.460 199.810 87.780 199.870 ;
        RECT 87.935 199.825 88.225 199.870 ;
        RECT 88.395 200.010 88.685 200.055 ;
        RECT 89.300 200.010 89.620 200.070 ;
        RECT 88.395 199.870 89.620 200.010 ;
        RECT 88.395 199.825 88.685 199.870 ;
        RECT 89.300 199.810 89.620 199.870 ;
        RECT 89.775 199.825 90.065 200.055 ;
        RECT 90.695 200.010 90.985 200.055 ;
        RECT 94.360 200.010 94.680 200.070 ;
        RECT 95.740 200.010 96.060 200.070 ;
        RECT 96.290 200.055 96.430 200.210 ;
        RECT 97.120 200.150 97.440 200.410 ;
        RECT 97.670 200.395 97.810 200.550 ;
        RECT 98.960 200.490 99.280 200.750 ;
        RECT 107.700 200.690 108.020 200.750 ;
        RECT 116.440 200.690 116.760 200.750 ;
        RECT 99.740 200.550 116.760 200.690 ;
        RECT 97.595 200.350 97.885 200.395 ;
        RECT 99.740 200.350 99.880 200.550 ;
        RECT 107.700 200.490 108.020 200.550 ;
        RECT 116.440 200.490 116.760 200.550 ;
        RECT 117.360 200.690 117.680 200.750 ;
        RECT 119.755 200.690 120.045 200.735 ;
        RECT 117.360 200.550 120.045 200.690 ;
        RECT 117.360 200.490 117.680 200.550 ;
        RECT 119.755 200.505 120.045 200.550 ;
        RECT 120.595 200.505 120.885 200.735 ;
        RECT 125.180 200.690 125.500 200.750 ;
        RECT 125.655 200.690 125.945 200.735 ;
        RECT 125.180 200.550 125.945 200.690 ;
        RECT 97.595 200.210 99.880 200.350 ;
        RECT 100.800 200.350 101.120 200.410 ;
        RECT 104.020 200.350 104.340 200.410 ;
        RECT 100.800 200.210 103.790 200.350 ;
        RECT 97.595 200.165 97.885 200.210 ;
        RECT 100.800 200.150 101.120 200.210 ;
        RECT 103.650 200.070 103.790 200.210 ;
        RECT 104.020 200.210 107.470 200.350 ;
        RECT 104.020 200.150 104.340 200.210 ;
        RECT 90.695 199.870 94.680 200.010 ;
        RECT 90.695 199.825 90.985 199.870 ;
        RECT 89.850 199.670 89.990 199.825 ;
        RECT 94.360 199.810 94.680 199.870 ;
        RECT 94.910 199.870 96.060 200.010 ;
        RECT 94.910 199.670 95.050 199.870 ;
        RECT 95.740 199.810 96.060 199.870 ;
        RECT 96.215 199.825 96.505 200.055 ;
        RECT 98.040 199.810 98.360 200.070 ;
        RECT 98.960 200.010 99.280 200.070 ;
        RECT 99.435 200.010 99.725 200.055 ;
        RECT 98.960 199.870 99.725 200.010 ;
        RECT 98.960 199.810 99.280 199.870 ;
        RECT 99.435 199.825 99.725 199.870 ;
        RECT 99.895 199.825 100.185 200.055 ;
        RECT 100.430 199.870 103.330 200.010 ;
        RECT 86.170 199.530 87.690 199.670 ;
        RECT 89.850 199.530 91.370 199.670 ;
        RECT 64.000 199.470 64.320 199.530 ;
        RECT 66.760 199.470 67.080 199.530 ;
        RECT 81.020 199.470 81.340 199.530 ;
        RECT 87.550 199.390 87.690 199.530 ;
        RECT 91.230 199.390 91.370 199.530 ;
        RECT 94.450 199.530 95.050 199.670 ;
        RECT 97.120 199.670 97.440 199.730 ;
        RECT 99.970 199.670 100.110 199.825 ;
        RECT 97.120 199.530 100.110 199.670 ;
        RECT 69.980 199.330 70.300 199.390 ;
        RECT 69.980 199.190 87.230 199.330 ;
        RECT 69.980 199.130 70.300 199.190 ;
        RECT 59.860 198.850 61.010 198.990 ;
        RECT 70.440 198.990 70.760 199.050 ;
        RECT 75.960 198.990 76.280 199.050 ;
        RECT 70.440 198.850 76.280 198.990 ;
        RECT 87.090 198.990 87.230 199.190 ;
        RECT 87.460 199.130 87.780 199.390 ;
        RECT 91.140 199.130 91.460 199.390 ;
        RECT 94.450 198.990 94.590 199.530 ;
        RECT 97.120 199.470 97.440 199.530 ;
        RECT 96.660 199.330 96.980 199.390 ;
        RECT 100.430 199.330 100.570 199.870 ;
        RECT 102.640 199.470 102.960 199.730 ;
        RECT 103.190 199.670 103.330 199.870 ;
        RECT 103.560 199.810 103.880 200.070 ;
        RECT 107.330 200.055 107.470 200.210 ;
        RECT 108.160 200.150 108.480 200.410 ;
        RECT 115.980 200.150 116.300 200.410 ;
        RECT 117.820 200.350 118.140 200.410 ;
        RECT 118.755 200.350 119.045 200.395 ;
        RECT 117.820 200.210 119.045 200.350 ;
        RECT 117.820 200.150 118.140 200.210 ;
        RECT 118.755 200.165 119.045 200.210 ;
        RECT 107.255 199.825 107.545 200.055 ;
        RECT 107.715 199.825 108.005 200.055 ;
        RECT 104.020 199.670 104.340 199.730 ;
        RECT 103.190 199.530 104.340 199.670 ;
        RECT 104.020 199.470 104.340 199.530 ;
        RECT 104.940 199.670 105.260 199.730 ;
        RECT 107.790 199.670 107.930 199.825 ;
        RECT 109.080 199.810 109.400 200.070 ;
        RECT 109.555 200.010 109.845 200.055 ;
        RECT 116.070 200.010 116.210 200.150 ;
        RECT 109.555 199.870 116.210 200.010 ;
        RECT 109.555 199.825 109.845 199.870 ;
        RECT 104.940 199.530 107.930 199.670 ;
        RECT 119.830 199.670 119.970 200.505 ;
        RECT 120.670 200.350 120.810 200.505 ;
        RECT 125.180 200.490 125.500 200.550 ;
        RECT 125.655 200.505 125.945 200.550 ;
        RECT 135.300 200.690 135.620 200.750 ;
        RECT 140.360 200.690 140.680 200.750 ;
        RECT 135.300 200.550 143.350 200.690 ;
        RECT 135.300 200.490 135.620 200.550 ;
        RECT 140.360 200.490 140.680 200.550 ;
        RECT 121.055 200.350 121.345 200.395 ;
        RECT 120.670 200.210 121.345 200.350 ;
        RECT 121.055 200.165 121.345 200.210 ;
        RECT 121.975 200.350 122.265 200.395 ;
        RECT 123.355 200.350 123.645 200.395 ;
        RECT 130.240 200.350 130.560 200.410 ;
        RECT 142.200 200.350 142.520 200.410 ;
        RECT 142.675 200.350 142.965 200.395 ;
        RECT 121.975 200.210 123.645 200.350 ;
        RECT 121.975 200.165 122.265 200.210 ;
        RECT 123.355 200.165 123.645 200.210 ;
        RECT 124.350 200.210 130.560 200.350 ;
        RECT 124.350 200.070 124.490 200.210 ;
        RECT 130.240 200.150 130.560 200.210 ;
        RECT 132.170 200.210 142.965 200.350 ;
        RECT 143.210 200.350 143.350 200.550 ;
        RECT 144.500 200.490 144.820 200.750 ;
        RECT 149.560 200.490 149.880 200.750 ;
        RECT 145.435 200.350 145.725 200.395 ;
        RECT 143.210 200.210 145.725 200.350 ;
        RECT 132.170 200.070 132.310 200.210 ;
        RECT 142.200 200.150 142.520 200.210 ;
        RECT 142.675 200.165 142.965 200.210 ;
        RECT 145.435 200.165 145.725 200.210 ;
        RECT 145.880 200.350 146.200 200.410 ;
        RECT 146.355 200.350 146.645 200.395 ;
        RECT 145.880 200.210 146.645 200.350 ;
        RECT 145.880 200.150 146.200 200.210 ;
        RECT 146.355 200.165 146.645 200.210 ;
        RECT 122.420 199.810 122.740 200.070 ;
        RECT 122.895 199.825 123.185 200.055 ;
        RECT 121.500 199.670 121.820 199.730 ;
        RECT 122.970 199.670 123.110 199.825 ;
        RECT 124.260 199.810 124.580 200.070 ;
        RECT 126.560 200.010 126.880 200.070 ;
        RECT 128.415 200.010 128.705 200.055 ;
        RECT 126.560 199.870 128.705 200.010 ;
        RECT 126.560 199.810 126.880 199.870 ;
        RECT 128.415 199.825 128.705 199.870 ;
        RECT 128.860 200.010 129.180 200.070 ;
        RECT 129.795 200.010 130.085 200.055 ;
        RECT 128.860 199.870 130.085 200.010 ;
        RECT 128.860 199.810 129.180 199.870 ;
        RECT 129.795 199.825 130.085 199.870 ;
        RECT 132.080 199.810 132.400 200.070 ;
        RECT 132.540 199.810 132.860 200.070 ;
        RECT 133.000 200.010 133.320 200.070 ;
        RECT 133.000 199.870 135.530 200.010 ;
        RECT 133.000 199.810 133.320 199.870 ;
        RECT 119.830 199.530 123.110 199.670 ;
        RECT 125.655 199.670 125.945 199.715 ;
        RECT 127.495 199.670 127.785 199.715 ;
        RECT 132.630 199.670 132.770 199.810 ;
        RECT 134.395 199.670 134.685 199.715 ;
        RECT 125.655 199.530 127.785 199.670 ;
        RECT 104.940 199.470 105.260 199.530 ;
        RECT 121.500 199.470 121.820 199.530 ;
        RECT 125.655 199.485 125.945 199.530 ;
        RECT 127.495 199.485 127.785 199.530 ;
        RECT 127.950 199.530 134.685 199.670 ;
        RECT 96.660 199.190 100.570 199.330 ;
        RECT 100.815 199.330 101.105 199.375 ;
        RECT 102.730 199.330 102.870 199.470 ;
        RECT 114.600 199.330 114.920 199.390 ;
        RECT 100.815 199.190 102.870 199.330 ;
        RECT 103.190 199.190 114.920 199.330 ;
        RECT 96.660 199.130 96.980 199.190 ;
        RECT 100.815 199.145 101.105 199.190 ;
        RECT 87.090 198.850 94.590 198.990 ;
        RECT 95.740 198.990 96.060 199.050 ;
        RECT 103.190 198.990 103.330 199.190 ;
        RECT 114.600 199.130 114.920 199.190 ;
        RECT 121.055 199.330 121.345 199.375 ;
        RECT 124.735 199.330 125.025 199.375 ;
        RECT 121.055 199.190 125.025 199.330 ;
        RECT 121.055 199.145 121.345 199.190 ;
        RECT 124.735 199.145 125.025 199.190 ;
        RECT 95.740 198.850 103.330 198.990 ;
        RECT 59.860 198.790 60.180 198.850 ;
        RECT 70.440 198.790 70.760 198.850 ;
        RECT 75.960 198.790 76.280 198.850 ;
        RECT 95.740 198.790 96.060 198.850 ;
        RECT 106.320 198.790 106.640 199.050 ;
        RECT 111.380 198.990 111.700 199.050 ;
        RECT 119.660 198.990 119.980 199.050 ;
        RECT 111.380 198.850 119.980 198.990 ;
        RECT 111.380 198.790 111.700 198.850 ;
        RECT 119.660 198.790 119.980 198.850 ;
        RECT 124.260 198.990 124.580 199.050 ;
        RECT 127.950 198.990 128.090 199.530 ;
        RECT 134.395 199.485 134.685 199.530 ;
        RECT 128.860 199.130 129.180 199.390 ;
        RECT 129.335 199.330 129.625 199.375 ;
        RECT 132.095 199.330 132.385 199.375 ;
        RECT 129.335 199.190 132.385 199.330 ;
        RECT 135.390 199.330 135.530 199.870 ;
        RECT 141.740 199.810 142.060 200.070 ;
        RECT 143.135 200.010 143.425 200.055 ;
        RECT 142.750 199.870 143.425 200.010 ;
        RECT 142.750 199.730 142.890 199.870 ;
        RECT 143.135 199.825 143.425 199.870 ;
        RECT 143.580 199.810 143.900 200.070 ;
        RECT 144.975 199.825 145.265 200.055 ;
        RECT 142.660 199.470 142.980 199.730 ;
        RECT 143.120 199.330 143.440 199.390 ;
        RECT 135.390 199.190 143.440 199.330 ;
        RECT 129.335 199.145 129.625 199.190 ;
        RECT 132.095 199.145 132.385 199.190 ;
        RECT 143.120 199.130 143.440 199.190 ;
        RECT 124.260 198.850 128.090 198.990 ;
        RECT 132.540 198.990 132.860 199.050 ;
        RECT 133.935 198.990 134.225 199.035 ;
        RECT 134.840 198.990 135.160 199.050 ;
        RECT 132.540 198.850 135.160 198.990 ;
        RECT 145.050 198.990 145.190 199.825 ;
        RECT 150.940 199.810 151.260 200.070 ;
        RECT 151.415 199.825 151.705 200.055 ;
        RECT 151.875 199.825 152.165 200.055 ;
        RECT 152.320 200.010 152.640 200.070 ;
        RECT 152.795 200.010 153.085 200.055 ;
        RECT 152.320 199.870 153.085 200.010 ;
        RECT 151.490 199.670 151.630 199.825 ;
        RECT 146.430 199.530 151.630 199.670 ;
        RECT 146.430 199.375 146.570 199.530 ;
        RECT 146.355 199.145 146.645 199.375 ;
        RECT 151.400 199.330 151.720 199.390 ;
        RECT 151.950 199.330 152.090 199.825 ;
        RECT 152.320 199.810 152.640 199.870 ;
        RECT 152.795 199.825 153.085 199.870 ;
        RECT 151.400 199.190 152.090 199.330 ;
        RECT 151.400 199.130 151.720 199.190 ;
        RECT 147.260 198.990 147.580 199.050 ;
        RECT 145.050 198.850 147.580 198.990 ;
        RECT 124.260 198.790 124.580 198.850 ;
        RECT 132.540 198.790 132.860 198.850 ;
        RECT 133.935 198.805 134.225 198.850 ;
        RECT 134.840 198.790 135.160 198.850 ;
        RECT 147.260 198.790 147.580 198.850 ;
        RECT 2.750 198.170 158.230 198.650 ;
        RECT 5.580 197.970 5.900 198.030 ;
        RECT 6.055 197.970 6.345 198.015 ;
        RECT 5.580 197.830 6.345 197.970 ;
        RECT 5.580 197.770 5.900 197.830 ;
        RECT 6.055 197.785 6.345 197.830 ;
        RECT 14.780 197.970 15.100 198.030 ;
        RECT 16.175 197.970 16.465 198.015 ;
        RECT 14.780 197.830 16.465 197.970 ;
        RECT 14.780 197.770 15.100 197.830 ;
        RECT 16.175 197.785 16.465 197.830 ;
        RECT 17.080 197.970 17.400 198.030 ;
        RECT 24.455 197.970 24.745 198.015 ;
        RECT 17.080 197.830 24.745 197.970 ;
        RECT 17.080 197.770 17.400 197.830 ;
        RECT 24.455 197.785 24.745 197.830 ;
        RECT 26.755 197.970 27.045 198.015 ;
        RECT 28.120 197.970 28.440 198.030 ;
        RECT 26.755 197.830 28.440 197.970 ;
        RECT 26.755 197.785 27.045 197.830 ;
        RECT 14.320 197.630 14.640 197.690 ;
        RECT 23.520 197.630 23.840 197.690 ;
        RECT 14.320 197.490 23.840 197.630 ;
        RECT 14.320 197.430 14.640 197.490 ;
        RECT 23.520 197.430 23.840 197.490 ;
        RECT 10.640 197.090 10.960 197.350 ;
        RECT 12.495 197.290 12.785 197.335 ;
        RECT 20.300 197.290 20.620 197.350 ;
        RECT 26.830 197.290 26.970 197.785 ;
        RECT 28.120 197.770 28.440 197.830 ;
        RECT 28.990 197.970 29.280 198.015 ;
        RECT 29.500 197.970 29.820 198.030 ;
        RECT 28.990 197.830 29.820 197.970 ;
        RECT 28.990 197.785 29.280 197.830 ;
        RECT 29.500 197.770 29.820 197.830 ;
        RECT 40.540 197.770 40.860 198.030 ;
        RECT 41.000 197.770 41.320 198.030 ;
        RECT 43.760 197.770 44.080 198.030 ;
        RECT 44.235 197.970 44.525 198.015 ;
        RECT 44.680 197.970 45.000 198.030 ;
        RECT 44.235 197.830 45.000 197.970 ;
        RECT 44.235 197.785 44.525 197.830 ;
        RECT 44.680 197.770 45.000 197.830 ;
        RECT 48.360 197.770 48.680 198.030 ;
        RECT 50.660 197.970 50.980 198.030 ;
        RECT 52.040 197.970 52.360 198.030 ;
        RECT 50.660 197.830 52.360 197.970 ;
        RECT 50.660 197.770 50.980 197.830 ;
        RECT 52.040 197.770 52.360 197.830 ;
        RECT 55.260 197.970 55.580 198.030 ;
        RECT 56.180 197.970 56.500 198.030 ;
        RECT 55.260 197.830 56.500 197.970 ;
        RECT 55.260 197.770 55.580 197.830 ;
        RECT 56.180 197.770 56.500 197.830 ;
        RECT 69.520 197.970 69.840 198.030 ;
        RECT 71.835 197.970 72.125 198.015 ;
        RECT 69.520 197.830 72.125 197.970 ;
        RECT 69.520 197.770 69.840 197.830 ;
        RECT 71.835 197.785 72.125 197.830 ;
        RECT 73.660 197.970 73.980 198.030 ;
        RECT 77.340 197.970 77.660 198.030 ;
        RECT 73.660 197.830 77.660 197.970 ;
        RECT 73.660 197.770 73.980 197.830 ;
        RECT 77.340 197.770 77.660 197.830 ;
        RECT 79.180 197.970 79.500 198.030 ;
        RECT 80.575 197.970 80.865 198.015 ;
        RECT 79.180 197.830 80.865 197.970 ;
        RECT 79.180 197.770 79.500 197.830 ;
        RECT 80.575 197.785 80.865 197.830 ;
        RECT 84.700 197.970 85.020 198.030 ;
        RECT 85.175 197.970 85.465 198.015 ;
        RECT 84.700 197.830 85.465 197.970 ;
        RECT 84.700 197.770 85.020 197.830 ;
        RECT 85.175 197.785 85.465 197.830 ;
        RECT 88.380 197.970 88.700 198.030 ;
        RECT 89.300 197.970 89.620 198.030 ;
        RECT 88.380 197.830 89.620 197.970 ;
        RECT 88.380 197.770 88.700 197.830 ;
        RECT 89.300 197.770 89.620 197.830 ;
        RECT 91.600 197.970 91.920 198.030 ;
        RECT 95.295 197.970 95.585 198.015 ;
        RECT 91.600 197.830 95.585 197.970 ;
        RECT 91.600 197.770 91.920 197.830 ;
        RECT 95.295 197.785 95.585 197.830 ;
        RECT 96.200 197.970 96.520 198.030 ;
        RECT 99.420 197.970 99.740 198.030 ;
        RECT 96.200 197.830 99.740 197.970 ;
        RECT 96.200 197.770 96.520 197.830 ;
        RECT 99.420 197.770 99.740 197.830 ;
        RECT 104.495 197.970 104.785 198.015 ;
        RECT 104.940 197.970 105.260 198.030 ;
        RECT 120.580 197.970 120.900 198.030 ;
        RECT 123.340 197.970 123.660 198.030 ;
        RECT 135.315 197.970 135.605 198.015 ;
        RECT 135.760 197.970 136.080 198.030 ;
        RECT 104.495 197.830 105.260 197.970 ;
        RECT 104.495 197.785 104.785 197.830 ;
        RECT 104.940 197.770 105.260 197.830 ;
        RECT 105.490 197.830 118.970 197.970 ;
        RECT 28.545 197.630 28.835 197.675 ;
        RECT 30.435 197.630 30.725 197.675 ;
        RECT 33.555 197.630 33.845 197.675 ;
        RECT 28.545 197.490 33.845 197.630 ;
        RECT 28.545 197.445 28.835 197.490 ;
        RECT 30.435 197.445 30.725 197.490 ;
        RECT 33.555 197.445 33.845 197.490 ;
        RECT 30.880 197.290 31.200 197.350 ;
        RECT 12.495 197.150 20.620 197.290 ;
        RECT 12.495 197.105 12.785 197.150 ;
        RECT 20.300 197.090 20.620 197.150 ;
        RECT 23.610 197.150 26.970 197.290 ;
        RECT 27.750 197.150 31.200 197.290 ;
        RECT 6.975 196.950 7.265 196.995 ;
        RECT 13.415 196.950 13.705 196.995 ;
        RECT 14.320 196.950 14.640 197.010 ;
        RECT 17.095 196.950 17.385 196.995 ;
        RECT 6.975 196.810 7.650 196.950 ;
        RECT 6.975 196.765 7.265 196.810 ;
        RECT 7.510 196.315 7.650 196.810 ;
        RECT 13.415 196.810 14.640 196.950 ;
        RECT 13.415 196.765 13.705 196.810 ;
        RECT 14.320 196.750 14.640 196.810 ;
        RECT 15.330 196.810 17.385 196.950 ;
        RECT 9.275 196.610 9.565 196.655 ;
        RECT 14.780 196.610 15.100 196.670 ;
        RECT 9.275 196.470 15.100 196.610 ;
        RECT 9.275 196.425 9.565 196.470 ;
        RECT 14.780 196.410 15.100 196.470 ;
        RECT 7.435 196.085 7.725 196.315 ;
        RECT 9.735 196.270 10.025 196.315 ;
        RECT 12.480 196.270 12.800 196.330 ;
        RECT 15.330 196.315 15.470 196.810 ;
        RECT 17.095 196.765 17.385 196.810 ;
        RECT 20.760 196.950 21.080 197.010 ;
        RECT 23.610 196.995 23.750 197.150 ;
        RECT 21.695 196.950 21.985 196.995 ;
        RECT 20.760 196.810 21.985 196.950 ;
        RECT 20.760 196.750 21.080 196.810 ;
        RECT 21.695 196.765 21.985 196.810 ;
        RECT 23.535 196.765 23.825 196.995 ;
        RECT 25.360 196.750 25.680 197.010 ;
        RECT 25.820 196.950 26.140 197.010 ;
        RECT 27.750 196.995 27.890 197.150 ;
        RECT 30.880 197.090 31.200 197.150 ;
        RECT 37.795 197.290 38.085 197.335 ;
        RECT 38.240 197.290 38.560 197.350 ;
        RECT 37.795 197.150 38.560 197.290 ;
        RECT 37.795 197.105 38.085 197.150 ;
        RECT 38.240 197.090 38.560 197.150 ;
        RECT 27.675 196.950 27.965 196.995 ;
        RECT 25.820 196.810 27.965 196.950 ;
        RECT 25.820 196.750 26.140 196.810 ;
        RECT 27.675 196.765 27.965 196.810 ;
        RECT 28.140 196.950 28.430 196.995 ;
        RECT 29.975 196.950 30.265 196.995 ;
        RECT 33.555 196.950 33.845 196.995 ;
        RECT 28.140 196.810 33.845 196.950 ;
        RECT 28.140 196.765 28.430 196.810 ;
        RECT 29.975 196.765 30.265 196.810 ;
        RECT 33.555 196.765 33.845 196.810 ;
        RECT 34.560 196.970 34.880 197.010 ;
        RECT 34.560 196.750 34.925 196.970 ;
        RECT 39.620 196.950 39.940 197.010 ;
        RECT 19.855 196.610 20.145 196.655 ;
        RECT 18.090 196.470 20.145 196.610 ;
        RECT 18.090 196.330 18.230 196.470 ;
        RECT 19.855 196.425 20.145 196.470 ;
        RECT 22.600 196.410 22.920 196.670 ;
        RECT 34.635 196.655 34.925 196.750 ;
        RECT 35.570 196.810 39.940 196.950 ;
        RECT 23.075 196.425 23.365 196.655 ;
        RECT 31.335 196.610 31.985 196.655 ;
        RECT 34.635 196.610 35.225 196.655 ;
        RECT 31.335 196.470 35.225 196.610 ;
        RECT 31.335 196.425 31.985 196.470 ;
        RECT 34.935 196.425 35.225 196.470 ;
        RECT 12.955 196.270 13.245 196.315 ;
        RECT 9.735 196.130 13.245 196.270 ;
        RECT 9.735 196.085 10.025 196.130 ;
        RECT 12.480 196.070 12.800 196.130 ;
        RECT 12.955 196.085 13.245 196.130 ;
        RECT 15.255 196.085 15.545 196.315 ;
        RECT 17.540 196.070 17.860 196.330 ;
        RECT 18.000 196.070 18.320 196.330 ;
        RECT 19.380 196.070 19.700 196.330 ;
        RECT 20.760 196.270 21.080 196.330 ;
        RECT 23.150 196.270 23.290 196.425 ;
        RECT 20.760 196.130 23.290 196.270 ;
        RECT 28.120 196.270 28.440 196.330 ;
        RECT 35.570 196.270 35.710 196.810 ;
        RECT 39.620 196.750 39.940 196.810 ;
        RECT 38.255 196.610 38.545 196.655 ;
        RECT 38.255 196.470 39.390 196.610 ;
        RECT 38.255 196.425 38.545 196.470 ;
        RECT 39.250 196.330 39.390 196.470 ;
        RECT 28.120 196.130 35.710 196.270 ;
        RECT 36.415 196.270 36.705 196.315 ;
        RECT 38.700 196.270 39.020 196.330 ;
        RECT 36.415 196.130 39.020 196.270 ;
        RECT 20.760 196.070 21.080 196.130 ;
        RECT 28.120 196.070 28.440 196.130 ;
        RECT 36.415 196.085 36.705 196.130 ;
        RECT 38.700 196.070 39.020 196.130 ;
        RECT 39.160 196.070 39.480 196.330 ;
        RECT 41.090 196.270 41.230 197.770 ;
        RECT 49.280 197.630 49.600 197.690 ;
        RECT 46.150 197.490 49.600 197.630 ;
        RECT 46.150 197.335 46.290 197.490 ;
        RECT 49.280 197.430 49.600 197.490 ;
        RECT 51.120 197.430 51.440 197.690 ;
        RECT 58.940 197.630 59.260 197.690 ;
        RECT 62.620 197.630 62.940 197.690 ;
        RECT 103.100 197.630 103.420 197.690 ;
        RECT 105.490 197.630 105.630 197.830 ;
        RECT 118.830 197.690 118.970 197.830 ;
        RECT 120.580 197.830 123.660 197.970 ;
        RECT 120.580 197.770 120.900 197.830 ;
        RECT 123.340 197.770 123.660 197.830 ;
        RECT 127.570 197.830 133.920 197.970 ;
        RECT 127.570 197.690 127.710 197.830 ;
        RECT 56.730 197.490 59.260 197.630 ;
        RECT 46.075 197.105 46.365 197.335 ;
        RECT 48.820 197.290 49.140 197.350 ;
        RECT 47.990 197.150 49.140 197.290 ;
        RECT 51.210 197.290 51.350 197.430 ;
        RECT 52.515 197.290 52.805 197.335 ;
        RECT 53.420 197.290 53.740 197.350 ;
        RECT 51.210 197.150 52.270 197.290 ;
        RECT 41.460 196.950 41.780 197.010 ;
        RECT 41.935 196.950 42.225 196.995 ;
        RECT 41.460 196.810 42.225 196.950 ;
        RECT 41.460 196.750 41.780 196.810 ;
        RECT 41.935 196.765 42.225 196.810 ;
        RECT 45.155 196.950 45.445 196.995 ;
        RECT 45.600 196.950 45.920 197.010 ;
        RECT 45.155 196.810 45.920 196.950 ;
        RECT 45.155 196.765 45.445 196.810 ;
        RECT 45.600 196.750 45.920 196.810 ;
        RECT 46.535 196.765 46.825 196.995 ;
        RECT 42.840 196.610 43.160 196.670 ;
        RECT 43.760 196.610 44.080 196.670 ;
        RECT 42.840 196.470 44.080 196.610 ;
        RECT 46.610 196.610 46.750 196.765 ;
        RECT 46.980 196.750 47.300 197.010 ;
        RECT 47.990 196.995 48.130 197.150 ;
        RECT 48.820 197.090 49.140 197.150 ;
        RECT 47.915 196.765 48.205 196.995 ;
        RECT 49.295 196.765 49.585 196.995 ;
        RECT 49.740 196.950 50.060 197.010 ;
        RECT 50.215 196.950 50.505 196.995 ;
        RECT 49.740 196.810 50.505 196.950 ;
        RECT 48.820 196.610 49.140 196.670 ;
        RECT 46.610 196.470 49.140 196.610 ;
        RECT 49.370 196.610 49.510 196.765 ;
        RECT 49.740 196.750 50.060 196.810 ;
        RECT 50.215 196.765 50.505 196.810 ;
        RECT 50.660 196.750 50.980 197.010 ;
        RECT 51.120 196.750 51.440 197.010 ;
        RECT 51.580 196.750 51.900 197.010 ;
        RECT 52.130 196.995 52.270 197.150 ;
        RECT 52.515 197.150 53.740 197.290 ;
        RECT 52.515 197.105 52.805 197.150 ;
        RECT 53.420 197.090 53.740 197.150 ;
        RECT 54.800 197.290 55.120 197.350 ;
        RECT 56.730 197.290 56.870 197.490 ;
        RECT 58.940 197.430 59.260 197.490 ;
        RECT 60.870 197.490 103.420 197.630 ;
        RECT 54.800 197.150 56.870 197.290 ;
        RECT 54.800 197.090 55.120 197.150 ;
        RECT 56.730 196.995 56.870 197.150 ;
        RECT 52.055 196.765 52.345 196.995 ;
        RECT 55.735 196.950 56.025 196.995 ;
        RECT 53.075 196.810 56.025 196.950 ;
        RECT 51.670 196.610 51.810 196.750 ;
        RECT 53.075 196.610 53.215 196.810 ;
        RECT 55.735 196.765 56.025 196.810 ;
        RECT 56.655 196.765 56.945 196.995 ;
        RECT 57.560 196.950 57.880 197.010 ;
        RECT 58.495 196.950 58.785 196.995 ;
        RECT 58.940 196.950 59.260 197.010 ;
        RECT 60.870 196.995 61.010 197.490 ;
        RECT 62.620 197.430 62.940 197.490 ;
        RECT 103.100 197.430 103.420 197.490 ;
        RECT 104.570 197.490 105.630 197.630 ;
        RECT 68.140 197.290 68.460 197.350 ;
        RECT 69.520 197.290 69.840 197.350 ;
        RECT 72.295 197.290 72.585 197.335 ;
        RECT 81.480 197.290 81.800 197.350 ;
        RECT 65.010 197.150 68.460 197.290 ;
        RECT 57.560 196.810 59.260 196.950 ;
        RECT 57.560 196.750 57.880 196.810 ;
        RECT 58.495 196.765 58.785 196.810 ;
        RECT 58.940 196.750 59.260 196.810 ;
        RECT 60.795 196.765 61.085 196.995 ;
        RECT 62.175 196.950 62.465 196.995 ;
        RECT 62.620 196.950 62.940 197.010 ;
        RECT 62.175 196.810 62.940 196.950 ;
        RECT 62.175 196.765 62.465 196.810 ;
        RECT 62.620 196.750 62.940 196.810 ;
        RECT 63.555 196.950 63.845 196.995 ;
        RECT 65.010 196.950 65.150 197.150 ;
        RECT 68.140 197.090 68.460 197.150 ;
        RECT 69.155 197.150 69.840 197.290 ;
        RECT 63.555 196.810 65.150 196.950 ;
        RECT 63.555 196.765 63.845 196.810 ;
        RECT 65.380 196.750 65.700 197.010 ;
        RECT 65.840 196.950 66.160 197.010 ;
        RECT 69.155 196.995 69.295 197.150 ;
        RECT 69.520 197.090 69.840 197.150 ;
        RECT 70.070 197.150 72.585 197.290 ;
        RECT 70.070 196.995 70.210 197.150 ;
        RECT 72.295 197.105 72.585 197.150 ;
        RECT 77.430 197.150 81.800 197.290 ;
        RECT 68.615 196.950 68.905 196.995 ;
        RECT 65.840 196.810 68.905 196.950 ;
        RECT 65.840 196.750 66.160 196.810 ;
        RECT 68.615 196.765 68.905 196.810 ;
        RECT 69.080 196.765 69.370 196.995 ;
        RECT 69.995 196.765 70.285 196.995 ;
        RECT 71.145 196.950 71.435 196.995 ;
        RECT 72.740 196.950 73.060 197.010 ;
        RECT 71.145 196.810 73.060 196.950 ;
        RECT 71.145 196.765 71.435 196.810 ;
        RECT 72.740 196.750 73.060 196.810 ;
        RECT 73.200 196.750 73.520 197.010 ;
        RECT 74.595 196.950 74.885 196.995 ;
        RECT 75.960 196.950 76.280 197.010 ;
        RECT 74.595 196.810 76.280 196.950 ;
        RECT 74.595 196.765 74.885 196.810 ;
        RECT 75.960 196.750 76.280 196.810 ;
        RECT 76.420 196.750 76.740 197.010 ;
        RECT 77.430 196.995 77.570 197.150 ;
        RECT 81.480 197.090 81.800 197.150 ;
        RECT 87.000 197.290 87.320 197.350 ;
        RECT 93.915 197.330 94.205 197.335 ;
        RECT 93.070 197.290 94.205 197.330 ;
        RECT 87.000 197.190 94.205 197.290 ;
        RECT 87.000 197.150 93.210 197.190 ;
        RECT 87.000 197.090 87.320 197.150 ;
        RECT 93.915 197.105 94.205 197.190 ;
        RECT 98.500 197.290 98.820 197.350 ;
        RECT 101.260 197.290 101.580 197.350 ;
        RECT 98.500 197.150 103.790 197.290 ;
        RECT 98.500 197.090 98.820 197.150 ;
        RECT 101.260 197.090 101.580 197.150 ;
        RECT 77.355 196.765 77.645 196.995 ;
        RECT 78.170 196.950 78.460 196.995 ;
        RECT 77.885 196.810 78.460 196.950 ;
        RECT 49.370 196.470 53.215 196.610 ;
        RECT 42.840 196.410 43.160 196.470 ;
        RECT 43.760 196.410 44.080 196.470 ;
        RECT 48.820 196.410 49.140 196.470 ;
        RECT 53.435 196.425 53.725 196.655 ;
        RECT 53.880 196.610 54.200 196.670 ;
        RECT 54.355 196.610 54.645 196.655 ;
        RECT 53.880 196.470 54.645 196.610 ;
        RECT 53.510 196.270 53.650 196.425 ;
        RECT 53.880 196.410 54.200 196.470 ;
        RECT 54.355 196.425 54.645 196.470 ;
        RECT 54.800 196.410 55.120 196.670 ;
        RECT 59.860 196.410 60.180 196.670 ;
        RECT 64.000 196.410 64.320 196.670 ;
        RECT 64.475 196.610 64.765 196.655 ;
        RECT 70.455 196.610 70.745 196.655 ;
        RECT 75.040 196.610 75.360 196.670 ;
        RECT 64.475 196.470 66.530 196.610 ;
        RECT 64.475 196.425 64.765 196.470 ;
        RECT 55.260 196.270 55.580 196.330 ;
        RECT 41.090 196.130 55.580 196.270 ;
        RECT 55.260 196.070 55.580 196.130 ;
        RECT 57.100 196.270 57.420 196.330 ;
        RECT 57.575 196.270 57.865 196.315 ;
        RECT 57.100 196.130 57.865 196.270 ;
        RECT 57.100 196.070 57.420 196.130 ;
        RECT 57.575 196.085 57.865 196.130 ;
        RECT 58.020 196.270 58.340 196.330 ;
        RECT 60.780 196.270 61.100 196.330 ;
        RECT 58.020 196.130 61.100 196.270 ;
        RECT 58.020 196.070 58.340 196.130 ;
        RECT 60.780 196.070 61.100 196.130 ;
        RECT 61.715 196.270 62.005 196.315 ;
        RECT 62.635 196.270 62.925 196.315 ;
        RECT 61.715 196.130 62.925 196.270 ;
        RECT 61.715 196.085 62.005 196.130 ;
        RECT 62.635 196.085 62.925 196.130 ;
        RECT 63.540 196.270 63.860 196.330 ;
        RECT 65.840 196.270 66.160 196.330 ;
        RECT 63.540 196.130 66.160 196.270 ;
        RECT 66.390 196.270 66.530 196.470 ;
        RECT 70.455 196.470 75.360 196.610 ;
        RECT 76.510 196.610 76.650 196.750 ;
        RECT 77.885 196.610 78.025 196.810 ;
        RECT 78.170 196.765 78.460 196.810 ;
        RECT 78.720 196.950 79.040 197.010 ;
        RECT 79.425 196.950 79.715 196.995 ;
        RECT 81.940 196.950 82.260 197.010 ;
        RECT 78.720 196.810 79.235 196.950 ;
        RECT 79.425 196.810 82.260 196.950 ;
        RECT 78.720 196.750 79.040 196.810 ;
        RECT 79.425 196.765 79.715 196.810 ;
        RECT 81.940 196.750 82.260 196.810 ;
        RECT 85.620 196.950 85.940 197.010 ;
        RECT 86.095 196.950 86.385 196.995 ;
        RECT 85.620 196.810 86.385 196.950 ;
        RECT 85.620 196.750 85.940 196.810 ;
        RECT 86.095 196.765 86.385 196.810 ;
        RECT 86.555 196.950 86.845 196.995 ;
        RECT 86.555 196.810 87.230 196.950 ;
        RECT 86.555 196.765 86.845 196.810 ;
        RECT 87.090 196.670 87.230 196.810 ;
        RECT 87.475 196.765 87.765 196.995 ;
        RECT 76.510 196.470 78.025 196.610 ;
        RECT 82.400 196.610 82.720 196.670 ;
        RECT 82.400 196.470 86.770 196.610 ;
        RECT 70.455 196.425 70.745 196.470 ;
        RECT 75.040 196.410 75.360 196.470 ;
        RECT 82.400 196.410 82.720 196.470 ;
        RECT 67.220 196.270 67.540 196.330 ;
        RECT 74.135 196.270 74.425 196.315 ;
        RECT 86.080 196.270 86.400 196.330 ;
        RECT 66.390 196.130 86.400 196.270 ;
        RECT 86.630 196.270 86.770 196.470 ;
        RECT 87.000 196.410 87.320 196.670 ;
        RECT 87.550 196.270 87.690 196.765 ;
        RECT 89.760 196.750 90.080 197.010 ;
        RECT 90.220 196.750 90.540 197.010 ;
        RECT 91.155 196.950 91.445 196.995 ;
        RECT 91.155 196.810 91.830 196.950 ;
        RECT 93.455 196.815 93.745 197.045 ;
        RECT 94.375 196.950 94.665 196.995 ;
        RECT 91.155 196.765 91.445 196.810 ;
        RECT 89.850 196.610 89.990 196.750 ;
        RECT 89.850 196.470 90.450 196.610 ;
        RECT 89.760 196.270 90.080 196.330 ;
        RECT 90.310 196.315 90.450 196.470 ;
        RECT 86.630 196.130 90.080 196.270 ;
        RECT 63.540 196.070 63.860 196.130 ;
        RECT 65.840 196.070 66.160 196.130 ;
        RECT 67.220 196.070 67.540 196.130 ;
        RECT 74.135 196.085 74.425 196.130 ;
        RECT 86.080 196.070 86.400 196.130 ;
        RECT 89.760 196.070 90.080 196.130 ;
        RECT 90.235 196.085 90.525 196.315 ;
        RECT 91.690 196.270 91.830 196.810 ;
        RECT 93.530 196.670 93.670 196.815 ;
        RECT 93.990 196.810 94.665 196.950 ;
        RECT 93.990 196.670 94.130 196.810 ;
        RECT 94.375 196.765 94.665 196.810 ;
        RECT 95.280 196.950 95.600 197.010 ;
        RECT 95.280 196.810 96.890 196.950 ;
        RECT 95.280 196.750 95.600 196.810 ;
        RECT 93.440 196.410 93.760 196.670 ;
        RECT 93.900 196.410 94.220 196.670 ;
        RECT 96.200 196.655 96.520 196.670 ;
        RECT 96.135 196.425 96.520 196.655 ;
        RECT 96.750 196.610 96.890 196.810 ;
        RECT 102.640 196.750 102.960 197.010 ;
        RECT 103.650 196.995 103.790 197.150 ;
        RECT 103.575 196.765 103.865 196.995 ;
        RECT 104.020 196.750 104.340 197.010 ;
        RECT 97.135 196.610 97.425 196.655 ;
        RECT 102.730 196.610 102.870 196.750 ;
        RECT 96.750 196.470 102.870 196.610 ;
        RECT 97.135 196.425 97.425 196.470 ;
        RECT 96.200 196.410 96.520 196.425 ;
        RECT 92.520 196.270 92.840 196.330 ;
        RECT 104.570 196.270 104.710 197.490 ;
        RECT 111.380 197.430 111.700 197.690 ;
        RECT 111.840 197.630 112.160 197.690 ;
        RECT 117.360 197.630 117.680 197.690 ;
        RECT 111.840 197.490 117.680 197.630 ;
        RECT 111.840 197.430 112.160 197.490 ;
        RECT 117.360 197.430 117.680 197.490 ;
        RECT 118.740 197.430 119.060 197.690 ;
        RECT 121.040 197.630 121.360 197.690 ;
        RECT 126.560 197.630 126.880 197.690 ;
        RECT 121.040 197.490 126.880 197.630 ;
        RECT 121.040 197.430 121.360 197.490 ;
        RECT 126.560 197.430 126.880 197.490 ;
        RECT 127.480 197.430 127.800 197.690 ;
        RECT 133.780 197.630 133.920 197.830 ;
        RECT 135.315 197.830 136.080 197.970 ;
        RECT 135.315 197.785 135.605 197.830 ;
        RECT 135.760 197.770 136.080 197.830 ;
        RECT 138.995 197.970 139.285 198.015 ;
        RECT 139.900 197.970 140.220 198.030 ;
        RECT 138.995 197.830 140.220 197.970 ;
        RECT 138.995 197.785 139.285 197.830 ;
        RECT 139.900 197.770 140.220 197.830 ;
        RECT 153.240 197.970 153.560 198.030 ;
        RECT 153.715 197.970 154.005 198.015 ;
        RECT 153.240 197.830 154.005 197.970 ;
        RECT 153.240 197.770 153.560 197.830 ;
        RECT 153.715 197.785 154.005 197.830 ;
        RECT 141.280 197.630 141.600 197.690 ;
        RECT 145.880 197.630 146.200 197.690 ;
        RECT 154.160 197.630 154.480 197.690 ;
        RECT 133.780 197.490 146.200 197.630 ;
        RECT 141.280 197.430 141.600 197.490 ;
        RECT 145.880 197.430 146.200 197.490 ;
        RECT 151.950 197.490 154.480 197.630 ;
        RECT 104.955 197.290 105.245 197.335 ;
        RECT 117.820 197.290 118.140 197.350 ;
        RECT 104.955 197.150 107.930 197.290 ;
        RECT 104.955 197.105 105.245 197.150 ;
        RECT 105.400 196.410 105.720 196.670 ;
        RECT 106.320 196.410 106.640 196.670 ;
        RECT 107.790 196.610 107.930 197.150 ;
        RECT 110.550 197.150 118.140 197.290 ;
        RECT 108.175 196.950 108.465 196.995 ;
        RECT 110.000 196.950 110.320 197.010 ;
        RECT 110.550 196.995 110.690 197.150 ;
        RECT 117.820 197.090 118.140 197.150 ;
        RECT 119.660 197.290 119.980 197.350 ;
        RECT 131.160 197.290 131.480 197.350 ;
        RECT 133.000 197.290 133.320 197.350 ;
        RECT 134.840 197.290 135.160 197.350 ;
        RECT 135.905 197.290 136.910 197.330 ;
        RECT 143.120 197.290 143.440 197.350 ;
        RECT 119.660 197.150 133.690 197.290 ;
        RECT 119.660 197.090 119.980 197.150 ;
        RECT 131.160 197.090 131.480 197.150 ;
        RECT 133.000 197.090 133.320 197.150 ;
        RECT 108.175 196.810 110.320 196.950 ;
        RECT 108.175 196.765 108.465 196.810 ;
        RECT 110.000 196.750 110.320 196.810 ;
        RECT 110.475 196.765 110.765 196.995 ;
        RECT 110.935 196.950 111.225 196.995 ;
        RECT 111.380 196.950 111.700 197.010 ;
        RECT 110.935 196.810 111.700 196.950 ;
        RECT 110.935 196.765 111.225 196.810 ;
        RECT 111.380 196.750 111.700 196.810 ;
        RECT 111.855 196.765 112.145 196.995 ;
        RECT 111.930 196.610 112.070 196.765 ;
        RECT 114.600 196.750 114.920 197.010 ;
        RECT 133.550 196.995 133.690 197.150 ;
        RECT 134.840 197.190 139.670 197.290 ;
        RECT 134.840 197.150 136.045 197.190 ;
        RECT 136.770 197.150 139.670 197.190 ;
        RECT 134.840 197.090 135.160 197.150 ;
        RECT 132.100 196.950 132.390 196.995 ;
        RECT 115.150 196.810 132.390 196.950 ;
        RECT 114.690 196.610 114.830 196.750 ;
        RECT 107.790 196.470 109.770 196.610 ;
        RECT 111.930 196.470 114.830 196.610 ;
        RECT 91.690 196.130 104.710 196.270 ;
        RECT 92.520 196.070 92.840 196.130 ;
        RECT 106.780 196.070 107.100 196.330 ;
        RECT 107.255 196.270 107.545 196.315 ;
        RECT 108.160 196.270 108.480 196.330 ;
        RECT 109.630 196.315 109.770 196.470 ;
        RECT 107.255 196.130 108.480 196.270 ;
        RECT 107.255 196.085 107.545 196.130 ;
        RECT 108.160 196.070 108.480 196.130 ;
        RECT 109.555 196.270 109.845 196.315 ;
        RECT 115.150 196.270 115.290 196.810 ;
        RECT 132.100 196.765 132.390 196.810 ;
        RECT 132.555 196.765 132.845 196.995 ;
        RECT 133.475 196.765 133.765 196.995 ;
        RECT 134.380 196.950 134.700 197.010 ;
        RECT 135.300 196.950 135.620 197.010 ;
        RECT 134.380 196.810 135.620 196.950 ;
        RECT 136.235 196.815 136.525 197.045 ;
        RECT 118.740 196.610 119.060 196.670 ;
        RECT 125.655 196.610 125.945 196.655 ;
        RECT 132.630 196.610 132.770 196.765 ;
        RECT 134.380 196.750 134.700 196.810 ;
        RECT 135.300 196.750 135.620 196.810 ;
        RECT 136.310 196.670 136.450 196.815 ;
        RECT 136.695 196.765 136.985 196.995 ;
        RECT 137.140 196.950 137.460 197.010 ;
        RECT 137.615 196.950 137.905 196.995 ;
        RECT 137.140 196.810 137.905 196.950 ;
        RECT 118.740 196.470 132.770 196.610 ;
        RECT 133.935 196.610 134.225 196.655 ;
        RECT 134.840 196.610 135.160 196.670 ;
        RECT 135.760 196.610 136.080 196.670 ;
        RECT 133.935 196.470 136.080 196.610 ;
        RECT 118.740 196.410 119.060 196.470 ;
        RECT 125.655 196.425 125.945 196.470 ;
        RECT 132.170 196.330 132.310 196.470 ;
        RECT 133.935 196.425 134.225 196.470 ;
        RECT 134.840 196.410 135.160 196.470 ;
        RECT 135.760 196.410 136.080 196.470 ;
        RECT 136.220 196.410 136.540 196.670 ;
        RECT 136.770 196.610 136.910 196.765 ;
        RECT 137.140 196.750 137.460 196.810 ;
        RECT 137.615 196.765 137.905 196.810 ;
        RECT 138.060 196.750 138.380 197.010 ;
        RECT 139.530 196.995 139.670 197.150 ;
        RECT 140.450 197.150 143.440 197.290 ;
        RECT 140.450 196.995 140.590 197.150 ;
        RECT 143.120 197.090 143.440 197.150 ;
        RECT 144.500 197.290 144.820 197.350 ;
        RECT 145.420 197.290 145.740 197.350 ;
        RECT 144.500 197.150 145.740 197.290 ;
        RECT 144.500 197.090 144.820 197.150 ;
        RECT 145.420 197.090 145.740 197.150 ;
        RECT 139.455 196.765 139.745 196.995 ;
        RECT 140.375 196.765 140.665 196.995 ;
        RECT 146.800 196.950 147.120 197.010 ;
        RECT 150.495 196.950 150.785 196.995 ;
        RECT 146.800 196.810 150.785 196.950 ;
        RECT 146.800 196.750 147.120 196.810 ;
        RECT 150.495 196.765 150.785 196.810 ;
        RECT 150.960 196.950 151.250 196.995 ;
        RECT 151.950 196.950 152.090 197.490 ;
        RECT 154.160 197.430 154.480 197.490 ;
        RECT 152.320 197.090 152.640 197.350 ;
        RECT 150.960 196.810 152.090 196.950 ;
        RECT 152.410 196.950 152.550 197.090 ;
        RECT 152.820 196.950 153.110 196.995 ;
        RECT 152.410 196.810 153.110 196.950 ;
        RECT 150.960 196.765 151.250 196.810 ;
        RECT 152.820 196.765 153.110 196.810 ;
        RECT 139.915 196.610 140.205 196.655 ;
        RECT 136.770 196.470 140.205 196.610 ;
        RECT 139.915 196.425 140.205 196.470 ;
        RECT 141.740 196.610 142.060 196.670 ;
        RECT 151.030 196.610 151.170 196.765 ;
        RECT 141.740 196.470 151.170 196.610 ;
        RECT 141.740 196.410 142.060 196.470 ;
        RECT 151.860 196.410 152.180 196.670 ;
        RECT 152.335 196.425 152.625 196.655 ;
        RECT 109.555 196.130 115.290 196.270 ;
        RECT 115.520 196.270 115.840 196.330 ;
        RECT 126.560 196.270 126.880 196.330 ;
        RECT 115.520 196.130 126.880 196.270 ;
        RECT 109.555 196.085 109.845 196.130 ;
        RECT 115.520 196.070 115.840 196.130 ;
        RECT 126.560 196.070 126.880 196.130 ;
        RECT 132.080 196.070 132.400 196.330 ;
        RECT 135.300 196.270 135.620 196.330 ;
        RECT 150.940 196.270 151.260 196.330 ;
        RECT 135.300 196.130 151.260 196.270 ;
        RECT 152.410 196.270 152.550 196.425 ;
        RECT 152.780 196.270 153.100 196.330 ;
        RECT 152.410 196.130 153.100 196.270 ;
        RECT 135.300 196.070 135.620 196.130 ;
        RECT 150.940 196.070 151.260 196.130 ;
        RECT 152.780 196.070 153.100 196.130 ;
        RECT 2.750 195.450 159.030 195.930 ;
        RECT 18.460 195.250 18.780 195.310 ;
        RECT 25.820 195.250 26.140 195.310 ;
        RECT 38.255 195.250 38.545 195.295 ;
        RECT 4.290 195.110 26.140 195.250 ;
        RECT 4.290 194.615 4.430 195.110 ;
        RECT 7.875 194.910 8.525 194.955 ;
        RECT 11.475 194.910 11.765 194.955 ;
        RECT 7.875 194.770 11.765 194.910 ;
        RECT 7.875 194.725 8.525 194.770 ;
        RECT 11.175 194.725 11.765 194.770 ;
        RECT 4.215 194.385 4.505 194.615 ;
        RECT 4.680 194.570 4.970 194.615 ;
        RECT 6.515 194.570 6.805 194.615 ;
        RECT 10.095 194.570 10.385 194.615 ;
        RECT 4.680 194.430 10.385 194.570 ;
        RECT 4.680 194.385 4.970 194.430 ;
        RECT 6.515 194.385 6.805 194.430 ;
        RECT 10.095 194.385 10.385 194.430 ;
        RECT 11.175 194.570 11.465 194.725 ;
        RECT 13.860 194.570 14.180 194.630 ;
        RECT 15.330 194.615 15.470 195.110 ;
        RECT 18.460 195.050 18.780 195.110 ;
        RECT 25.820 195.050 26.140 195.110 ;
        RECT 29.065 195.110 38.545 195.250 ;
        RECT 18.915 194.910 19.565 194.955 ;
        RECT 22.515 194.910 22.805 194.955 ;
        RECT 18.915 194.770 22.805 194.910 ;
        RECT 18.915 194.725 19.565 194.770 ;
        RECT 22.215 194.725 22.805 194.770 ;
        RECT 11.175 194.430 14.180 194.570 ;
        RECT 11.175 194.410 11.465 194.430 ;
        RECT 13.860 194.370 14.180 194.430 ;
        RECT 15.255 194.385 15.545 194.615 ;
        RECT 15.720 194.570 16.010 194.615 ;
        RECT 17.555 194.570 17.845 194.615 ;
        RECT 21.135 194.570 21.425 194.615 ;
        RECT 15.720 194.430 21.425 194.570 ;
        RECT 15.720 194.385 16.010 194.430 ;
        RECT 17.555 194.385 17.845 194.430 ;
        RECT 21.135 194.385 21.425 194.430 ;
        RECT 22.215 194.570 22.505 194.725 ;
        RECT 23.520 194.570 23.840 194.630 ;
        RECT 24.455 194.570 24.745 194.615 ;
        RECT 22.215 194.430 24.745 194.570 ;
        RECT 25.910 194.570 26.050 195.050 ;
        RECT 26.295 194.910 26.585 194.955 ;
        RECT 28.120 194.910 28.440 194.970 ;
        RECT 26.295 194.770 28.440 194.910 ;
        RECT 26.295 194.725 26.585 194.770 ;
        RECT 28.120 194.710 28.440 194.770 ;
        RECT 27.215 194.570 27.505 194.615 ;
        RECT 29.065 194.570 29.205 195.110 ;
        RECT 38.255 195.065 38.545 195.110 ;
        RECT 38.700 195.250 39.020 195.310 ;
        RECT 42.840 195.250 43.160 195.310 ;
        RECT 47.900 195.250 48.220 195.310 ;
        RECT 38.700 195.110 48.220 195.250 ;
        RECT 38.700 195.050 39.020 195.110 ;
        RECT 42.840 195.050 43.160 195.110 ;
        RECT 47.900 195.050 48.220 195.110 ;
        RECT 48.820 195.250 49.140 195.310 ;
        RECT 50.200 195.250 50.520 195.310 ;
        RECT 48.820 195.110 50.520 195.250 ;
        RECT 48.820 195.050 49.140 195.110 ;
        RECT 50.200 195.050 50.520 195.110 ;
        RECT 50.675 195.065 50.965 195.295 ;
        RECT 32.715 194.910 33.365 194.955 ;
        RECT 36.315 194.910 36.605 194.955 ;
        RECT 36.860 194.910 37.180 194.970 ;
        RECT 50.750 194.910 50.890 195.065 ;
        RECT 52.960 195.050 53.280 195.310 ;
        RECT 65.380 195.250 65.700 195.310 ;
        RECT 71.835 195.250 72.125 195.295 ;
        RECT 59.030 195.110 65.150 195.250 ;
        RECT 32.715 194.770 46.750 194.910 ;
        RECT 32.715 194.725 33.365 194.770 ;
        RECT 36.015 194.725 36.605 194.770 ;
        RECT 25.910 194.430 26.970 194.570 ;
        RECT 22.215 194.410 22.505 194.430 ;
        RECT 23.520 194.370 23.840 194.430 ;
        RECT 24.455 194.385 24.745 194.430 ;
        RECT 5.580 194.030 5.900 194.290 ;
        RECT 16.635 194.230 16.925 194.275 ;
        RECT 17.080 194.230 17.400 194.290 ;
        RECT 16.635 194.090 17.400 194.230 ;
        RECT 16.635 194.045 16.925 194.090 ;
        RECT 17.080 194.030 17.400 194.090 ;
        RECT 18.920 194.230 19.240 194.290 ;
        RECT 26.830 194.230 26.970 194.430 ;
        RECT 27.215 194.560 28.350 194.570 ;
        RECT 28.670 194.560 29.205 194.570 ;
        RECT 27.215 194.430 29.205 194.560 ;
        RECT 29.520 194.570 29.810 194.615 ;
        RECT 31.355 194.570 31.645 194.615 ;
        RECT 34.935 194.570 35.225 194.615 ;
        RECT 29.520 194.430 35.225 194.570 ;
        RECT 27.215 194.385 27.505 194.430 ;
        RECT 28.210 194.420 28.810 194.430 ;
        RECT 29.520 194.385 29.810 194.430 ;
        RECT 31.355 194.385 31.645 194.430 ;
        RECT 34.935 194.385 35.225 194.430 ;
        RECT 36.015 194.410 36.305 194.725 ;
        RECT 36.860 194.710 37.180 194.770 ;
        RECT 39.160 194.570 39.480 194.630 ;
        RECT 40.095 194.570 40.385 194.615 ;
        RECT 37.870 194.430 40.385 194.570 ;
        RECT 29.055 194.230 29.345 194.275 ;
        RECT 30.435 194.230 30.725 194.275 ;
        RECT 18.920 194.090 26.510 194.230 ;
        RECT 26.830 194.090 29.345 194.230 ;
        RECT 18.920 194.030 19.240 194.090 ;
        RECT 26.370 193.950 26.510 194.090 ;
        RECT 29.055 194.045 29.345 194.090 ;
        RECT 29.590 194.090 30.725 194.230 ;
        RECT 5.085 193.890 5.375 193.935 ;
        RECT 6.975 193.890 7.265 193.935 ;
        RECT 10.095 193.890 10.385 193.935 ;
        RECT 5.085 193.750 10.385 193.890 ;
        RECT 5.085 193.705 5.375 193.750 ;
        RECT 6.975 193.705 7.265 193.750 ;
        RECT 10.095 193.705 10.385 193.750 ;
        RECT 16.125 193.890 16.415 193.935 ;
        RECT 18.015 193.890 18.305 193.935 ;
        RECT 21.135 193.890 21.425 193.935 ;
        RECT 16.125 193.750 21.425 193.890 ;
        RECT 16.125 193.705 16.415 193.750 ;
        RECT 18.015 193.705 18.305 193.750 ;
        RECT 21.135 193.705 21.425 193.750 ;
        RECT 26.280 193.690 26.600 193.950 ;
        RECT 28.135 193.890 28.425 193.935 ;
        RECT 29.590 193.890 29.730 194.090 ;
        RECT 30.435 194.045 30.725 194.090 ;
        RECT 35.480 194.030 35.800 194.290 ;
        RECT 37.870 194.275 38.010 194.430 ;
        RECT 39.160 194.370 39.480 194.430 ;
        RECT 40.095 194.385 40.385 194.430 ;
        RECT 40.555 194.570 40.845 194.615 ;
        RECT 40.555 194.430 41.690 194.570 ;
        RECT 40.555 194.385 40.845 194.430 ;
        RECT 37.795 194.045 38.085 194.275 ;
        RECT 41.015 194.045 41.305 194.275 ;
        RECT 28.135 193.750 29.730 193.890 ;
        RECT 29.925 193.890 30.215 193.935 ;
        RECT 31.815 193.890 32.105 193.935 ;
        RECT 34.935 193.890 35.225 193.935 ;
        RECT 29.925 193.750 35.225 193.890 ;
        RECT 35.570 193.890 35.710 194.030 ;
        RECT 41.090 193.890 41.230 194.045 ;
        RECT 35.570 193.750 41.230 193.890 ;
        RECT 41.550 193.890 41.690 194.430 ;
        RECT 46.610 194.290 46.750 194.770 ;
        RECT 50.290 194.770 50.890 194.910 ;
        RECT 53.050 194.910 53.190 195.050 ;
        RECT 57.100 194.910 57.420 194.970 ;
        RECT 53.050 194.770 57.420 194.910 ;
        RECT 47.455 194.385 47.745 194.615 ;
        RECT 49.295 194.580 49.585 194.615 ;
        RECT 49.740 194.580 50.060 194.630 ;
        RECT 50.290 194.615 50.430 194.770 ;
        RECT 51.580 194.615 51.900 194.630 ;
        RECT 49.295 194.440 50.060 194.580 ;
        RECT 49.295 194.385 49.585 194.440 ;
        RECT 42.855 194.230 43.145 194.275 ;
        RECT 43.760 194.230 44.080 194.290 ;
        RECT 42.855 194.090 44.080 194.230 ;
        RECT 42.855 194.045 43.145 194.090 ;
        RECT 43.760 194.030 44.080 194.090 ;
        RECT 44.680 194.030 45.000 194.290 ;
        RECT 46.520 194.030 46.840 194.290 ;
        RECT 44.770 193.890 44.910 194.030 ;
        RECT 41.550 193.750 44.910 193.890 ;
        RECT 28.135 193.705 28.425 193.750 ;
        RECT 29.925 193.705 30.215 193.750 ;
        RECT 31.815 193.705 32.105 193.750 ;
        RECT 34.935 193.705 35.225 193.750 ;
        RECT 12.940 193.550 13.260 193.610 ;
        RECT 18.920 193.550 19.240 193.610 ;
        RECT 12.940 193.410 19.240 193.550 ;
        RECT 12.940 193.350 13.260 193.410 ;
        RECT 18.920 193.350 19.240 193.410 ;
        RECT 19.380 193.550 19.700 193.610 ;
        RECT 23.980 193.550 24.300 193.610 ;
        RECT 19.380 193.410 24.300 193.550 ;
        RECT 19.380 193.350 19.700 193.410 ;
        RECT 23.980 193.350 24.300 193.410 ;
        RECT 25.820 193.550 26.140 193.610 ;
        RECT 26.740 193.550 27.060 193.610 ;
        RECT 25.820 193.410 27.060 193.550 ;
        RECT 25.820 193.350 26.140 193.410 ;
        RECT 26.740 193.350 27.060 193.410 ;
        RECT 45.600 193.350 45.920 193.610 ;
        RECT 46.535 193.550 46.825 193.595 ;
        RECT 46.980 193.550 47.300 193.610 ;
        RECT 46.535 193.410 47.300 193.550 ;
        RECT 47.530 193.550 47.670 194.385 ;
        RECT 49.740 194.370 50.060 194.440 ;
        RECT 50.215 194.385 50.505 194.615 ;
        RECT 51.570 194.570 51.900 194.615 ;
        RECT 51.385 194.430 51.900 194.570 ;
        RECT 51.570 194.385 51.900 194.430 ;
        RECT 51.580 194.370 51.900 194.385 ;
        RECT 52.040 194.370 52.360 194.630 ;
        RECT 52.500 194.370 52.820 194.630 ;
        RECT 52.960 194.615 53.280 194.630 ;
        RECT 53.970 194.615 54.110 194.770 ;
        RECT 57.100 194.710 57.420 194.770 ;
        RECT 52.960 194.385 53.445 194.615 ;
        RECT 53.895 194.385 54.185 194.615 ;
        RECT 54.815 194.385 55.105 194.615 ;
        RECT 55.260 194.570 55.580 194.630 ;
        RECT 59.030 194.615 59.170 195.110 ;
        RECT 59.400 194.710 59.720 194.970 ;
        RECT 60.780 194.910 61.100 194.970 ;
        RECT 65.010 194.910 65.150 195.110 ;
        RECT 65.380 195.110 72.125 195.250 ;
        RECT 65.380 195.050 65.700 195.110 ;
        RECT 71.835 195.065 72.125 195.110 ;
        RECT 72.280 195.250 72.600 195.310 ;
        RECT 77.800 195.250 78.120 195.310 ;
        RECT 92.060 195.250 92.380 195.310 ;
        RECT 72.280 195.110 92.380 195.250 ;
        RECT 72.280 195.050 72.600 195.110 ;
        RECT 77.800 195.050 78.120 195.110 ;
        RECT 69.520 194.910 69.840 194.970 ;
        RECT 60.780 194.770 61.930 194.910 ;
        RECT 65.010 194.770 71.130 194.910 ;
        RECT 60.780 194.710 61.100 194.770 ;
        RECT 57.575 194.570 57.865 194.615 ;
        RECT 55.260 194.430 57.865 194.570 ;
        RECT 52.960 194.370 53.280 194.385 ;
        RECT 48.360 194.030 48.680 194.290 ;
        RECT 48.820 194.030 49.140 194.290 ;
        RECT 54.890 194.230 55.030 194.385 ;
        RECT 55.260 194.370 55.580 194.430 ;
        RECT 57.575 194.385 57.865 194.430 ;
        RECT 58.495 194.385 58.785 194.615 ;
        RECT 58.955 194.385 59.245 194.615 ;
        RECT 49.830 194.090 55.030 194.230 ;
        RECT 58.570 194.230 58.710 194.385 ;
        RECT 59.490 194.230 59.630 194.710 ;
        RECT 59.875 194.385 60.165 194.615 ;
        RECT 58.570 194.090 59.630 194.230 ;
        RECT 59.950 194.230 60.090 194.385 ;
        RECT 60.320 194.370 60.640 194.630 ;
        RECT 61.790 194.615 61.930 194.770 ;
        RECT 69.520 194.710 69.840 194.770 ;
        RECT 61.715 194.385 62.005 194.615 ;
        RECT 62.635 194.570 62.925 194.615 ;
        RECT 66.760 194.570 67.080 194.630 ;
        RECT 62.635 194.430 67.080 194.570 ;
        RECT 62.635 194.385 62.925 194.430 ;
        RECT 66.760 194.370 67.080 194.430 ;
        RECT 70.455 194.385 70.745 194.615 ;
        RECT 63.080 194.230 63.400 194.290 ;
        RECT 59.950 194.090 63.400 194.230 ;
        RECT 49.830 193.890 49.970 194.090 ;
        RECT 63.080 194.030 63.400 194.090 ;
        RECT 63.540 194.030 63.860 194.290 ;
        RECT 64.475 194.045 64.765 194.275 ;
        RECT 64.935 194.045 65.225 194.275 ;
        RECT 48.935 193.750 49.970 193.890 ;
        RECT 51.120 193.890 51.440 193.950 ;
        RECT 54.800 193.890 55.120 193.950 ;
        RECT 51.120 193.750 55.120 193.890 ;
        RECT 48.935 193.550 49.075 193.750 ;
        RECT 51.120 193.690 51.440 193.750 ;
        RECT 54.800 193.690 55.120 193.750 ;
        RECT 62.175 193.890 62.465 193.935 ;
        RECT 64.550 193.890 64.690 194.045 ;
        RECT 62.175 193.750 64.690 193.890 ;
        RECT 65.010 193.890 65.150 194.045 ;
        RECT 65.380 194.030 65.700 194.290 ;
        RECT 65.855 194.230 66.145 194.275 ;
        RECT 65.855 194.090 66.990 194.230 ;
        RECT 65.855 194.045 66.145 194.090 ;
        RECT 66.850 193.950 66.990 194.090 ;
        RECT 65.010 193.750 66.530 193.890 ;
        RECT 62.175 193.705 62.465 193.750 ;
        RECT 47.530 193.410 49.075 193.550 ;
        RECT 61.255 193.550 61.545 193.595 ;
        RECT 65.840 193.550 66.160 193.610 ;
        RECT 61.255 193.410 66.160 193.550 ;
        RECT 66.390 193.550 66.530 193.750 ;
        RECT 66.760 193.690 67.080 193.950 ;
        RECT 70.530 193.890 70.670 194.385 ;
        RECT 70.990 194.230 71.130 194.770 ;
        RECT 71.450 194.770 73.890 194.910 ;
        RECT 71.450 194.615 71.590 194.770 ;
        RECT 73.750 194.630 73.890 194.770 ;
        RECT 71.375 194.385 71.665 194.615 ;
        RECT 71.820 194.570 72.140 194.630 ;
        RECT 72.755 194.570 73.045 194.615 ;
        RECT 73.200 194.570 73.520 194.630 ;
        RECT 71.820 194.430 73.520 194.570 ;
        RECT 71.820 194.370 72.140 194.430 ;
        RECT 72.755 194.385 73.045 194.430 ;
        RECT 73.200 194.370 73.520 194.430 ;
        RECT 73.660 194.370 73.980 194.630 ;
        RECT 74.135 194.570 74.425 194.615 ;
        RECT 74.580 194.570 74.900 194.630 ;
        RECT 81.570 194.615 81.710 195.110 ;
        RECT 92.060 195.050 92.380 195.110 ;
        RECT 98.515 195.250 98.805 195.295 ;
        RECT 100.815 195.250 101.105 195.295 ;
        RECT 98.515 195.110 101.105 195.250 ;
        RECT 98.515 195.065 98.805 195.110 ;
        RECT 100.815 195.065 101.105 195.110 ;
        RECT 103.100 195.250 103.420 195.310 ;
        RECT 106.320 195.250 106.640 195.310 ;
        RECT 103.100 195.110 106.640 195.250 ;
        RECT 103.100 195.050 103.420 195.110 ;
        RECT 106.320 195.050 106.640 195.110 ;
        RECT 108.160 195.250 108.480 195.310 ;
        RECT 123.340 195.250 123.660 195.310 ;
        RECT 126.575 195.250 126.865 195.295 ;
        RECT 108.160 195.110 123.110 195.250 ;
        RECT 108.160 195.050 108.480 195.110 ;
        RECT 82.860 194.710 83.180 194.970 ;
        RECT 89.300 194.910 89.620 194.970 ;
        RECT 111.380 194.910 111.700 194.970 ;
        RECT 111.855 194.910 112.145 194.955 ;
        RECT 83.410 194.770 88.150 194.910 ;
        RECT 74.135 194.430 74.900 194.570 ;
        RECT 74.135 194.385 74.425 194.430 ;
        RECT 74.580 194.370 74.900 194.430 ;
        RECT 81.495 194.385 81.785 194.615 ;
        RECT 81.940 194.570 82.260 194.630 ;
        RECT 83.410 194.570 83.550 194.770 ;
        RECT 84.790 194.615 84.930 194.770 ;
        RECT 81.940 194.430 83.550 194.570 ;
        RECT 81.940 194.370 82.260 194.430 ;
        RECT 83.795 194.385 84.085 194.615 ;
        RECT 84.715 194.385 85.005 194.615 ;
        RECT 80.575 194.230 80.865 194.275 ;
        RECT 82.030 194.230 82.170 194.370 ;
        RECT 70.990 194.090 74.810 194.230 ;
        RECT 74.670 193.950 74.810 194.090 ;
        RECT 80.575 194.090 82.170 194.230 ;
        RECT 80.575 194.045 80.865 194.090 ;
        RECT 83.320 194.030 83.640 194.290 ;
        RECT 83.870 194.230 84.010 194.385 ;
        RECT 86.080 194.370 86.400 194.630 ;
        RECT 87.015 194.570 87.305 194.615 ;
        RECT 87.460 194.570 87.780 194.630 ;
        RECT 87.015 194.430 87.780 194.570 ;
        RECT 88.010 194.570 88.150 194.770 ;
        RECT 89.300 194.770 110.230 194.910 ;
        RECT 89.300 194.710 89.620 194.770 ;
        RECT 97.595 194.570 97.885 194.615 ;
        RECT 98.500 194.570 98.820 194.630 ;
        RECT 88.010 194.430 97.350 194.570 ;
        RECT 87.015 194.385 87.305 194.430 ;
        RECT 87.460 194.370 87.780 194.430 ;
        RECT 84.240 194.230 84.560 194.290 ;
        RECT 92.980 194.230 93.300 194.290 ;
        RECT 83.870 194.090 84.560 194.230 ;
        RECT 72.280 193.890 72.600 193.950 ;
        RECT 70.530 193.750 72.600 193.890 ;
        RECT 72.280 193.690 72.600 193.750 ;
        RECT 73.215 193.705 73.505 193.935 ;
        RECT 70.440 193.550 70.760 193.610 ;
        RECT 66.390 193.410 70.760 193.550 ;
        RECT 46.535 193.365 46.825 193.410 ;
        RECT 46.980 193.350 47.300 193.410 ;
        RECT 61.255 193.365 61.545 193.410 ;
        RECT 65.840 193.350 66.160 193.410 ;
        RECT 70.440 193.350 70.760 193.410 ;
        RECT 71.375 193.550 71.665 193.595 ;
        RECT 71.820 193.550 72.140 193.610 ;
        RECT 71.375 193.410 72.140 193.550 ;
        RECT 73.290 193.550 73.430 193.705 ;
        RECT 73.660 193.690 73.980 193.950 ;
        RECT 74.580 193.690 74.900 193.950 ;
        RECT 81.480 193.890 81.800 193.950 ;
        RECT 83.870 193.890 84.010 194.090 ;
        RECT 84.240 194.030 84.560 194.090 ;
        RECT 87.090 194.090 93.300 194.230 ;
        RECT 97.210 194.230 97.350 194.430 ;
        RECT 97.595 194.430 98.820 194.570 ;
        RECT 97.595 194.385 97.885 194.430 ;
        RECT 98.500 194.370 98.820 194.430 ;
        RECT 98.975 194.385 99.265 194.615 ;
        RECT 97.210 194.090 98.730 194.230 ;
        RECT 87.090 193.890 87.230 194.090 ;
        RECT 92.980 194.030 93.300 194.090 ;
        RECT 98.590 193.950 98.730 194.090 ;
        RECT 81.480 193.750 87.230 193.890 ;
        RECT 90.220 193.890 90.540 193.950 ;
        RECT 95.740 193.890 96.060 193.950 ;
        RECT 90.220 193.750 96.060 193.890 ;
        RECT 81.480 193.690 81.800 193.750 ;
        RECT 90.220 193.690 90.540 193.750 ;
        RECT 95.740 193.690 96.060 193.750 ;
        RECT 96.675 193.890 96.965 193.935 ;
        RECT 97.120 193.890 97.440 193.950 ;
        RECT 96.675 193.750 97.440 193.890 ;
        RECT 96.675 193.705 96.965 193.750 ;
        RECT 97.120 193.690 97.440 193.750 ;
        RECT 98.500 193.690 98.820 193.950 ;
        RECT 99.100 193.890 99.240 194.385 ;
        RECT 99.420 194.370 99.740 194.630 ;
        RECT 100.430 194.615 100.570 194.770 ;
        RECT 100.355 194.385 100.645 194.615 ;
        RECT 100.800 194.370 101.120 194.630 ;
        RECT 101.735 194.570 102.025 194.615 ;
        RECT 102.640 194.570 102.960 194.630 ;
        RECT 101.735 194.430 102.960 194.570 ;
        RECT 101.735 194.385 102.025 194.430 ;
        RECT 102.640 194.370 102.960 194.430 ;
        RECT 104.480 194.570 104.800 194.630 ;
        RECT 107.700 194.570 108.020 194.630 ;
        RECT 110.090 194.615 110.230 194.770 ;
        RECT 111.380 194.770 112.145 194.910 ;
        RECT 111.380 194.710 111.700 194.770 ;
        RECT 111.855 194.725 112.145 194.770 ;
        RECT 113.680 194.910 114.000 194.970 ;
        RECT 121.040 194.910 121.360 194.970 ;
        RECT 113.680 194.770 117.130 194.910 ;
        RECT 113.680 194.710 114.000 194.770 ;
        RECT 104.480 194.430 108.020 194.570 ;
        RECT 104.480 194.370 104.800 194.430 ;
        RECT 107.700 194.370 108.020 194.430 ;
        RECT 110.015 194.385 110.305 194.615 ;
        RECT 112.760 194.570 113.080 194.630 ;
        RECT 115.075 194.570 115.365 194.615 ;
        RECT 112.760 194.430 115.365 194.570 ;
        RECT 112.760 194.370 113.080 194.430 ;
        RECT 115.075 194.385 115.365 194.430 ;
        RECT 115.520 194.370 115.840 194.630 ;
        RECT 115.995 194.570 116.285 194.615 ;
        RECT 116.440 194.570 116.760 194.630 ;
        RECT 116.990 194.615 117.130 194.770 ;
        RECT 117.450 194.770 121.360 194.910 ;
        RECT 117.450 194.615 117.590 194.770 ;
        RECT 121.040 194.710 121.360 194.770 ;
        RECT 121.500 194.710 121.820 194.970 ;
        RECT 121.960 194.710 122.280 194.970 ;
        RECT 115.995 194.430 116.760 194.570 ;
        RECT 115.995 194.385 116.285 194.430 ;
        RECT 116.440 194.370 116.760 194.430 ;
        RECT 116.915 194.385 117.205 194.615 ;
        RECT 117.375 194.385 117.665 194.615 ;
        RECT 121.590 194.565 121.730 194.710 ;
        RECT 121.515 194.335 121.805 194.565 ;
        RECT 122.435 194.385 122.725 194.615 ;
        RECT 122.970 194.570 123.110 195.110 ;
        RECT 123.340 195.110 126.865 195.250 ;
        RECT 123.340 195.050 123.660 195.110 ;
        RECT 126.575 195.065 126.865 195.110 ;
        RECT 128.860 195.250 129.180 195.310 ;
        RECT 132.095 195.250 132.385 195.295 ;
        RECT 128.860 195.110 132.385 195.250 ;
        RECT 128.860 195.050 129.180 195.110 ;
        RECT 132.095 195.065 132.385 195.110 ;
        RECT 133.000 195.250 133.320 195.310 ;
        RECT 134.840 195.250 135.160 195.310 ;
        RECT 133.000 195.110 135.160 195.250 ;
        RECT 133.000 195.050 133.320 195.110 ;
        RECT 134.840 195.050 135.160 195.110 ;
        RECT 135.760 195.050 136.080 195.310 ;
        RECT 137.140 195.250 137.460 195.310 ;
        RECT 140.835 195.250 141.125 195.295 ;
        RECT 152.780 195.250 153.100 195.310 ;
        RECT 137.140 195.110 153.100 195.250 ;
        RECT 137.140 195.050 137.460 195.110 ;
        RECT 140.835 195.065 141.125 195.110 ;
        RECT 152.780 195.050 153.100 195.110 ;
        RECT 124.735 194.910 125.025 194.955 ;
        RECT 125.180 194.910 125.500 194.970 ;
        RECT 125.655 194.910 125.945 194.955 ;
        RECT 124.735 194.770 125.945 194.910 ;
        RECT 124.735 194.725 125.025 194.770 ;
        RECT 125.180 194.710 125.500 194.770 ;
        RECT 125.655 194.725 125.945 194.770 ;
        RECT 126.100 194.910 126.420 194.970 ;
        RECT 128.415 194.910 128.705 194.955 ;
        RECT 126.100 194.770 127.710 194.910 ;
        RECT 126.100 194.710 126.420 194.770 ;
        RECT 127.570 194.570 127.710 194.770 ;
        RECT 128.415 194.770 141.050 194.910 ;
        RECT 128.415 194.725 128.705 194.770 ;
        RECT 129.795 194.570 130.085 194.615 ;
        RECT 122.970 194.430 127.250 194.570 ;
        RECT 127.570 194.430 130.085 194.570 ;
        RECT 99.880 194.030 100.200 194.290 ;
        RECT 106.780 194.230 107.100 194.290 ;
        RECT 122.510 194.230 122.650 194.385 ;
        RECT 127.110 194.230 127.250 194.430 ;
        RECT 129.795 194.385 130.085 194.430 ;
        RECT 131.160 194.570 131.480 194.630 ;
        RECT 133.475 194.570 133.765 194.615 ;
        RECT 131.160 194.430 133.765 194.570 ;
        RECT 131.160 194.370 131.480 194.430 ;
        RECT 133.475 194.385 133.765 194.430 ;
        RECT 133.935 194.385 134.225 194.615 ;
        RECT 128.415 194.230 128.705 194.275 ;
        RECT 106.780 194.090 121.270 194.230 ;
        RECT 106.780 194.030 107.100 194.090 ;
        RECT 100.800 193.890 101.120 193.950 ;
        RECT 99.100 193.750 101.120 193.890 ;
        RECT 100.800 193.690 101.120 193.750 ;
        RECT 103.560 193.890 103.880 193.950 ;
        RECT 114.600 193.890 114.920 193.950 ;
        RECT 103.560 193.750 114.920 193.890 ;
        RECT 103.560 193.690 103.880 193.750 ;
        RECT 114.600 193.690 114.920 193.750 ;
        RECT 117.820 193.690 118.140 193.950 ;
        RECT 121.130 193.890 121.270 194.090 ;
        RECT 122.510 194.090 126.790 194.230 ;
        RECT 127.110 194.090 128.705 194.230 ;
        RECT 134.010 194.230 134.150 194.385 ;
        RECT 134.380 194.370 134.700 194.630 ;
        RECT 134.840 194.570 135.160 194.630 ;
        RECT 135.315 194.570 135.605 194.615 ;
        RECT 134.840 194.430 135.605 194.570 ;
        RECT 134.840 194.370 135.160 194.430 ;
        RECT 135.315 194.385 135.605 194.430 ;
        RECT 135.775 194.385 136.065 194.615 ;
        RECT 136.220 194.570 136.540 194.630 ;
        RECT 136.695 194.570 136.985 194.615 ;
        RECT 136.220 194.430 136.985 194.570 ;
        RECT 135.905 194.230 136.045 194.385 ;
        RECT 136.220 194.370 136.540 194.430 ;
        RECT 136.695 194.385 136.985 194.430 ;
        RECT 139.915 194.385 140.205 194.615 ;
        RECT 134.010 194.090 136.045 194.230 ;
        RECT 122.510 193.890 122.650 194.090 ;
        RECT 121.130 193.750 122.650 193.890 ;
        RECT 83.780 193.550 84.100 193.610 ;
        RECT 73.290 193.410 84.100 193.550 ;
        RECT 71.375 193.365 71.665 193.410 ;
        RECT 71.820 193.350 72.140 193.410 ;
        RECT 83.780 193.350 84.100 193.410 ;
        RECT 84.255 193.550 84.545 193.595 ;
        RECT 84.700 193.550 85.020 193.610 ;
        RECT 85.620 193.550 85.940 193.610 ;
        RECT 84.255 193.410 85.940 193.550 ;
        RECT 84.255 193.365 84.545 193.410 ;
        RECT 84.700 193.350 85.020 193.410 ;
        RECT 85.620 193.350 85.940 193.410 ;
        RECT 87.000 193.350 87.320 193.610 ;
        RECT 89.760 193.550 90.080 193.610 ;
        RECT 92.980 193.550 93.300 193.610 ;
        RECT 89.760 193.410 93.300 193.550 ;
        RECT 89.760 193.350 90.080 193.410 ;
        RECT 92.980 193.350 93.300 193.410 ;
        RECT 98.040 193.550 98.360 193.610 ;
        RECT 106.320 193.550 106.640 193.610 ;
        RECT 98.040 193.410 106.640 193.550 ;
        RECT 98.040 193.350 98.360 193.410 ;
        RECT 106.320 193.350 106.640 193.410 ;
        RECT 110.920 193.550 111.240 193.610 ;
        RECT 111.855 193.550 112.145 193.595 ;
        RECT 110.920 193.410 112.145 193.550 ;
        RECT 110.920 193.350 111.240 193.410 ;
        RECT 111.855 193.365 112.145 193.410 ;
        RECT 112.775 193.550 113.065 193.595 ;
        RECT 113.680 193.550 114.000 193.610 ;
        RECT 112.775 193.410 114.000 193.550 ;
        RECT 112.775 193.365 113.065 193.410 ;
        RECT 113.680 193.350 114.000 193.410 ;
        RECT 114.140 193.350 114.460 193.610 ;
        RECT 117.910 193.550 118.050 193.690 ;
        RECT 122.880 193.550 123.200 193.610 ;
        RECT 123.355 193.550 123.645 193.595 ;
        RECT 126.100 193.550 126.420 193.610 ;
        RECT 126.650 193.595 126.790 194.090 ;
        RECT 128.415 194.045 128.705 194.090 ;
        RECT 134.930 193.950 135.070 194.090 ;
        RECT 127.480 193.690 127.800 193.950 ;
        RECT 128.860 193.890 129.180 193.950 ;
        RECT 129.335 193.890 129.625 193.935 ;
        RECT 128.860 193.750 129.625 193.890 ;
        RECT 128.860 193.690 129.180 193.750 ;
        RECT 129.335 193.705 129.625 193.750 ;
        RECT 134.840 193.690 135.160 193.950 ;
        RECT 135.760 193.890 136.080 193.950 ;
        RECT 138.060 193.890 138.380 193.950 ;
        RECT 135.760 193.750 138.380 193.890 ;
        RECT 135.760 193.690 136.080 193.750 ;
        RECT 138.060 193.690 138.380 193.750 ;
        RECT 117.910 193.410 126.420 193.550 ;
        RECT 122.880 193.350 123.200 193.410 ;
        RECT 123.355 193.365 123.645 193.410 ;
        RECT 126.100 193.350 126.420 193.410 ;
        RECT 126.575 193.550 126.865 193.595 ;
        RECT 139.990 193.550 140.130 194.385 ;
        RECT 140.910 194.230 141.050 194.770 ;
        RECT 141.370 194.770 144.270 194.910 ;
        RECT 141.370 194.630 141.510 194.770 ;
        RECT 141.280 194.370 141.600 194.630 ;
        RECT 142.660 194.570 142.980 194.630 ;
        RECT 144.130 194.615 144.270 194.770 ;
        RECT 144.590 194.770 146.570 194.910 ;
        RECT 143.135 194.570 143.425 194.615 ;
        RECT 142.660 194.430 143.425 194.570 ;
        RECT 142.660 194.370 142.980 194.430 ;
        RECT 143.135 194.385 143.425 194.430 ;
        RECT 144.055 194.385 144.345 194.615 ;
        RECT 144.590 194.230 144.730 194.770 ;
        RECT 145.435 194.385 145.725 194.615 ;
        RECT 140.910 194.090 144.730 194.230 ;
        RECT 144.040 193.690 144.360 193.950 ;
        RECT 144.500 193.690 144.820 193.950 ;
        RECT 141.740 193.550 142.060 193.610 ;
        RECT 126.575 193.410 142.060 193.550 ;
        RECT 145.510 193.550 145.650 194.385 ;
        RECT 145.880 194.370 146.200 194.630 ;
        RECT 146.430 194.615 146.570 194.770 ;
        RECT 146.355 194.385 146.645 194.615 ;
        RECT 146.800 194.370 147.120 194.630 ;
        RECT 147.720 194.370 148.040 194.630 ;
        RECT 151.860 194.570 152.180 194.630 ;
        RECT 153.240 194.570 153.560 194.630 ;
        RECT 151.860 194.430 153.560 194.570 ;
        RECT 151.860 194.370 152.180 194.430 ;
        RECT 153.240 194.370 153.560 194.430 ;
        RECT 145.970 193.935 146.110 194.370 ;
        RECT 145.895 193.705 146.185 193.935 ;
        RECT 146.340 193.550 146.660 193.610 ;
        RECT 145.510 193.410 146.660 193.550 ;
        RECT 126.575 193.365 126.865 193.410 ;
        RECT 141.740 193.350 142.060 193.410 ;
        RECT 146.340 193.350 146.660 193.410 ;
        RECT 2.750 192.730 158.230 193.210 ;
        RECT 5.580 192.530 5.900 192.590 ;
        RECT 6.055 192.530 6.345 192.575 ;
        RECT 37.795 192.530 38.085 192.575 ;
        RECT 43.760 192.530 44.080 192.590 ;
        RECT 5.580 192.390 6.345 192.530 ;
        RECT 5.580 192.330 5.900 192.390 ;
        RECT 6.055 192.345 6.345 192.390 ;
        RECT 12.110 192.390 20.990 192.530 ;
        RECT 5.120 192.190 5.440 192.250 ;
        RECT 11.575 192.190 11.865 192.235 ;
        RECT 5.120 192.050 11.865 192.190 ;
        RECT 5.120 191.990 5.440 192.050 ;
        RECT 11.575 192.005 11.865 192.050 ;
        RECT 10.640 191.850 10.960 191.910 ;
        RECT 12.110 191.850 12.250 192.390 ;
        RECT 20.300 192.190 20.620 192.250 ;
        RECT 14.870 192.050 20.620 192.190 ;
        RECT 14.870 191.895 15.010 192.050 ;
        RECT 20.300 191.990 20.620 192.050 ;
        RECT 10.640 191.710 12.250 191.850 ;
        RECT 10.640 191.650 10.960 191.710 ;
        RECT 14.795 191.665 15.085 191.895 ;
        RECT 15.700 191.850 16.020 191.910 ;
        RECT 19.855 191.850 20.145 191.895 ;
        RECT 20.850 191.850 20.990 192.390 ;
        RECT 24.555 192.390 36.630 192.530 ;
        RECT 21.695 191.850 21.985 191.895 ;
        RECT 24.555 191.850 24.695 192.390 ;
        RECT 29.925 192.190 30.215 192.235 ;
        RECT 31.815 192.190 32.105 192.235 ;
        RECT 34.935 192.190 35.225 192.235 ;
        RECT 24.990 192.050 26.510 192.190 ;
        RECT 24.990 191.910 25.130 192.050 ;
        RECT 15.700 191.710 18.690 191.850 ;
        RECT 15.700 191.650 16.020 191.710 ;
        RECT 6.975 191.510 7.265 191.555 ;
        RECT 9.275 191.510 9.565 191.555 ;
        RECT 12.940 191.510 13.260 191.570 ;
        RECT 6.975 191.370 7.650 191.510 ;
        RECT 6.975 191.325 7.265 191.370 ;
        RECT 7.510 190.875 7.650 191.370 ;
        RECT 9.275 191.370 13.260 191.510 ;
        RECT 9.275 191.325 9.565 191.370 ;
        RECT 12.940 191.310 13.260 191.370 ;
        RECT 13.415 191.510 13.705 191.555 ;
        RECT 14.320 191.510 14.640 191.570 ;
        RECT 18.000 191.510 18.320 191.570 ;
        RECT 18.550 191.555 18.690 191.710 ;
        RECT 19.855 191.710 24.695 191.850 ;
        RECT 19.855 191.665 20.145 191.710 ;
        RECT 21.695 191.665 21.985 191.710 ;
        RECT 24.900 191.650 25.220 191.910 ;
        RECT 25.820 191.650 26.140 191.910 ;
        RECT 26.370 191.895 26.510 192.050 ;
        RECT 29.925 192.050 35.225 192.190 ;
        RECT 29.925 192.005 30.215 192.050 ;
        RECT 31.815 192.005 32.105 192.050 ;
        RECT 34.935 192.005 35.225 192.050 ;
        RECT 36.490 191.910 36.630 192.390 ;
        RECT 37.795 192.390 44.080 192.530 ;
        RECT 37.795 192.345 38.085 192.390 ;
        RECT 26.295 191.665 26.585 191.895 ;
        RECT 27.660 191.850 27.980 191.910 ;
        RECT 29.055 191.850 29.345 191.895 ;
        RECT 27.660 191.710 29.345 191.850 ;
        RECT 27.660 191.650 27.980 191.710 ;
        RECT 29.055 191.665 29.345 191.710 ;
        RECT 36.400 191.850 36.720 191.910 ;
        RECT 38.700 191.850 39.020 191.910 ;
        RECT 39.250 191.895 39.390 192.390 ;
        RECT 43.760 192.330 44.080 192.390 ;
        RECT 44.335 192.390 45.370 192.530 ;
        RECT 41.935 192.190 42.225 192.235 ;
        RECT 43.300 192.190 43.620 192.250 ;
        RECT 41.935 192.050 43.620 192.190 ;
        RECT 41.935 192.005 42.225 192.050 ;
        RECT 43.300 191.990 43.620 192.050 ;
        RECT 36.400 191.710 39.020 191.850 ;
        RECT 36.400 191.650 36.720 191.710 ;
        RECT 38.700 191.650 39.020 191.710 ;
        RECT 39.175 191.665 39.465 191.895 ;
        RECT 44.335 191.850 44.475 192.390 ;
        RECT 45.230 191.895 45.370 192.390 ;
        RECT 46.520 192.330 46.840 192.590 ;
        RECT 46.980 192.330 47.300 192.590 ;
        RECT 48.360 192.530 48.680 192.590 ;
        RECT 49.280 192.530 49.600 192.590 ;
        RECT 48.360 192.390 49.600 192.530 ;
        RECT 48.360 192.330 48.680 192.390 ;
        RECT 49.280 192.330 49.600 192.390 ;
        RECT 54.340 192.330 54.660 192.590 ;
        RECT 56.640 192.530 56.960 192.590 ;
        RECT 57.115 192.530 57.405 192.575 ;
        RECT 56.640 192.390 57.405 192.530 ;
        RECT 56.640 192.330 56.960 192.390 ;
        RECT 57.115 192.345 57.405 192.390 ;
        RECT 59.860 192.530 60.180 192.590 ;
        RECT 61.255 192.530 61.545 192.575 ;
        RECT 59.860 192.390 61.545 192.530 ;
        RECT 59.860 192.330 60.180 192.390 ;
        RECT 61.255 192.345 61.545 192.390 ;
        RECT 66.760 192.530 67.080 192.590 ;
        RECT 72.740 192.530 73.060 192.590 ;
        RECT 73.215 192.530 73.505 192.575 ;
        RECT 66.760 192.390 72.510 192.530 ;
        RECT 66.760 192.330 67.080 192.390 ;
        RECT 47.070 192.190 47.210 192.330 ;
        RECT 48.785 192.190 49.075 192.235 ;
        RECT 50.675 192.190 50.965 192.235 ;
        RECT 53.795 192.190 54.085 192.235 ;
        RECT 47.070 192.050 48.360 192.190 ;
        RECT 39.710 191.710 44.475 191.850 ;
        RECT 13.415 191.370 14.640 191.510 ;
        RECT 13.415 191.325 13.705 191.370 ;
        RECT 14.320 191.310 14.640 191.370 ;
        RECT 15.790 191.370 18.320 191.510 ;
        RECT 9.735 191.170 10.025 191.215 ;
        RECT 15.790 191.170 15.930 191.370 ;
        RECT 18.000 191.310 18.320 191.370 ;
        RECT 18.475 191.510 18.765 191.555 ;
        RECT 26.740 191.510 27.060 191.570 ;
        RECT 18.475 191.370 27.060 191.510 ;
        RECT 18.475 191.325 18.765 191.370 ;
        RECT 26.740 191.310 27.060 191.370 ;
        RECT 29.520 191.510 29.810 191.555 ;
        RECT 31.355 191.510 31.645 191.555 ;
        RECT 34.935 191.510 35.225 191.555 ;
        RECT 29.520 191.370 35.225 191.510 ;
        RECT 29.520 191.325 29.810 191.370 ;
        RECT 31.355 191.325 31.645 191.370 ;
        RECT 34.935 191.325 35.225 191.370 ;
        RECT 36.015 191.510 36.305 191.530 ;
        RECT 36.860 191.510 37.180 191.570 ;
        RECT 36.015 191.370 37.180 191.510 ;
        RECT 38.790 191.510 38.930 191.650 ;
        RECT 39.710 191.510 39.850 191.710 ;
        RECT 45.155 191.665 45.445 191.895 ;
        RECT 48.220 191.850 48.360 192.050 ;
        RECT 48.785 192.050 54.085 192.190 ;
        RECT 54.430 192.190 54.570 192.330 ;
        RECT 64.000 192.190 64.320 192.250 ;
        RECT 69.980 192.190 70.300 192.250 ;
        RECT 54.430 192.050 61.470 192.190 ;
        RECT 48.785 192.005 49.075 192.050 ;
        RECT 50.675 192.005 50.965 192.050 ;
        RECT 53.795 192.005 54.085 192.050 ;
        RECT 49.295 191.850 49.585 191.895 ;
        RECT 48.220 191.710 49.585 191.850 ;
        RECT 49.295 191.665 49.585 191.710 ;
        RECT 55.260 191.850 55.580 191.910 ;
        RECT 56.655 191.850 56.945 191.895 ;
        RECT 59.400 191.850 59.720 191.910 ;
        RECT 59.875 191.850 60.165 191.895 ;
        RECT 55.260 191.710 59.170 191.850 ;
        RECT 55.260 191.650 55.580 191.710 ;
        RECT 56.655 191.665 56.945 191.710 ;
        RECT 38.790 191.370 39.850 191.510 ;
        RECT 18.935 191.170 19.225 191.215 ;
        RECT 9.735 191.030 15.930 191.170 ;
        RECT 16.250 191.030 19.225 191.170 ;
        RECT 9.735 190.985 10.025 191.030 ;
        RECT 16.250 190.890 16.390 191.030 ;
        RECT 18.935 190.985 19.225 191.030 ;
        RECT 22.155 191.170 22.445 191.215 ;
        RECT 28.120 191.170 28.440 191.230 ;
        RECT 22.155 191.030 28.440 191.170 ;
        RECT 22.155 190.985 22.445 191.030 ;
        RECT 28.120 190.970 28.440 191.030 ;
        RECT 30.420 190.970 30.740 191.230 ;
        RECT 36.015 191.215 36.305 191.370 ;
        RECT 36.860 191.310 37.180 191.370 ;
        RECT 40.080 191.310 40.400 191.570 ;
        RECT 41.015 191.510 41.305 191.555 ;
        RECT 42.380 191.510 42.700 191.570 ;
        RECT 41.015 191.370 42.700 191.510 ;
        RECT 41.015 191.325 41.305 191.370 ;
        RECT 42.380 191.310 42.700 191.370 ;
        RECT 46.520 191.560 46.840 191.570 ;
        RECT 46.520 191.510 47.210 191.560 ;
        RECT 47.900 191.510 48.220 191.570 ;
        RECT 59.030 191.555 59.170 191.710 ;
        RECT 59.400 191.710 60.165 191.850 ;
        RECT 59.400 191.650 59.720 191.710 ;
        RECT 59.875 191.665 60.165 191.710 ;
        RECT 61.330 191.555 61.470 192.050 ;
        RECT 64.000 192.050 70.300 192.190 ;
        RECT 64.000 191.990 64.320 192.050 ;
        RECT 69.980 191.990 70.300 192.050 ;
        RECT 64.920 191.850 65.240 191.910 ;
        RECT 65.395 191.850 65.685 191.895 ;
        RECT 64.920 191.710 65.685 191.850 ;
        RECT 64.920 191.650 65.240 191.710 ;
        RECT 65.395 191.665 65.685 191.710 ;
        RECT 66.775 191.850 67.065 191.895 ;
        RECT 68.140 191.850 68.460 191.910 ;
        RECT 66.775 191.710 68.460 191.850 ;
        RECT 66.775 191.665 67.065 191.710 ;
        RECT 68.140 191.650 68.460 191.710 ;
        RECT 46.520 191.420 48.220 191.510 ;
        RECT 46.520 191.310 46.840 191.420 ;
        RECT 47.070 191.370 48.220 191.420 ;
        RECT 47.900 191.310 48.220 191.370 ;
        RECT 48.380 191.510 48.670 191.555 ;
        RECT 50.215 191.510 50.505 191.555 ;
        RECT 53.795 191.510 54.085 191.555 ;
        RECT 48.380 191.370 54.085 191.510 ;
        RECT 48.380 191.325 48.670 191.370 ;
        RECT 50.215 191.325 50.505 191.370 ;
        RECT 53.795 191.325 54.085 191.370 ;
        RECT 32.715 191.170 33.365 191.215 ;
        RECT 36.015 191.170 36.605 191.215 ;
        RECT 46.980 191.170 47.300 191.230 ;
        RECT 49.740 191.170 50.060 191.230 ;
        RECT 54.875 191.215 55.165 191.530 ;
        RECT 58.955 191.325 59.245 191.555 ;
        RECT 61.255 191.325 61.545 191.555 ;
        RECT 62.175 191.325 62.465 191.555 ;
        RECT 51.575 191.170 52.225 191.215 ;
        RECT 54.875 191.170 55.465 191.215 ;
        RECT 59.415 191.170 59.705 191.215 ;
        RECT 32.715 191.030 36.605 191.170 ;
        RECT 32.715 190.985 33.365 191.030 ;
        RECT 36.315 190.985 36.605 191.030 ;
        RECT 42.470 191.030 46.750 191.170 ;
        RECT 7.435 190.645 7.725 190.875 ;
        RECT 13.875 190.830 14.165 190.875 ;
        RECT 16.160 190.830 16.480 190.890 ;
        RECT 13.875 190.690 16.480 190.830 ;
        RECT 13.875 190.645 14.165 190.690 ;
        RECT 16.160 190.630 16.480 190.690 ;
        RECT 16.620 190.630 16.940 190.890 ;
        RECT 22.615 190.830 22.905 190.875 ;
        RECT 23.060 190.830 23.380 190.890 ;
        RECT 22.615 190.690 23.380 190.830 ;
        RECT 22.615 190.645 22.905 190.690 ;
        RECT 23.060 190.630 23.380 190.690 ;
        RECT 24.455 190.830 24.745 190.875 ;
        RECT 25.820 190.830 26.140 190.890 ;
        RECT 24.455 190.690 26.140 190.830 ;
        RECT 24.455 190.645 24.745 190.690 ;
        RECT 25.820 190.630 26.140 190.690 ;
        RECT 28.595 190.830 28.885 190.875 ;
        RECT 42.470 190.830 42.610 191.030 ;
        RECT 28.595 190.690 42.610 190.830 ;
        RECT 42.840 190.830 43.160 190.890 ;
        RECT 43.775 190.830 44.065 190.875 ;
        RECT 42.840 190.690 44.065 190.830 ;
        RECT 28.595 190.645 28.885 190.690 ;
        RECT 42.840 190.630 43.160 190.690 ;
        RECT 43.775 190.645 44.065 190.690 ;
        RECT 44.235 190.830 44.525 190.875 ;
        RECT 44.680 190.830 45.000 190.890 ;
        RECT 44.235 190.690 45.000 190.830 ;
        RECT 46.610 190.830 46.750 191.030 ;
        RECT 46.980 191.030 55.465 191.170 ;
        RECT 46.980 190.970 47.300 191.030 ;
        RECT 49.740 190.970 50.060 191.030 ;
        RECT 51.575 190.985 52.225 191.030 ;
        RECT 55.175 190.985 55.465 191.030 ;
        RECT 55.810 191.030 59.705 191.170 ;
        RECT 55.810 190.830 55.950 191.030 ;
        RECT 59.415 190.985 59.705 191.030 ;
        RECT 46.610 190.690 55.950 190.830 ;
        RECT 56.180 190.830 56.500 190.890 ;
        RECT 62.250 190.830 62.390 191.325 ;
        RECT 64.350 191.170 64.640 191.215 ;
        RECT 71.820 191.170 72.140 191.230 ;
        RECT 64.350 191.030 72.140 191.170 ;
        RECT 72.370 191.170 72.510 192.390 ;
        RECT 72.740 192.390 73.505 192.530 ;
        RECT 72.740 192.330 73.060 192.390 ;
        RECT 73.215 192.345 73.505 192.390 ;
        RECT 74.135 192.530 74.425 192.575 ;
        RECT 74.580 192.530 74.900 192.590 ;
        RECT 74.135 192.390 74.900 192.530 ;
        RECT 74.135 192.345 74.425 192.390 ;
        RECT 74.580 192.330 74.900 192.390 ;
        RECT 81.480 192.530 81.800 192.590 ;
        RECT 86.540 192.530 86.860 192.590 ;
        RECT 81.480 192.390 86.860 192.530 ;
        RECT 81.480 192.330 81.800 192.390 ;
        RECT 86.540 192.330 86.860 192.390 ;
        RECT 89.315 192.530 89.605 192.575 ;
        RECT 89.315 192.390 94.590 192.530 ;
        RECT 89.315 192.345 89.605 192.390 ;
        RECT 76.880 192.190 77.200 192.250 ;
        RECT 81.940 192.190 82.260 192.250 ;
        RECT 72.830 192.050 82.260 192.190 ;
        RECT 72.830 191.555 72.970 192.050 ;
        RECT 76.880 191.990 77.200 192.050 ;
        RECT 81.940 191.990 82.260 192.050 ;
        RECT 83.780 192.190 84.100 192.250 ;
        RECT 87.000 192.190 87.320 192.250 ;
        RECT 87.935 192.190 88.225 192.235 ;
        RECT 83.780 192.050 88.225 192.190 ;
        RECT 83.780 191.990 84.100 192.050 ;
        RECT 87.000 191.990 87.320 192.050 ;
        RECT 87.935 192.005 88.225 192.050 ;
        RECT 89.760 192.190 90.080 192.250 ;
        RECT 90.680 192.190 91.000 192.250 ;
        RECT 89.760 192.050 91.000 192.190 ;
        RECT 89.760 191.990 90.080 192.050 ;
        RECT 90.680 191.990 91.000 192.050 ;
        RECT 93.440 191.990 93.760 192.250 ;
        RECT 78.720 191.850 79.040 191.910 ;
        RECT 93.530 191.850 93.670 191.990 ;
        RECT 74.210 191.710 93.670 191.850 ;
        RECT 72.755 191.325 73.045 191.555 ;
        RECT 73.660 191.310 73.980 191.570 ;
        RECT 74.210 191.555 74.350 191.710 ;
        RECT 78.720 191.650 79.040 191.710 ;
        RECT 74.135 191.325 74.425 191.555 ;
        RECT 75.055 191.510 75.345 191.555 ;
        RECT 76.420 191.510 76.740 191.570 ;
        RECT 75.055 191.370 76.740 191.510 ;
        RECT 75.055 191.325 75.345 191.370 ;
        RECT 76.420 191.310 76.740 191.370 ;
        RECT 86.095 191.510 86.385 191.555 ;
        RECT 86.540 191.510 86.860 191.570 ;
        RECT 86.095 191.370 86.860 191.510 ;
        RECT 86.095 191.325 86.385 191.370 ;
        RECT 86.540 191.310 86.860 191.370 ;
        RECT 87.000 191.310 87.320 191.570 ;
        RECT 87.460 191.310 87.780 191.570 ;
        RECT 88.395 191.510 88.685 191.555 ;
        RECT 88.840 191.510 89.160 191.570 ;
        RECT 88.395 191.370 89.160 191.510 ;
        RECT 88.395 191.325 88.685 191.370 ;
        RECT 88.840 191.310 89.160 191.370 ;
        RECT 89.760 191.510 90.080 191.570 ;
        RECT 92.980 191.510 93.300 191.570 ;
        RECT 94.450 191.555 94.590 192.390 ;
        RECT 94.820 192.330 95.140 192.590 ;
        RECT 96.200 192.530 96.520 192.590 ;
        RECT 97.135 192.530 97.425 192.575 ;
        RECT 96.200 192.390 97.425 192.530 ;
        RECT 96.200 192.330 96.520 192.390 ;
        RECT 97.135 192.345 97.425 192.390 ;
        RECT 104.480 192.530 104.800 192.590 ;
        RECT 105.875 192.530 106.165 192.575 ;
        RECT 109.080 192.530 109.400 192.590 ;
        RECT 104.480 192.390 106.165 192.530 ;
        RECT 104.480 192.330 104.800 192.390 ;
        RECT 105.875 192.345 106.165 192.390 ;
        RECT 106.410 192.390 109.400 192.530 ;
        RECT 94.910 191.850 95.050 192.330 ;
        RECT 96.675 192.190 96.965 192.235 ;
        RECT 106.410 192.190 106.550 192.390 ;
        RECT 109.080 192.330 109.400 192.390 ;
        RECT 109.540 192.530 109.860 192.590 ;
        RECT 114.615 192.530 114.905 192.575 ;
        RECT 115.060 192.530 115.380 192.590 ;
        RECT 109.540 192.390 113.450 192.530 ;
        RECT 109.540 192.330 109.860 192.390 ;
        RECT 96.675 192.050 106.550 192.190 ;
        RECT 108.175 192.190 108.465 192.235 ;
        RECT 113.310 192.190 113.450 192.390 ;
        RECT 114.615 192.390 115.380 192.530 ;
        RECT 114.615 192.345 114.905 192.390 ;
        RECT 115.060 192.330 115.380 192.390 ;
        RECT 115.520 192.530 115.840 192.590 ;
        RECT 116.900 192.530 117.220 192.590 ;
        RECT 115.520 192.390 117.220 192.530 ;
        RECT 115.520 192.330 115.840 192.390 ;
        RECT 116.900 192.330 117.220 192.390 ;
        RECT 121.040 192.330 121.360 192.590 ;
        RECT 121.960 192.530 122.280 192.590 ;
        RECT 128.860 192.530 129.180 192.590 ;
        RECT 121.960 192.390 129.180 192.530 ;
        RECT 121.960 192.330 122.280 192.390 ;
        RECT 128.860 192.330 129.180 192.390 ;
        RECT 130.240 192.530 130.560 192.590 ;
        RECT 146.800 192.530 147.120 192.590 ;
        RECT 148.180 192.530 148.500 192.590 ;
        RECT 130.240 192.390 148.500 192.530 ;
        RECT 130.240 192.330 130.560 192.390 ;
        RECT 146.800 192.330 147.120 192.390 ;
        RECT 148.180 192.330 148.500 192.390 ;
        RECT 150.940 192.330 151.260 192.590 ;
        RECT 151.875 192.345 152.165 192.575 ;
        RECT 121.130 192.190 121.270 192.330 ;
        RECT 108.175 192.050 112.990 192.190 ;
        RECT 113.310 192.050 121.270 192.190 ;
        RECT 96.675 192.005 96.965 192.050 ;
        RECT 108.175 192.005 108.465 192.050 ;
        RECT 96.200 191.850 96.520 191.910 ;
        RECT 100.340 191.850 100.660 191.910 ;
        RECT 94.910 191.710 98.730 191.850 ;
        RECT 96.200 191.650 96.520 191.710 ;
        RECT 89.760 191.370 93.300 191.510 ;
        RECT 89.760 191.310 90.080 191.370 ;
        RECT 92.980 191.310 93.300 191.370 ;
        RECT 93.455 191.325 93.745 191.555 ;
        RECT 94.375 191.325 94.665 191.555 ;
        RECT 91.600 191.170 91.920 191.230 ;
        RECT 93.530 191.170 93.670 191.325 ;
        RECT 94.820 191.310 95.140 191.570 ;
        RECT 95.280 191.310 95.600 191.570 ;
        RECT 98.590 191.555 98.730 191.710 ;
        RECT 100.340 191.710 103.790 191.850 ;
        RECT 100.340 191.650 100.660 191.710 ;
        RECT 98.060 191.230 98.350 191.445 ;
        RECT 98.515 191.325 98.805 191.555 ;
        RECT 98.975 191.510 99.265 191.555 ;
        RECT 98.975 191.370 101.950 191.510 ;
        RECT 98.975 191.325 99.265 191.370 ;
        RECT 97.120 191.170 97.440 191.230 ;
        RECT 72.370 191.030 93.670 191.170 ;
        RECT 93.990 191.030 97.440 191.170 ;
        RECT 64.350 190.985 64.640 191.030 ;
        RECT 71.820 190.970 72.140 191.030 ;
        RECT 91.600 190.970 91.920 191.030 ;
        RECT 56.180 190.690 62.390 190.830 ;
        RECT 44.235 190.645 44.525 190.690 ;
        RECT 44.680 190.630 45.000 190.690 ;
        RECT 56.180 190.630 56.500 190.690 ;
        RECT 63.540 190.630 63.860 190.890 ;
        RECT 64.935 190.830 65.225 190.875 ;
        RECT 65.380 190.830 65.700 190.890 ;
        RECT 67.220 190.830 67.540 190.890 ;
        RECT 64.935 190.690 67.540 190.830 ;
        RECT 64.935 190.645 65.225 190.690 ;
        RECT 65.380 190.630 65.700 190.690 ;
        RECT 67.220 190.630 67.540 190.690 ;
        RECT 87.920 190.830 88.240 190.890 ;
        RECT 93.990 190.830 94.130 191.030 ;
        RECT 97.120 190.970 97.440 191.030 ;
        RECT 98.040 190.970 98.360 191.230 ;
        RECT 87.920 190.690 94.130 190.830 ;
        RECT 94.360 190.830 94.680 190.890 ;
        RECT 99.050 190.830 99.190 191.325 ;
        RECT 101.810 191.230 101.950 191.370 ;
        RECT 102.655 191.325 102.945 191.555 ;
        RECT 99.665 191.170 99.955 191.215 ;
        RECT 100.800 191.170 101.120 191.230 ;
        RECT 99.665 191.030 101.120 191.170 ;
        RECT 99.665 190.985 99.955 191.030 ;
        RECT 100.800 190.970 101.120 191.030 ;
        RECT 101.720 190.970 102.040 191.230 ;
        RECT 102.730 191.170 102.870 191.325 ;
        RECT 103.100 191.310 103.420 191.570 ;
        RECT 103.650 191.510 103.790 191.710 ;
        RECT 104.020 191.650 104.340 191.910 ;
        RECT 104.940 191.650 105.260 191.910 ;
        RECT 105.860 191.650 106.180 191.910 ;
        RECT 106.320 191.650 106.640 191.910 ;
        RECT 105.030 191.510 105.170 191.650 ;
        RECT 105.950 191.510 106.090 191.650 ;
        RECT 103.650 191.370 105.170 191.510 ;
        RECT 105.490 191.370 106.090 191.510 ;
        RECT 107.255 191.510 107.545 191.555 ;
        RECT 109.540 191.510 109.860 191.570 ;
        RECT 112.850 191.555 112.990 192.050 ;
        RECT 135.300 191.990 135.620 192.250 ;
        RECT 143.120 192.190 143.440 192.250 ;
        RECT 135.850 192.050 143.440 192.190 ;
        RECT 113.695 191.850 113.985 191.895 ;
        RECT 114.140 191.850 114.460 191.910 ;
        RECT 128.400 191.850 128.720 191.910 ;
        RECT 113.695 191.710 114.460 191.850 ;
        RECT 113.695 191.665 113.985 191.710 ;
        RECT 114.140 191.650 114.460 191.710 ;
        RECT 115.150 191.710 128.720 191.850 ;
        RECT 114.600 191.555 114.920 191.570 ;
        RECT 107.255 191.370 109.860 191.510 ;
        RECT 102.730 191.030 103.330 191.170 ;
        RECT 94.360 190.690 99.190 190.830 ;
        RECT 103.190 190.830 103.330 191.030 ;
        RECT 104.940 190.830 105.260 190.890 ;
        RECT 105.490 190.830 105.630 191.370 ;
        RECT 107.255 191.325 107.545 191.370 ;
        RECT 109.540 191.310 109.860 191.370 ;
        RECT 112.775 191.325 113.065 191.555 ;
        RECT 114.600 191.510 114.965 191.555 ;
        RECT 115.150 191.510 115.290 191.710 ;
        RECT 128.400 191.650 128.720 191.710 ;
        RECT 128.860 191.850 129.180 191.910 ;
        RECT 135.850 191.850 135.990 192.050 ;
        RECT 143.120 191.990 143.440 192.050 ;
        RECT 128.860 191.710 135.990 191.850 ;
        RECT 128.860 191.650 129.180 191.710 ;
        RECT 137.600 191.650 137.920 191.910 ;
        RECT 138.075 191.850 138.365 191.895 ;
        RECT 140.820 191.850 141.140 191.910 ;
        RECT 138.075 191.710 141.140 191.850 ;
        RECT 138.075 191.665 138.365 191.710 ;
        RECT 140.820 191.650 141.140 191.710 ;
        RECT 150.940 191.850 151.260 191.910 ;
        RECT 151.950 191.850 152.090 192.345 ;
        RECT 150.940 191.710 152.090 191.850 ;
        RECT 150.940 191.650 151.260 191.710 ;
        RECT 114.600 191.370 115.290 191.510 ;
        RECT 117.820 191.510 118.140 191.570 ;
        RECT 120.135 191.510 120.425 191.555 ;
        RECT 117.820 191.370 120.425 191.510 ;
        RECT 114.600 191.325 114.965 191.370 ;
        RECT 114.600 191.310 114.920 191.325 ;
        RECT 117.820 191.310 118.140 191.370 ;
        RECT 120.135 191.325 120.425 191.370 ;
        RECT 120.595 191.510 120.885 191.555 ;
        RECT 143.580 191.510 143.900 191.570 ;
        RECT 120.595 191.370 143.900 191.510 ;
        RECT 120.595 191.325 120.885 191.370 ;
        RECT 105.860 191.170 106.180 191.230 ;
        RECT 107.700 191.170 108.020 191.230 ;
        RECT 105.860 191.030 108.020 191.170 ;
        RECT 105.860 190.970 106.180 191.030 ;
        RECT 107.700 190.970 108.020 191.030 ;
        RECT 113.235 191.170 113.525 191.215 ;
        RECT 119.660 191.170 119.980 191.230 ;
        RECT 120.670 191.170 120.810 191.325 ;
        RECT 143.580 191.310 143.900 191.370 ;
        RECT 151.860 191.310 152.180 191.570 ;
        RECT 152.335 191.510 152.625 191.555 ;
        RECT 153.700 191.510 154.020 191.570 ;
        RECT 152.335 191.370 154.020 191.510 ;
        RECT 152.335 191.325 152.625 191.370 ;
        RECT 113.235 191.030 119.430 191.170 ;
        RECT 113.235 190.985 113.525 191.030 ;
        RECT 103.190 190.690 105.630 190.830 ;
        RECT 106.320 190.830 106.640 190.890 ;
        RECT 116.440 190.830 116.760 190.890 ;
        RECT 119.290 190.875 119.430 191.030 ;
        RECT 119.660 191.030 120.810 191.170 ;
        RECT 121.515 191.170 121.805 191.215 ;
        RECT 133.460 191.170 133.780 191.230 ;
        RECT 137.140 191.170 137.460 191.230 ;
        RECT 121.515 191.030 122.190 191.170 ;
        RECT 119.660 190.970 119.980 191.030 ;
        RECT 121.515 190.985 121.805 191.030 ;
        RECT 122.050 190.890 122.190 191.030 ;
        RECT 133.460 191.030 137.460 191.170 ;
        RECT 133.460 190.970 133.780 191.030 ;
        RECT 137.140 190.970 137.460 191.030 ;
        RECT 148.640 191.170 148.960 191.230 ;
        RECT 152.410 191.170 152.550 191.325 ;
        RECT 153.700 191.310 154.020 191.370 ;
        RECT 148.640 191.030 152.550 191.170 ;
        RECT 148.640 190.970 148.960 191.030 ;
        RECT 153.255 190.985 153.545 191.215 ;
        RECT 106.320 190.690 116.760 190.830 ;
        RECT 87.920 190.630 88.240 190.690 ;
        RECT 94.360 190.630 94.680 190.690 ;
        RECT 104.940 190.630 105.260 190.690 ;
        RECT 106.320 190.630 106.640 190.690 ;
        RECT 116.440 190.630 116.760 190.690 ;
        RECT 119.215 190.645 119.505 190.875 ;
        RECT 121.960 190.630 122.280 190.890 ;
        RECT 137.600 190.630 137.920 190.890 ;
        RECT 152.320 190.830 152.640 190.890 ;
        RECT 153.330 190.830 153.470 190.985 ;
        RECT 152.320 190.690 153.470 190.830 ;
        RECT 152.320 190.630 152.640 190.690 ;
        RECT 2.750 190.010 159.030 190.490 ;
        RECT 5.120 189.610 5.440 189.870 ;
        RECT 5.595 189.625 5.885 189.855 ;
        RECT 25.835 189.810 26.125 189.855 ;
        RECT 26.740 189.810 27.060 189.870 ;
        RECT 16.710 189.670 24.210 189.810 ;
        RECT 4.675 189.130 4.965 189.175 ;
        RECT 5.210 189.130 5.350 189.610 ;
        RECT 5.670 189.470 5.810 189.625 ;
        RECT 7.435 189.470 7.725 189.515 ;
        RECT 5.670 189.330 7.725 189.470 ;
        RECT 7.435 189.285 7.725 189.330 ;
        RECT 9.715 189.470 10.365 189.515 ;
        RECT 13.315 189.470 13.605 189.515 ;
        RECT 13.860 189.470 14.180 189.530 ;
        RECT 16.710 189.470 16.850 189.670 ;
        RECT 9.715 189.330 16.850 189.470 ;
        RECT 20.755 189.470 21.405 189.515 ;
        RECT 24.070 189.470 24.210 189.670 ;
        RECT 25.835 189.670 27.060 189.810 ;
        RECT 25.835 189.625 26.125 189.670 ;
        RECT 26.740 189.610 27.060 189.670 ;
        RECT 30.420 189.610 30.740 189.870 ;
        RECT 30.880 189.610 31.200 189.870 ;
        RECT 32.735 189.810 33.025 189.855 ;
        RECT 33.180 189.810 33.500 189.870 ;
        RECT 46.520 189.810 46.840 189.870 ;
        RECT 32.735 189.670 33.500 189.810 ;
        RECT 32.735 189.625 33.025 189.670 ;
        RECT 33.180 189.610 33.500 189.670 ;
        RECT 36.490 189.670 46.840 189.810 ;
        RECT 24.355 189.470 24.645 189.515 ;
        RECT 20.755 189.330 24.645 189.470 ;
        RECT 9.715 189.285 10.365 189.330 ;
        RECT 13.015 189.285 13.605 189.330 ;
        RECT 4.675 188.990 5.350 189.130 ;
        RECT 6.520 189.130 6.810 189.175 ;
        RECT 8.355 189.130 8.645 189.175 ;
        RECT 11.935 189.130 12.225 189.175 ;
        RECT 6.520 188.990 12.225 189.130 ;
        RECT 4.675 188.945 4.965 188.990 ;
        RECT 6.520 188.945 6.810 188.990 ;
        RECT 8.355 188.945 8.645 188.990 ;
        RECT 11.935 188.945 12.225 188.990 ;
        RECT 13.015 188.970 13.305 189.285 ;
        RECT 13.860 189.270 14.180 189.330 ;
        RECT 20.755 189.285 21.405 189.330 ;
        RECT 24.055 189.285 24.645 189.330 ;
        RECT 24.055 189.190 24.345 189.285 ;
        RECT 15.715 189.130 16.005 189.175 ;
        RECT 16.620 189.130 16.940 189.190 ;
        RECT 15.715 188.990 16.940 189.130 ;
        RECT 15.715 188.945 16.005 188.990 ;
        RECT 16.620 188.930 16.940 188.990 ;
        RECT 17.560 189.130 17.850 189.175 ;
        RECT 19.395 189.130 19.685 189.175 ;
        RECT 22.975 189.130 23.265 189.175 ;
        RECT 17.560 188.990 23.265 189.130 ;
        RECT 17.560 188.945 17.850 188.990 ;
        RECT 19.395 188.945 19.685 188.990 ;
        RECT 22.975 188.945 23.265 188.990 ;
        RECT 23.980 188.970 24.345 189.190 ;
        RECT 23.980 188.930 24.300 188.970 ;
        RECT 6.055 188.790 6.345 188.835 ;
        RECT 13.400 188.790 13.720 188.850 ;
        RECT 17.095 188.790 17.385 188.835 ;
        RECT 18.475 188.790 18.765 188.835 ;
        RECT 4.750 188.650 17.385 188.790 ;
        RECT 4.750 188.170 4.890 188.650 ;
        RECT 6.055 188.605 6.345 188.650 ;
        RECT 13.400 188.590 13.720 188.650 ;
        RECT 17.095 188.605 17.385 188.650 ;
        RECT 17.630 188.650 18.765 188.790 ;
        RECT 6.925 188.450 7.215 188.495 ;
        RECT 8.815 188.450 9.105 188.495 ;
        RECT 11.935 188.450 12.225 188.495 ;
        RECT 6.925 188.310 12.225 188.450 ;
        RECT 6.925 188.265 7.215 188.310 ;
        RECT 8.815 188.265 9.105 188.310 ;
        RECT 11.935 188.265 12.225 188.310 ;
        RECT 16.635 188.450 16.925 188.495 ;
        RECT 17.630 188.450 17.770 188.650 ;
        RECT 18.475 188.605 18.765 188.650 ;
        RECT 18.920 188.790 19.240 188.850 ;
        RECT 20.300 188.790 20.620 188.850 ;
        RECT 18.920 188.650 25.590 188.790 ;
        RECT 18.920 188.590 19.240 188.650 ;
        RECT 20.300 188.590 20.620 188.650 ;
        RECT 16.635 188.310 17.770 188.450 ;
        RECT 17.965 188.450 18.255 188.495 ;
        RECT 19.855 188.450 20.145 188.495 ;
        RECT 22.975 188.450 23.265 188.495 ;
        RECT 17.965 188.310 23.265 188.450 ;
        RECT 16.635 188.265 16.925 188.310 ;
        RECT 17.965 188.265 18.255 188.310 ;
        RECT 19.855 188.265 20.145 188.310 ;
        RECT 22.975 188.265 23.265 188.310 ;
        RECT 4.660 187.910 4.980 188.170 ;
        RECT 14.320 188.110 14.640 188.170 ;
        RECT 14.795 188.110 15.085 188.155 ;
        RECT 24.900 188.110 25.220 188.170 ;
        RECT 14.320 187.970 25.220 188.110 ;
        RECT 25.450 188.110 25.590 188.650 ;
        RECT 30.510 188.450 30.650 189.610 ;
        RECT 30.970 189.470 31.110 189.610 ;
        RECT 36.490 189.515 36.630 189.670 ;
        RECT 46.520 189.610 46.840 189.670 ;
        RECT 46.980 189.610 47.300 189.870 ;
        RECT 47.440 189.610 47.760 189.870 ;
        RECT 47.900 189.810 48.220 189.870 ;
        RECT 55.260 189.810 55.580 189.870 ;
        RECT 47.900 189.670 55.580 189.810 ;
        RECT 47.900 189.610 48.220 189.670 ;
        RECT 55.260 189.610 55.580 189.670 ;
        RECT 58.480 189.810 58.800 189.870 ;
        RECT 59.875 189.810 60.165 189.855 ;
        RECT 58.480 189.670 60.165 189.810 ;
        RECT 58.480 189.610 58.800 189.670 ;
        RECT 59.875 189.625 60.165 189.670 ;
        RECT 62.620 189.610 62.940 189.870 ;
        RECT 63.540 189.610 63.860 189.870 ;
        RECT 68.155 189.810 68.445 189.855 ;
        RECT 70.900 189.810 71.220 189.870 ;
        RECT 68.155 189.670 71.220 189.810 ;
        RECT 68.155 189.625 68.445 189.670 ;
        RECT 70.900 189.610 71.220 189.670 ;
        RECT 71.820 189.810 72.140 189.870 ;
        RECT 76.435 189.810 76.725 189.855 ;
        RECT 81.480 189.810 81.800 189.870 ;
        RECT 71.820 189.670 81.800 189.810 ;
        RECT 71.820 189.610 72.140 189.670 ;
        RECT 76.435 189.625 76.725 189.670 ;
        RECT 81.480 189.610 81.800 189.670 ;
        RECT 82.400 189.810 82.720 189.870 ;
        RECT 86.095 189.810 86.385 189.855 ;
        RECT 87.460 189.810 87.780 189.870 ;
        RECT 82.400 189.670 87.780 189.810 ;
        RECT 82.400 189.610 82.720 189.670 ;
        RECT 86.095 189.625 86.385 189.670 ;
        RECT 87.460 189.610 87.780 189.670 ;
        RECT 87.920 189.810 88.240 189.870 ;
        RECT 91.155 189.810 91.445 189.855 ;
        RECT 87.920 189.670 91.445 189.810 ;
        RECT 87.920 189.610 88.240 189.670 ;
        RECT 91.155 189.625 91.445 189.670 ;
        RECT 91.600 189.610 91.920 189.870 ;
        RECT 92.520 189.610 92.840 189.870 ;
        RECT 93.915 189.810 94.205 189.855 ;
        RECT 94.820 189.810 95.140 189.870 ;
        RECT 97.120 189.810 97.440 189.870 ;
        RECT 112.760 189.810 113.080 189.870 ;
        RECT 93.915 189.670 95.140 189.810 ;
        RECT 93.915 189.625 94.205 189.670 ;
        RECT 94.820 189.610 95.140 189.670 ;
        RECT 95.830 189.670 113.080 189.810 ;
        RECT 36.415 189.470 36.705 189.515 ;
        RECT 30.970 189.330 36.705 189.470 ;
        RECT 36.415 189.285 36.705 189.330 ;
        RECT 39.620 189.470 39.940 189.530 ;
        RECT 47.070 189.470 47.210 189.610 ;
        RECT 39.620 189.330 47.210 189.470 ;
        RECT 47.530 189.470 47.670 189.610 ;
        RECT 49.740 189.470 50.060 189.530 ;
        RECT 54.340 189.470 54.660 189.530 ;
        RECT 47.530 189.330 49.510 189.470 ;
        RECT 39.620 189.270 39.940 189.330 ;
        RECT 32.275 188.945 32.565 189.175 ;
        RECT 33.195 189.130 33.485 189.175 ;
        RECT 33.640 189.130 33.960 189.190 ;
        RECT 33.195 188.990 33.960 189.130 ;
        RECT 33.195 188.945 33.485 188.990 ;
        RECT 32.350 188.790 32.490 188.945 ;
        RECT 33.640 188.930 33.960 188.990 ;
        RECT 34.100 188.930 34.420 189.190 ;
        RECT 34.575 189.130 34.865 189.175 ;
        RECT 35.020 189.130 35.340 189.190 ;
        RECT 34.575 188.990 35.340 189.130 ;
        RECT 34.575 188.945 34.865 188.990 ;
        RECT 35.020 188.930 35.340 188.990 ;
        RECT 40.080 188.930 40.400 189.190 ;
        RECT 42.380 189.130 42.700 189.190 ;
        RECT 45.155 189.130 45.445 189.175 ;
        RECT 42.380 188.990 45.445 189.130 ;
        RECT 42.380 188.930 42.700 188.990 ;
        RECT 45.155 188.945 45.445 188.990 ;
        RECT 45.600 189.130 45.920 189.190 ;
        RECT 49.370 189.175 49.510 189.330 ;
        RECT 49.740 189.330 54.660 189.470 ;
        RECT 49.740 189.270 50.060 189.330 ;
        RECT 54.340 189.270 54.660 189.330 ;
        RECT 58.940 189.470 59.260 189.530 ;
        RECT 61.095 189.470 61.385 189.515 ;
        RECT 58.940 189.330 61.385 189.470 ;
        RECT 58.940 189.270 59.260 189.330 ;
        RECT 61.095 189.285 61.385 189.330 ;
        RECT 62.175 189.285 62.465 189.515 ;
        RECT 63.630 189.470 63.770 189.610 ;
        RECT 81.020 189.470 81.340 189.530 ;
        RECT 84.255 189.470 84.545 189.515 ;
        RECT 84.700 189.470 85.020 189.530 ;
        RECT 63.630 189.330 64.230 189.470 ;
        RECT 46.535 189.130 46.825 189.175 ;
        RECT 48.375 189.130 48.665 189.175 ;
        RECT 45.600 188.990 46.825 189.130 ;
        RECT 45.600 188.930 45.920 188.990 ;
        RECT 46.535 188.945 46.825 188.990 ;
        RECT 47.070 188.990 48.665 189.130 ;
        RECT 34.190 188.790 34.330 188.930 ;
        RECT 32.350 188.650 34.330 188.790 ;
        RECT 40.170 188.790 40.310 188.930 ;
        RECT 40.170 188.650 46.750 188.790 ;
        RECT 46.610 188.510 46.750 188.650 ;
        RECT 47.070 188.510 47.210 188.990 ;
        RECT 48.375 188.945 48.665 188.990 ;
        RECT 49.295 188.945 49.585 189.175 ;
        RECT 54.815 189.130 55.105 189.175 ;
        RECT 49.830 188.990 55.105 189.130 ;
        RECT 47.455 188.605 47.745 188.835 ;
        RECT 47.915 188.790 48.205 188.835 ;
        RECT 48.820 188.790 49.140 188.850 ;
        RECT 47.915 188.650 49.140 188.790 ;
        RECT 47.915 188.605 48.205 188.650 ;
        RECT 45.615 188.450 45.905 188.495 ;
        RECT 30.510 188.310 45.905 188.450 ;
        RECT 45.615 188.265 45.905 188.310 ;
        RECT 46.520 188.250 46.840 188.510 ;
        RECT 46.980 188.250 47.300 188.510 ;
        RECT 47.530 188.450 47.670 188.605 ;
        RECT 48.820 188.590 49.140 188.650 ;
        RECT 49.280 188.450 49.600 188.510 ;
        RECT 47.530 188.310 49.600 188.450 ;
        RECT 49.280 188.250 49.600 188.310 ;
        RECT 34.115 188.110 34.405 188.155 ;
        RECT 25.450 187.970 34.405 188.110 ;
        RECT 14.320 187.910 14.640 187.970 ;
        RECT 14.795 187.925 15.085 187.970 ;
        RECT 24.900 187.910 25.220 187.970 ;
        RECT 34.115 187.925 34.405 187.970 ;
        RECT 43.300 188.110 43.620 188.170 ;
        RECT 49.830 188.110 49.970 188.990 ;
        RECT 54.815 188.945 55.105 188.990 ;
        RECT 55.720 188.930 56.040 189.190 ;
        RECT 58.020 189.130 58.340 189.190 ;
        RECT 62.250 189.130 62.390 189.285 ;
        RECT 63.540 189.130 63.860 189.190 ;
        RECT 64.090 189.175 64.230 189.330 ;
        RECT 76.970 189.330 83.550 189.470 ;
        RECT 58.020 188.990 62.390 189.130 ;
        RECT 63.360 188.990 63.860 189.130 ;
        RECT 58.020 188.930 58.340 188.990 ;
        RECT 63.540 188.930 63.860 188.990 ;
        RECT 64.015 188.945 64.305 189.175 ;
        RECT 65.840 188.930 66.160 189.190 ;
        RECT 66.760 188.930 67.080 189.190 ;
        RECT 70.900 188.930 71.220 189.190 ;
        RECT 73.200 189.130 73.520 189.190 ;
        RECT 73.675 189.130 73.965 189.175 ;
        RECT 73.200 188.990 73.965 189.130 ;
        RECT 73.200 188.930 73.520 188.990 ;
        RECT 73.675 188.945 73.965 188.990 ;
        RECT 74.120 189.130 74.440 189.190 ;
        RECT 76.970 189.175 77.110 189.330 ;
        RECT 81.020 189.270 81.340 189.330 ;
        RECT 74.595 189.130 74.885 189.175 ;
        RECT 74.120 188.990 74.885 189.130 ;
        RECT 74.120 188.930 74.440 188.990 ;
        RECT 74.595 188.945 74.885 188.990 ;
        RECT 76.895 188.945 77.185 189.175 ;
        RECT 77.815 189.130 78.105 189.175 ;
        RECT 80.100 189.130 80.420 189.190 ;
        RECT 77.815 188.990 80.420 189.130 ;
        RECT 77.815 188.945 78.105 188.990 ;
        RECT 80.100 188.930 80.420 188.990 ;
        RECT 81.495 188.945 81.785 189.175 ;
        RECT 51.120 188.590 51.440 188.850 ;
        RECT 53.880 188.790 54.200 188.850 ;
        RECT 56.655 188.790 56.945 188.835 ;
        RECT 53.880 188.650 56.945 188.790 ;
        RECT 53.880 188.590 54.200 188.650 ;
        RECT 56.655 188.605 56.945 188.650 ;
        RECT 52.500 188.450 52.820 188.510 ;
        RECT 54.815 188.450 55.105 188.495 ;
        RECT 52.500 188.310 55.105 188.450 ;
        RECT 52.500 188.250 52.820 188.310 ;
        RECT 54.815 188.265 55.105 188.310 ;
        RECT 55.260 188.250 55.580 188.510 ;
        RECT 56.730 188.450 56.870 188.605 ;
        RECT 57.560 188.590 57.880 188.850 ;
        RECT 80.575 188.790 80.865 188.835 ;
        RECT 65.470 188.650 80.865 188.790 ;
        RECT 81.570 188.790 81.710 188.945 ;
        RECT 82.400 188.930 82.720 189.190 ;
        RECT 82.860 188.930 83.180 189.190 ;
        RECT 83.410 189.130 83.550 189.330 ;
        RECT 84.255 189.330 85.020 189.470 ;
        RECT 84.255 189.285 84.545 189.330 ;
        RECT 84.700 189.270 85.020 189.330 ;
        RECT 85.335 189.470 85.625 189.515 ;
        RECT 87.000 189.470 87.320 189.530 ;
        RECT 92.610 189.470 92.750 189.610 ;
        RECT 94.360 189.470 94.680 189.530 ;
        RECT 85.335 189.330 87.320 189.470 ;
        RECT 85.335 189.285 85.625 189.330 ;
        RECT 87.000 189.270 87.320 189.330 ;
        RECT 89.390 189.330 92.750 189.470 ;
        RECT 93.990 189.330 94.680 189.470 ;
        RECT 95.830 189.470 95.970 189.670 ;
        RECT 97.120 189.610 97.440 189.670 ;
        RECT 112.760 189.610 113.080 189.670 ;
        RECT 115.980 189.610 116.300 189.870 ;
        RECT 116.900 189.810 117.220 189.870 ;
        RECT 120.120 189.810 120.440 189.870 ;
        RECT 121.500 189.810 121.820 189.870 ;
        RECT 116.900 189.670 120.440 189.810 ;
        RECT 116.900 189.610 117.220 189.670 ;
        RECT 120.120 189.610 120.440 189.670 ;
        RECT 120.670 189.670 121.820 189.810 ;
        RECT 98.500 189.470 98.820 189.530 ;
        RECT 107.700 189.470 108.020 189.530 ;
        RECT 114.155 189.470 114.445 189.515 ;
        RECT 95.830 189.330 96.350 189.470 ;
        RECT 83.795 189.130 84.085 189.175 ;
        RECT 89.390 189.130 89.530 189.330 ;
        RECT 92.535 189.130 92.825 189.175 ;
        RECT 93.990 189.130 94.130 189.330 ;
        RECT 94.360 189.270 94.680 189.330 ;
        RECT 96.210 189.175 96.350 189.330 ;
        RECT 98.500 189.330 108.020 189.470 ;
        RECT 98.500 189.270 98.820 189.330 ;
        RECT 107.700 189.270 108.020 189.330 ;
        RECT 108.250 189.330 114.445 189.470 ;
        RECT 83.410 188.990 89.530 189.130 ;
        RECT 89.850 188.990 94.130 189.130 ;
        RECT 83.795 188.945 84.085 188.990 ;
        RECT 89.850 188.790 89.990 188.990 ;
        RECT 92.535 188.945 92.825 188.990 ;
        RECT 95.295 188.945 95.585 189.175 ;
        RECT 95.755 188.945 96.045 189.175 ;
        RECT 96.210 188.990 96.530 189.175 ;
        RECT 96.240 188.945 96.530 188.990 ;
        RECT 97.135 189.120 97.425 189.175 ;
        RECT 97.580 189.120 97.900 189.190 ;
        RECT 97.135 188.980 97.900 189.120 ;
        RECT 97.135 188.945 97.425 188.980 ;
        RECT 81.570 188.650 89.990 188.790 ;
        RECT 90.220 188.790 90.540 188.850 ;
        RECT 92.980 188.835 93.300 188.850 ;
        RECT 90.695 188.790 90.985 188.835 ;
        RECT 90.220 188.650 90.985 188.790 ;
        RECT 59.400 188.450 59.720 188.510 ;
        RECT 56.730 188.310 59.720 188.450 ;
        RECT 59.400 188.250 59.720 188.310 ;
        RECT 59.860 188.450 60.180 188.510 ;
        RECT 59.860 188.310 61.470 188.450 ;
        RECT 59.860 188.250 60.180 188.310 ;
        RECT 43.300 187.970 49.970 188.110 ;
        RECT 53.420 188.110 53.740 188.170 ;
        RECT 53.895 188.110 54.185 188.155 ;
        RECT 53.420 187.970 54.185 188.110 ;
        RECT 55.350 188.110 55.490 188.250 ;
        RECT 61.330 188.155 61.470 188.310 ;
        RECT 60.335 188.110 60.625 188.155 ;
        RECT 55.350 187.970 60.625 188.110 ;
        RECT 43.300 187.910 43.620 187.970 ;
        RECT 53.420 187.910 53.740 187.970 ;
        RECT 53.895 187.925 54.185 187.970 ;
        RECT 60.335 187.925 60.625 187.970 ;
        RECT 61.255 188.110 61.545 188.155 ;
        RECT 64.920 188.110 65.240 188.170 ;
        RECT 65.470 188.155 65.610 188.650 ;
        RECT 80.575 188.605 80.865 188.650 ;
        RECT 83.870 188.510 84.010 188.650 ;
        RECT 90.220 188.590 90.540 188.650 ;
        RECT 90.695 188.605 90.985 188.650 ;
        RECT 92.975 188.790 93.300 188.835 ;
        RECT 92.975 188.650 93.475 188.790 ;
        RECT 92.975 188.605 93.300 188.650 ;
        RECT 81.955 188.265 82.245 188.495 ;
        RECT 61.255 187.970 65.240 188.110 ;
        RECT 61.255 187.925 61.545 187.970 ;
        RECT 64.920 187.910 65.240 187.970 ;
        RECT 65.395 187.925 65.685 188.155 ;
        RECT 71.820 187.910 72.140 188.170 ;
        RECT 75.515 188.110 75.805 188.155 ;
        RECT 78.720 188.110 79.040 188.170 ;
        RECT 75.515 187.970 79.040 188.110 ;
        RECT 82.030 188.110 82.170 188.265 ;
        RECT 83.780 188.250 84.100 188.510 ;
        RECT 88.840 188.450 89.160 188.510 ;
        RECT 84.840 188.310 89.160 188.450 ;
        RECT 90.770 188.450 90.910 188.605 ;
        RECT 92.980 188.590 93.300 188.605 ;
        RECT 94.820 188.590 95.140 188.850 ;
        RECT 95.370 188.450 95.510 188.945 ;
        RECT 90.770 188.310 95.510 188.450 ;
        RECT 95.830 188.450 95.970 188.945 ;
        RECT 97.580 188.930 97.900 188.980 ;
        RECT 98.055 188.945 98.345 189.175 ;
        RECT 103.100 189.130 103.420 189.190 ;
        RECT 103.575 189.130 103.865 189.175 ;
        RECT 103.100 188.990 103.865 189.130 ;
        RECT 98.135 188.790 98.275 188.945 ;
        RECT 103.100 188.930 103.420 188.990 ;
        RECT 103.575 188.945 103.865 188.990 ;
        RECT 104.940 188.930 105.260 189.190 ;
        RECT 106.780 188.930 107.100 189.190 ;
        RECT 107.240 189.130 107.560 189.190 ;
        RECT 108.250 189.130 108.390 189.330 ;
        RECT 114.155 189.285 114.445 189.330 ;
        RECT 115.060 189.470 115.380 189.530 ;
        RECT 116.070 189.470 116.210 189.610 ;
        RECT 118.740 189.470 119.060 189.530 ;
        RECT 120.670 189.515 120.810 189.670 ;
        RECT 121.500 189.610 121.820 189.670 ;
        RECT 122.435 189.810 122.725 189.855 ;
        RECT 123.340 189.810 123.660 189.870 ;
        RECT 122.435 189.670 123.660 189.810 ;
        RECT 122.435 189.625 122.725 189.670 ;
        RECT 123.340 189.610 123.660 189.670 ;
        RECT 124.260 189.810 124.580 189.870 ;
        RECT 124.735 189.810 125.025 189.855 ;
        RECT 124.260 189.670 125.025 189.810 ;
        RECT 124.260 189.610 124.580 189.670 ;
        RECT 124.735 189.625 125.025 189.670 ;
        RECT 130.700 189.810 131.020 189.870 ;
        RECT 137.600 189.810 137.920 189.870 ;
        RECT 139.915 189.810 140.205 189.855 ;
        RECT 130.700 189.670 135.990 189.810 ;
        RECT 130.700 189.610 131.020 189.670 ;
        RECT 120.595 189.470 120.885 189.515 ;
        RECT 115.060 189.330 118.510 189.470 ;
        RECT 115.060 189.270 115.380 189.330 ;
        RECT 107.240 188.990 108.390 189.130 ;
        RECT 107.240 188.930 107.560 188.990 ;
        RECT 110.920 188.930 111.240 189.190 ;
        RECT 113.680 188.930 114.000 189.190 ;
        RECT 114.615 189.130 114.905 189.175 ;
        RECT 115.980 189.130 116.300 189.190 ;
        RECT 114.230 188.990 116.300 189.130 ;
        RECT 118.370 189.130 118.510 189.330 ;
        RECT 118.740 189.330 120.885 189.470 ;
        RECT 118.740 189.270 119.060 189.330 ;
        RECT 120.595 189.285 120.885 189.330 ;
        RECT 121.040 189.470 121.360 189.530 ;
        RECT 126.115 189.470 126.405 189.515 ;
        RECT 121.040 189.330 125.410 189.470 ;
        RECT 121.040 189.270 121.360 189.330 ;
        RECT 125.270 189.190 125.410 189.330 ;
        RECT 125.730 189.330 126.405 189.470 ;
        RECT 119.215 189.130 119.505 189.175 ;
        RECT 118.370 188.990 119.505 189.130 ;
        RECT 102.180 188.790 102.500 188.850 ;
        RECT 98.135 188.650 102.500 188.790 ;
        RECT 102.180 188.590 102.500 188.650 ;
        RECT 102.640 188.790 102.960 188.850 ;
        RECT 106.870 188.790 107.010 188.930 ;
        RECT 102.640 188.650 107.010 188.790 ;
        RECT 102.640 188.590 102.960 188.650 ;
        RECT 97.595 188.450 97.885 188.495 ;
        RECT 104.020 188.450 104.340 188.510 ;
        RECT 104.495 188.450 104.785 188.495 ;
        RECT 107.330 188.450 107.470 188.930 ;
        RECT 111.395 188.605 111.685 188.835 ;
        RECT 95.830 188.310 97.885 188.450 ;
        RECT 84.840 188.110 84.980 188.310 ;
        RECT 88.840 188.250 89.160 188.310 ;
        RECT 82.030 187.970 84.980 188.110 ;
        RECT 85.175 188.110 85.465 188.155 ;
        RECT 87.920 188.110 88.240 188.170 ;
        RECT 89.300 188.110 89.620 188.170 ;
        RECT 85.175 187.970 89.620 188.110 ;
        RECT 75.515 187.925 75.805 187.970 ;
        RECT 78.720 187.910 79.040 187.970 ;
        RECT 85.175 187.925 85.465 187.970 ;
        RECT 87.920 187.910 88.240 187.970 ;
        RECT 89.300 187.910 89.620 187.970 ;
        RECT 91.600 188.110 91.920 188.170 ;
        RECT 95.830 188.110 95.970 188.310 ;
        RECT 97.595 188.265 97.885 188.310 ;
        RECT 98.130 188.310 104.785 188.450 ;
        RECT 91.600 187.970 95.970 188.110 ;
        RECT 96.200 188.110 96.520 188.170 ;
        RECT 98.130 188.110 98.270 188.310 ;
        RECT 104.020 188.250 104.340 188.310 ;
        RECT 104.495 188.265 104.785 188.310 ;
        RECT 105.030 188.310 107.470 188.450 ;
        RECT 111.470 188.450 111.610 188.605 ;
        RECT 114.230 188.450 114.370 188.990 ;
        RECT 114.615 188.945 114.905 188.990 ;
        RECT 115.980 188.930 116.300 188.990 ;
        RECT 119.215 188.945 119.505 188.990 ;
        RECT 119.660 189.130 119.980 189.190 ;
        RECT 121.960 189.175 122.280 189.190 ;
        RECT 119.660 188.990 120.175 189.130 ;
        RECT 119.660 188.930 119.980 188.990 ;
        RECT 121.745 188.945 122.280 189.175 ;
        RECT 121.960 188.930 122.280 188.945 ;
        RECT 125.180 188.930 125.500 189.190 ;
        RECT 117.360 188.790 117.680 188.850 ;
        RECT 119.750 188.790 119.890 188.930 ;
        RECT 125.730 188.790 125.870 189.330 ;
        RECT 126.115 189.285 126.405 189.330 ;
        RECT 128.415 189.470 128.705 189.515 ;
        RECT 132.080 189.470 132.400 189.530 ;
        RECT 128.415 189.330 132.400 189.470 ;
        RECT 128.415 189.285 128.705 189.330 ;
        RECT 127.040 189.055 127.330 189.285 ;
        RECT 132.080 189.270 132.400 189.330 ;
        RECT 127.110 188.990 127.255 189.055 ;
        RECT 127.110 188.850 127.250 188.990 ;
        RECT 128.875 188.945 129.165 189.175 ;
        RECT 129.335 188.945 129.625 189.175 ;
        RECT 130.255 188.945 130.545 189.175 ;
        RECT 126.100 188.790 126.420 188.850 ;
        RECT 117.360 188.650 119.890 188.790 ;
        RECT 121.130 188.650 126.420 188.790 ;
        RECT 117.360 188.590 117.680 188.650 ;
        RECT 121.130 188.510 121.270 188.650 ;
        RECT 126.100 188.590 126.420 188.650 ;
        RECT 127.020 188.590 127.340 188.850 ;
        RECT 128.400 188.590 128.720 188.850 ;
        RECT 111.470 188.310 114.370 188.450 ;
        RECT 96.200 187.970 98.270 188.110 ;
        RECT 100.340 188.110 100.660 188.170 ;
        RECT 105.030 188.110 105.170 188.310 ;
        RECT 121.040 188.250 121.360 188.510 ;
        RECT 122.880 188.250 123.200 188.510 ;
        RECT 123.340 188.450 123.660 188.510 ;
        RECT 128.950 188.450 129.090 188.945 ;
        RECT 123.340 188.310 129.090 188.450 ;
        RECT 123.340 188.250 123.660 188.310 ;
        RECT 100.340 187.970 105.170 188.110 ;
        RECT 111.855 188.110 112.145 188.155 ;
        RECT 112.760 188.110 113.080 188.170 ;
        RECT 111.855 187.970 113.080 188.110 ;
        RECT 91.600 187.910 91.920 187.970 ;
        RECT 96.200 187.910 96.520 187.970 ;
        RECT 100.340 187.910 100.660 187.970 ;
        RECT 111.855 187.925 112.145 187.970 ;
        RECT 112.760 187.910 113.080 187.970 ;
        RECT 117.820 188.110 118.140 188.170 ;
        RECT 122.970 188.110 123.110 188.250 ;
        RECT 117.820 187.970 123.110 188.110 ;
        RECT 126.560 188.110 126.880 188.170 ;
        RECT 127.495 188.110 127.785 188.155 ;
        RECT 126.560 187.970 127.785 188.110 ;
        RECT 129.410 188.110 129.550 188.945 ;
        RECT 130.330 188.510 130.470 188.945 ;
        RECT 130.700 188.930 131.020 189.190 ;
        RECT 131.175 189.130 131.465 189.175 ;
        RECT 133.015 189.130 133.305 189.175 ;
        RECT 131.175 188.990 133.305 189.130 ;
        RECT 131.175 188.945 131.465 188.990 ;
        RECT 133.015 188.945 133.305 188.990 ;
        RECT 133.920 188.930 134.240 189.190 ;
        RECT 135.850 189.175 135.990 189.670 ;
        RECT 137.600 189.670 140.205 189.810 ;
        RECT 137.600 189.610 137.920 189.670 ;
        RECT 139.915 189.625 140.205 189.670 ;
        RECT 147.720 189.810 148.040 189.870 ;
        RECT 149.575 189.810 149.865 189.855 ;
        RECT 147.720 189.670 149.865 189.810 ;
        RECT 147.720 189.610 148.040 189.670 ;
        RECT 149.575 189.625 149.865 189.670 ;
        RECT 136.695 189.470 136.985 189.515 ;
        RECT 138.075 189.470 138.365 189.515 ;
        RECT 136.695 189.330 138.365 189.470 ;
        RECT 136.695 189.285 136.985 189.330 ;
        RECT 138.075 189.285 138.365 189.330 ;
        RECT 138.520 189.270 138.840 189.530 ;
        RECT 140.835 189.470 141.125 189.515 ;
        RECT 147.810 189.470 147.950 189.610 ;
        RECT 140.835 189.330 143.350 189.470 ;
        RECT 140.835 189.285 141.125 189.330 ;
        RECT 143.210 189.190 143.350 189.330 ;
        RECT 146.430 189.330 147.950 189.470 ;
        RECT 135.775 188.945 136.065 189.175 ;
        RECT 137.140 188.930 137.460 189.190 ;
        RECT 137.600 189.130 137.920 189.190 ;
        RECT 138.995 189.130 139.285 189.175 ;
        RECT 137.600 188.990 139.285 189.130 ;
        RECT 137.600 188.930 137.920 188.990 ;
        RECT 138.995 188.945 139.285 188.990 ;
        RECT 139.900 189.130 140.220 189.190 ;
        RECT 140.375 189.130 140.665 189.175 ;
        RECT 139.900 188.990 140.665 189.130 ;
        RECT 139.900 188.930 140.220 188.990 ;
        RECT 140.375 188.945 140.665 188.990 ;
        RECT 141.280 189.130 141.600 189.190 ;
        RECT 141.755 189.130 142.045 189.175 ;
        RECT 141.280 188.990 142.045 189.130 ;
        RECT 141.280 188.930 141.600 188.990 ;
        RECT 141.755 188.945 142.045 188.990 ;
        RECT 143.120 188.930 143.440 189.190 ;
        RECT 146.430 189.175 146.570 189.330 ;
        RECT 151.860 189.270 152.180 189.530 ;
        RECT 146.355 188.945 146.645 189.175 ;
        RECT 146.800 188.930 147.120 189.190 ;
        RECT 147.275 188.945 147.565 189.175 ;
        RECT 130.790 188.790 130.930 188.930 ;
        RECT 134.395 188.790 134.685 188.835 ;
        RECT 130.790 188.650 134.685 188.790 ;
        RECT 134.395 188.605 134.685 188.650 ;
        RECT 134.855 188.790 135.145 188.835 ;
        RECT 144.975 188.790 145.265 188.835 ;
        RECT 134.855 188.650 145.265 188.790 ;
        RECT 147.350 188.790 147.490 188.945 ;
        RECT 148.180 188.930 148.500 189.190 ;
        RECT 148.640 189.130 148.960 189.190 ;
        RECT 150.495 189.130 150.785 189.175 ;
        RECT 148.640 188.990 150.785 189.130 ;
        RECT 148.640 188.930 148.960 188.990 ;
        RECT 150.495 188.945 150.785 188.990 ;
        RECT 150.940 188.930 151.260 189.190 ;
        RECT 151.415 189.130 151.705 189.175 ;
        RECT 151.950 189.130 152.090 189.270 ;
        RECT 152.780 189.130 153.100 189.190 ;
        RECT 151.415 188.990 153.100 189.130 ;
        RECT 151.415 188.945 151.705 188.990 ;
        RECT 152.780 188.930 153.100 188.990 ;
        RECT 149.100 188.790 149.420 188.850 ;
        RECT 147.350 188.650 149.420 188.790 ;
        RECT 134.855 188.605 135.145 188.650 ;
        RECT 144.975 188.605 145.265 188.650 ;
        RECT 149.100 188.590 149.420 188.650 ;
        RECT 151.860 188.590 152.180 188.850 ;
        RECT 130.240 188.250 130.560 188.510 ;
        RECT 142.660 188.110 142.980 188.170 ;
        RECT 129.410 187.970 142.980 188.110 ;
        RECT 117.820 187.910 118.140 187.970 ;
        RECT 126.560 187.910 126.880 187.970 ;
        RECT 127.495 187.925 127.785 187.970 ;
        RECT 142.660 187.910 142.980 187.970 ;
        RECT 2.750 187.290 158.230 187.770 ;
        RECT 16.635 187.090 16.925 187.135 ;
        RECT 17.080 187.090 17.400 187.150 ;
        RECT 16.635 186.950 17.400 187.090 ;
        RECT 16.635 186.905 16.925 186.950 ;
        RECT 17.080 186.890 17.400 186.950 ;
        RECT 18.460 186.890 18.780 187.150 ;
        RECT 27.660 187.090 27.980 187.150 ;
        RECT 33.195 187.090 33.485 187.135 ;
        RECT 27.660 186.950 33.485 187.090 ;
        RECT 27.660 186.890 27.980 186.950 ;
        RECT 33.195 186.905 33.485 186.950 ;
        RECT 41.935 187.090 42.225 187.135 ;
        RECT 44.220 187.090 44.540 187.150 ;
        RECT 41.935 186.950 44.540 187.090 ;
        RECT 41.935 186.905 42.225 186.950 ;
        RECT 44.220 186.890 44.540 186.950 ;
        RECT 51.120 186.890 51.440 187.150 ;
        RECT 59.400 187.090 59.720 187.150 ;
        RECT 80.575 187.090 80.865 187.135 ;
        RECT 81.020 187.090 81.340 187.150 ;
        RECT 52.130 186.950 59.170 187.090 ;
        RECT 4.680 186.750 4.970 186.795 ;
        RECT 6.540 186.750 6.830 186.795 ;
        RECT 9.320 186.750 9.610 186.795 ;
        RECT 15.700 186.750 16.020 186.810 ;
        RECT 18.550 186.750 18.690 186.890 ;
        RECT 23.485 186.750 23.775 186.795 ;
        RECT 25.375 186.750 25.665 186.795 ;
        RECT 28.495 186.750 28.785 186.795 ;
        RECT 4.680 186.610 9.610 186.750 ;
        RECT 4.680 186.565 4.970 186.610 ;
        RECT 6.540 186.565 6.830 186.610 ;
        RECT 9.320 186.565 9.610 186.610 ;
        RECT 13.030 186.610 16.020 186.750 ;
        RECT 3.740 186.410 4.060 186.470 ;
        RECT 13.030 186.410 13.170 186.610 ;
        RECT 15.700 186.550 16.020 186.610 ;
        RECT 17.250 186.610 18.230 186.750 ;
        RECT 18.550 186.610 22.830 186.750 ;
        RECT 3.740 186.270 13.170 186.410 ;
        RECT 13.400 186.410 13.720 186.470 ;
        RECT 17.250 186.410 17.390 186.610 ;
        RECT 13.400 186.270 17.390 186.410 ;
        RECT 3.740 186.210 4.060 186.270 ;
        RECT 13.400 186.210 13.720 186.270 ;
        RECT 17.540 186.210 17.860 186.470 ;
        RECT 18.090 186.410 18.230 186.610 ;
        RECT 22.690 186.455 22.830 186.610 ;
        RECT 23.485 186.610 28.785 186.750 ;
        RECT 23.485 186.565 23.775 186.610 ;
        RECT 25.375 186.565 25.665 186.610 ;
        RECT 28.495 186.565 28.785 186.610 ;
        RECT 45.600 186.750 45.920 186.810 ;
        RECT 52.130 186.750 52.270 186.950 ;
        RECT 59.030 186.810 59.170 186.950 ;
        RECT 59.400 186.950 63.310 187.090 ;
        RECT 59.400 186.890 59.720 186.950 ;
        RECT 45.600 186.610 52.270 186.750 ;
        RECT 52.465 186.750 52.755 186.795 ;
        RECT 54.355 186.750 54.645 186.795 ;
        RECT 57.475 186.750 57.765 186.795 ;
        RECT 52.465 186.610 57.765 186.750 ;
        RECT 45.600 186.550 45.920 186.610 ;
        RECT 52.465 186.565 52.755 186.610 ;
        RECT 54.355 186.565 54.645 186.610 ;
        RECT 57.475 186.565 57.765 186.610 ;
        RECT 58.940 186.550 59.260 186.810 ;
        RECT 62.160 186.550 62.480 186.810 ;
        RECT 21.235 186.410 21.525 186.455 ;
        RECT 18.090 186.270 21.525 186.410 ;
        RECT 21.235 186.225 21.525 186.270 ;
        RECT 22.615 186.225 22.905 186.455 ;
        RECT 34.100 186.410 34.420 186.470 ;
        RECT 42.840 186.410 43.160 186.470 ;
        RECT 44.235 186.410 44.525 186.455 ;
        RECT 45.155 186.410 45.445 186.455 ;
        RECT 47.900 186.410 48.220 186.470 ;
        RECT 34.100 186.270 43.160 186.410 ;
        RECT 34.100 186.210 34.420 186.270 ;
        RECT 42.840 186.210 43.160 186.270 ;
        RECT 43.390 186.270 44.525 186.410 ;
        RECT 4.215 186.070 4.505 186.115 ;
        RECT 4.660 186.070 4.980 186.130 ;
        RECT 4.215 185.930 4.980 186.070 ;
        RECT 4.215 185.885 4.505 185.930 ;
        RECT 4.660 185.870 4.980 185.930 ;
        RECT 6.040 185.870 6.360 186.130 ;
        RECT 9.320 186.070 9.610 186.115 ;
        RECT 7.075 185.930 9.610 186.070 ;
        RECT 17.630 185.995 17.770 186.210 ;
        RECT 18.000 186.070 18.320 186.130 ;
        RECT 20.775 186.070 21.065 186.115 ;
        RECT 7.075 185.775 7.290 185.930 ;
        RECT 9.320 185.885 9.610 185.930 ;
        RECT 11.100 185.775 11.420 185.790 ;
        RECT 5.140 185.730 5.430 185.775 ;
        RECT 7.000 185.730 7.290 185.775 ;
        RECT 5.140 185.590 7.290 185.730 ;
        RECT 5.140 185.545 5.430 185.590 ;
        RECT 7.000 185.545 7.290 185.590 ;
        RECT 7.920 185.730 8.210 185.775 ;
        RECT 11.100 185.730 11.470 185.775 ;
        RECT 13.860 185.730 14.180 185.790 ;
        RECT 17.555 185.765 17.845 185.995 ;
        RECT 18.000 185.930 21.065 186.070 ;
        RECT 18.000 185.870 18.320 185.930 ;
        RECT 20.775 185.885 21.065 185.930 ;
        RECT 23.080 186.070 23.370 186.115 ;
        RECT 24.915 186.070 25.205 186.115 ;
        RECT 28.495 186.070 28.785 186.115 ;
        RECT 23.080 185.930 28.785 186.070 ;
        RECT 23.080 185.885 23.370 185.930 ;
        RECT 24.915 185.885 25.205 185.930 ;
        RECT 28.495 185.885 28.785 185.930 ;
        RECT 29.575 186.070 29.865 186.090 ;
        RECT 34.560 186.070 34.880 186.130 ;
        RECT 36.860 186.070 37.180 186.130 ;
        RECT 29.575 185.930 37.180 186.070 ;
        RECT 7.920 185.590 14.180 185.730 ;
        RECT 7.920 185.545 8.210 185.590 ;
        RECT 11.100 185.545 11.470 185.590 ;
        RECT 11.100 185.530 11.420 185.545 ;
        RECT 13.860 185.530 14.180 185.590 ;
        RECT 23.980 185.530 24.300 185.790 ;
        RECT 29.575 185.775 29.865 185.930 ;
        RECT 34.560 185.870 34.880 185.930 ;
        RECT 36.860 185.870 37.180 185.930 ;
        RECT 39.620 186.070 39.940 186.130 ;
        RECT 43.390 186.070 43.530 186.270 ;
        RECT 44.235 186.225 44.525 186.270 ;
        RECT 44.770 186.270 45.445 186.410 ;
        RECT 44.770 186.130 44.910 186.270 ;
        RECT 45.155 186.225 45.445 186.270 ;
        RECT 46.150 186.270 48.220 186.410 ;
        RECT 39.620 185.930 43.530 186.070 ;
        RECT 39.620 185.870 39.940 185.930 ;
        RECT 43.760 185.870 44.080 186.130 ;
        RECT 44.680 185.870 45.000 186.130 ;
        RECT 46.150 186.115 46.290 186.270 ;
        RECT 47.900 186.210 48.220 186.270 ;
        RECT 49.740 186.410 50.060 186.470 ;
        RECT 51.595 186.410 51.885 186.455 ;
        RECT 49.740 186.270 51.885 186.410 ;
        RECT 49.740 186.210 50.060 186.270 ;
        RECT 51.595 186.225 51.885 186.270 ;
        RECT 52.975 186.410 53.265 186.455 ;
        RECT 53.420 186.410 53.740 186.470 ;
        RECT 52.975 186.270 53.740 186.410 ;
        RECT 52.975 186.225 53.265 186.270 ;
        RECT 53.420 186.210 53.740 186.270 ;
        RECT 55.260 186.410 55.580 186.470 ;
        RECT 58.020 186.410 58.340 186.470 ;
        RECT 60.335 186.410 60.625 186.455 ;
        RECT 55.260 186.270 60.625 186.410 ;
        RECT 55.260 186.210 55.580 186.270 ;
        RECT 58.020 186.210 58.340 186.270 ;
        RECT 60.335 186.225 60.625 186.270 ;
        RECT 63.170 186.410 63.310 186.950 ;
        RECT 80.575 186.950 81.340 187.090 ;
        RECT 80.575 186.905 80.865 186.950 ;
        RECT 81.020 186.890 81.340 186.950 ;
        RECT 83.335 187.090 83.625 187.135 ;
        RECT 83.780 187.090 84.100 187.150 ;
        RECT 83.335 186.950 84.100 187.090 ;
        RECT 83.335 186.905 83.625 186.950 ;
        RECT 83.780 186.890 84.100 186.950 ;
        RECT 87.920 187.090 88.240 187.150 ;
        RECT 92.060 187.090 92.380 187.150 ;
        RECT 93.915 187.090 94.205 187.135 ;
        RECT 87.920 186.950 91.370 187.090 ;
        RECT 87.920 186.890 88.240 186.950 ;
        RECT 64.000 186.750 64.320 186.810 ;
        RECT 66.760 186.750 67.080 186.810 ;
        RECT 85.160 186.750 85.480 186.810 ;
        RECT 89.300 186.750 89.620 186.810 ;
        RECT 64.000 186.610 89.620 186.750 ;
        RECT 91.230 186.750 91.370 186.950 ;
        RECT 92.060 186.950 94.205 187.090 ;
        RECT 92.060 186.890 92.380 186.950 ;
        RECT 93.915 186.905 94.205 186.950 ;
        RECT 97.580 186.890 97.900 187.150 ;
        RECT 98.515 186.905 98.805 187.135 ;
        RECT 99.435 187.090 99.725 187.135 ;
        RECT 100.800 187.090 101.120 187.150 ;
        RECT 112.760 187.090 113.080 187.150 ;
        RECT 113.235 187.090 113.525 187.135 ;
        RECT 113.680 187.090 114.000 187.150 ;
        RECT 99.435 186.950 101.120 187.090 ;
        RECT 99.435 186.905 99.725 186.950 ;
        RECT 97.670 186.750 97.810 186.890 ;
        RECT 91.230 186.610 97.810 186.750 ;
        RECT 98.590 186.750 98.730 186.905 ;
        RECT 100.800 186.890 101.120 186.950 ;
        RECT 101.350 186.950 114.000 187.090 ;
        RECT 99.880 186.750 100.200 186.810 ;
        RECT 98.590 186.610 100.200 186.750 ;
        RECT 64.000 186.550 64.320 186.610 ;
        RECT 66.760 186.550 67.080 186.610 ;
        RECT 85.160 186.550 85.480 186.610 ;
        RECT 89.300 186.550 89.620 186.610 ;
        RECT 99.880 186.550 100.200 186.610 ;
        RECT 74.135 186.410 74.425 186.455 ;
        RECT 63.170 186.270 74.425 186.410 ;
        RECT 46.075 185.885 46.365 186.115 ;
        RECT 46.520 186.070 46.840 186.130 ;
        RECT 46.995 186.070 47.285 186.115 ;
        RECT 46.520 185.930 47.285 186.070 ;
        RECT 46.520 185.870 46.840 185.930 ;
        RECT 46.995 185.885 47.285 185.930 ;
        RECT 47.440 185.870 47.760 186.130 ;
        RECT 48.375 185.885 48.665 186.115 ;
        RECT 26.275 185.730 26.925 185.775 ;
        RECT 29.575 185.730 30.165 185.775 ;
        RECT 40.080 185.730 40.400 185.790 ;
        RECT 40.555 185.730 40.845 185.775 ;
        RECT 42.380 185.730 42.700 185.790 ;
        RECT 26.275 185.590 30.165 185.730 ;
        RECT 26.275 185.545 26.925 185.590 ;
        RECT 29.875 185.545 30.165 185.590 ;
        RECT 30.510 185.590 35.710 185.730 ;
        RECT 12.940 185.435 13.260 185.450 ;
        RECT 12.940 185.205 13.475 185.435 ;
        RECT 18.000 185.390 18.320 185.450 ;
        RECT 18.475 185.390 18.765 185.435 ;
        RECT 18.000 185.250 18.765 185.390 ;
        RECT 12.940 185.190 13.260 185.205 ;
        RECT 18.000 185.190 18.320 185.250 ;
        RECT 18.475 185.205 18.765 185.250 ;
        RECT 20.300 185.190 20.620 185.450 ;
        RECT 21.220 185.390 21.540 185.450 ;
        RECT 23.060 185.390 23.380 185.450 ;
        RECT 30.510 185.390 30.650 185.590 ;
        RECT 35.570 185.450 35.710 185.590 ;
        RECT 40.080 185.590 42.700 185.730 ;
        RECT 40.080 185.530 40.400 185.590 ;
        RECT 40.555 185.545 40.845 185.590 ;
        RECT 42.380 185.530 42.700 185.590 ;
        RECT 21.220 185.250 30.650 185.390 ;
        RECT 21.220 185.190 21.540 185.250 ;
        RECT 23.060 185.190 23.380 185.250 ;
        RECT 31.340 185.190 31.660 185.450 ;
        RECT 35.480 185.390 35.800 185.450 ;
        RECT 45.140 185.390 45.460 185.450 ;
        RECT 35.480 185.250 45.460 185.390 ;
        RECT 35.480 185.190 35.800 185.250 ;
        RECT 45.140 185.190 45.460 185.250 ;
        RECT 46.520 185.190 46.840 185.450 ;
        RECT 48.450 185.390 48.590 185.885 ;
        RECT 48.820 185.870 49.140 186.130 ;
        RECT 49.280 185.870 49.600 186.130 ;
        RECT 50.200 185.870 50.520 186.130 ;
        RECT 52.060 186.070 52.350 186.115 ;
        RECT 53.895 186.070 54.185 186.115 ;
        RECT 57.475 186.070 57.765 186.115 ;
        RECT 52.060 185.930 57.765 186.070 ;
        RECT 52.060 185.885 52.350 185.930 ;
        RECT 53.895 185.885 54.185 185.930 ;
        RECT 57.475 185.885 57.765 185.930 ;
        RECT 48.910 185.730 49.050 185.870 ;
        RECT 52.960 185.730 53.280 185.790 ;
        RECT 48.910 185.590 53.280 185.730 ;
        RECT 52.960 185.530 53.280 185.590 ;
        RECT 54.340 185.730 54.660 185.790 ;
        RECT 58.555 185.775 58.845 186.090 ;
        RECT 62.160 185.870 62.480 186.130 ;
        RECT 63.170 186.070 63.310 186.270 ;
        RECT 64.015 186.070 64.305 186.115 ;
        RECT 63.170 185.930 64.305 186.070 ;
        RECT 64.015 185.885 64.305 185.930 ;
        RECT 64.920 186.070 65.240 186.130 ;
        RECT 68.690 186.115 68.830 186.270 ;
        RECT 74.135 186.225 74.425 186.270 ;
        RECT 76.420 186.410 76.740 186.470 ;
        RECT 101.350 186.410 101.490 186.950 ;
        RECT 112.760 186.890 113.080 186.950 ;
        RECT 113.235 186.905 113.525 186.950 ;
        RECT 113.680 186.890 114.000 186.950 ;
        RECT 114.140 187.090 114.460 187.150 ;
        RECT 115.060 187.090 115.380 187.150 ;
        RECT 114.140 186.950 115.380 187.090 ;
        RECT 114.140 186.890 114.460 186.950 ;
        RECT 115.060 186.890 115.380 186.950 ;
        RECT 117.360 187.090 117.680 187.150 ;
        RECT 127.955 187.090 128.245 187.135 ;
        RECT 137.600 187.090 137.920 187.150 ;
        RECT 117.360 186.950 127.710 187.090 ;
        RECT 117.360 186.890 117.680 186.950 ;
        RECT 102.180 186.750 102.500 186.810 ;
        RECT 114.615 186.750 114.905 186.795 ;
        RECT 127.020 186.750 127.340 186.810 ;
        RECT 102.180 186.610 111.150 186.750 ;
        RECT 102.180 186.550 102.500 186.610 ;
        RECT 111.010 186.470 111.150 186.610 ;
        RECT 114.615 186.610 127.340 186.750 ;
        RECT 114.615 186.565 114.905 186.610 ;
        RECT 127.020 186.550 127.340 186.610 ;
        RECT 104.480 186.410 104.800 186.470 ;
        RECT 108.620 186.410 108.940 186.470 ;
        RECT 76.420 186.270 101.490 186.410 ;
        RECT 101.810 186.270 108.940 186.410 ;
        RECT 76.420 186.210 76.740 186.270 ;
        RECT 65.855 186.070 66.145 186.115 ;
        RECT 67.695 186.070 67.985 186.115 ;
        RECT 64.920 185.930 67.985 186.070 ;
        RECT 64.920 185.870 65.240 185.930 ;
        RECT 65.855 185.885 66.145 185.930 ;
        RECT 67.695 185.885 67.985 185.930 ;
        RECT 68.615 185.885 68.905 186.115 ;
        RECT 69.995 185.885 70.285 186.115 ;
        RECT 71.360 186.070 71.680 186.130 ;
        RECT 72.755 186.070 73.045 186.115 ;
        RECT 71.360 185.930 73.045 186.070 ;
        RECT 55.255 185.730 55.905 185.775 ;
        RECT 58.555 185.730 59.145 185.775 ;
        RECT 54.340 185.590 59.145 185.730 ;
        RECT 62.250 185.730 62.390 185.870 ;
        RECT 70.070 185.730 70.210 185.885 ;
        RECT 71.360 185.870 71.680 185.930 ;
        RECT 72.755 185.885 73.045 185.930 ;
        RECT 73.215 185.885 73.505 186.115 ;
        RECT 77.355 186.070 77.645 186.115 ;
        RECT 73.750 185.930 77.645 186.070 ;
        RECT 62.250 185.590 70.210 185.730 ;
        RECT 54.340 185.530 54.660 185.590 ;
        RECT 55.255 185.545 55.905 185.590 ;
        RECT 58.855 185.545 59.145 185.590 ;
        RECT 59.400 185.390 59.720 185.450 ;
        RECT 48.450 185.250 59.720 185.390 ;
        RECT 59.400 185.190 59.720 185.250 ;
        RECT 69.520 185.390 69.840 185.450 ;
        RECT 73.290 185.390 73.430 185.885 ;
        RECT 73.750 185.450 73.890 185.930 ;
        RECT 77.355 185.885 77.645 185.930 ;
        RECT 77.430 185.730 77.570 185.885 ;
        RECT 78.260 185.870 78.580 186.130 ;
        RECT 78.720 186.070 79.040 186.130 ;
        RECT 79.195 186.070 79.485 186.115 ;
        RECT 78.720 185.930 79.485 186.070 ;
        RECT 78.720 185.870 79.040 185.930 ;
        RECT 79.195 185.885 79.485 185.930 ;
        RECT 80.100 186.070 80.420 186.130 ;
        RECT 81.480 186.070 81.800 186.130 ;
        RECT 81.955 186.070 82.245 186.115 ;
        RECT 80.100 185.930 82.245 186.070 ;
        RECT 80.100 185.870 80.420 185.930 ;
        RECT 81.480 185.870 81.800 185.930 ;
        RECT 81.955 185.885 82.245 185.930 ;
        RECT 83.780 186.070 84.100 186.130 ;
        RECT 86.080 186.070 86.400 186.130 ;
        RECT 83.780 185.930 100.570 186.070 ;
        RECT 83.780 185.870 84.100 185.930 ;
        RECT 86.080 185.870 86.400 185.930 ;
        RECT 87.000 185.730 87.320 185.790 ;
        RECT 77.430 185.590 87.320 185.730 ;
        RECT 87.000 185.530 87.320 185.590 ;
        RECT 95.295 185.545 95.585 185.775 ;
        RECT 95.740 185.730 96.060 185.790 ;
        RECT 97.595 185.730 97.885 185.775 ;
        RECT 95.740 185.590 97.885 185.730 ;
        RECT 69.520 185.250 73.430 185.390 ;
        RECT 69.520 185.190 69.840 185.250 ;
        RECT 73.660 185.190 73.980 185.450 ;
        RECT 77.340 185.390 77.660 185.450 ;
        RECT 86.080 185.390 86.400 185.450 ;
        RECT 77.340 185.250 86.400 185.390 ;
        RECT 77.340 185.190 77.660 185.250 ;
        RECT 86.080 185.190 86.400 185.250 ;
        RECT 86.540 185.390 86.860 185.450 ;
        RECT 90.220 185.390 90.540 185.450 ;
        RECT 86.540 185.250 90.540 185.390 ;
        RECT 95.370 185.390 95.510 185.545 ;
        RECT 95.740 185.530 96.060 185.590 ;
        RECT 97.595 185.545 97.885 185.590 ;
        RECT 98.040 185.730 98.360 185.790 ;
        RECT 98.040 185.590 100.110 185.730 ;
        RECT 98.040 185.530 98.360 185.590 ;
        RECT 99.970 185.450 100.110 185.590 ;
        RECT 97.120 185.390 97.440 185.450 ;
        RECT 95.370 185.250 97.440 185.390 ;
        RECT 86.540 185.190 86.860 185.250 ;
        RECT 90.220 185.190 90.540 185.250 ;
        RECT 97.120 185.190 97.440 185.250 ;
        RECT 98.645 185.390 98.935 185.435 ;
        RECT 99.420 185.390 99.740 185.450 ;
        RECT 98.645 185.250 99.740 185.390 ;
        RECT 98.645 185.205 98.935 185.250 ;
        RECT 99.420 185.190 99.740 185.250 ;
        RECT 99.880 185.190 100.200 185.450 ;
        RECT 100.430 185.390 100.570 185.930 ;
        RECT 100.800 185.870 101.120 186.130 ;
        RECT 101.810 186.115 101.950 186.270 ;
        RECT 104.480 186.210 104.800 186.270 ;
        RECT 108.620 186.210 108.940 186.270 ;
        RECT 110.920 186.210 111.240 186.470 ;
        RECT 112.775 186.410 113.065 186.455 ;
        RECT 118.740 186.410 119.060 186.470 ;
        RECT 112.775 186.270 119.060 186.410 ;
        RECT 112.775 186.225 113.065 186.270 ;
        RECT 101.735 185.885 102.025 186.115 ;
        RECT 102.195 186.070 102.485 186.115 ;
        RECT 102.195 185.930 104.710 186.070 ;
        RECT 102.195 185.885 102.485 185.930 ;
        RECT 100.890 185.730 101.030 185.870 ;
        RECT 103.100 185.730 103.420 185.790 ;
        RECT 100.890 185.590 103.420 185.730 ;
        RECT 103.100 185.530 103.420 185.590 ;
        RECT 104.570 185.450 104.710 185.930 ;
        RECT 104.940 185.870 105.260 186.130 ;
        RECT 105.415 186.070 105.705 186.115 ;
        RECT 105.860 186.070 106.180 186.130 ;
        RECT 108.160 186.070 108.480 186.130 ;
        RECT 105.415 185.930 108.480 186.070 ;
        RECT 105.415 185.885 105.705 185.930 ;
        RECT 105.860 185.870 106.180 185.930 ;
        RECT 108.160 185.870 108.480 185.930 ;
        RECT 111.840 185.870 112.160 186.130 ;
        RECT 113.235 186.070 113.525 186.115 ;
        RECT 114.140 186.070 114.460 186.130 ;
        RECT 113.235 185.930 114.460 186.070 ;
        RECT 113.235 185.885 113.525 185.930 ;
        RECT 114.140 185.870 114.460 185.930 ;
        RECT 115.060 186.070 115.380 186.130 ;
        RECT 115.535 186.070 115.825 186.115 ;
        RECT 115.060 185.930 115.825 186.070 ;
        RECT 115.060 185.870 115.380 185.930 ;
        RECT 115.535 185.885 115.825 185.930 ;
        RECT 115.995 185.885 116.285 186.115 ;
        RECT 106.320 185.530 106.640 185.790 ;
        RECT 113.680 185.730 114.000 185.790 ;
        RECT 114.600 185.730 114.920 185.790 ;
        RECT 113.680 185.590 114.920 185.730 ;
        RECT 116.070 185.730 116.210 185.885 ;
        RECT 116.440 185.870 116.760 186.130 ;
        RECT 117.450 186.115 117.590 186.270 ;
        RECT 118.740 186.210 119.060 186.270 ;
        RECT 119.660 186.410 119.980 186.470 ;
        RECT 121.055 186.410 121.345 186.455 ;
        RECT 119.660 186.270 121.345 186.410 ;
        RECT 119.660 186.210 119.980 186.270 ;
        RECT 121.055 186.225 121.345 186.270 ;
        RECT 121.500 186.410 121.820 186.470 ;
        RECT 123.815 186.410 124.105 186.455 ;
        RECT 126.115 186.410 126.405 186.455 ;
        RECT 121.500 186.270 123.110 186.410 ;
        RECT 121.500 186.210 121.820 186.270 ;
        RECT 117.375 186.070 117.665 186.115 ;
        RECT 120.120 186.070 120.440 186.130 ;
        RECT 122.970 186.115 123.110 186.270 ;
        RECT 123.815 186.270 126.405 186.410 ;
        RECT 123.815 186.225 124.105 186.270 ;
        RECT 126.115 186.225 126.405 186.270 ;
        RECT 121.975 186.070 122.265 186.115 ;
        RECT 117.375 185.930 117.775 186.070 ;
        RECT 120.120 185.930 122.265 186.070 ;
        RECT 117.375 185.885 117.665 185.930 ;
        RECT 120.120 185.870 120.440 185.930 ;
        RECT 121.130 185.790 121.270 185.930 ;
        RECT 121.975 185.885 122.265 185.930 ;
        RECT 122.895 185.885 123.185 186.115 ;
        RECT 125.640 185.870 125.960 186.130 ;
        RECT 126.560 185.870 126.880 186.130 ;
        RECT 127.110 186.115 127.250 186.550 ;
        RECT 127.570 186.410 127.710 186.950 ;
        RECT 127.955 186.950 137.920 187.090 ;
        RECT 127.955 186.905 128.245 186.950 ;
        RECT 137.600 186.890 137.920 186.950 ;
        RECT 140.820 187.090 141.140 187.150 ;
        RECT 141.295 187.090 141.585 187.135 ;
        RECT 140.820 186.950 141.585 187.090 ;
        RECT 140.820 186.890 141.140 186.950 ;
        RECT 141.295 186.905 141.585 186.950 ;
        RECT 142.215 187.090 142.505 187.135 ;
        RECT 146.800 187.090 147.120 187.150 ;
        RECT 142.215 186.950 147.120 187.090 ;
        RECT 142.215 186.905 142.505 186.950 ;
        RECT 146.800 186.890 147.120 186.950 ;
        RECT 150.940 186.890 151.260 187.150 ;
        RECT 154.160 186.890 154.480 187.150 ;
        RECT 128.400 186.750 128.720 186.810 ;
        RECT 151.030 186.750 151.170 186.890 ;
        RECT 128.400 186.610 151.170 186.750 ;
        RECT 128.400 186.550 128.720 186.610 ;
        RECT 135.760 186.410 136.080 186.470 ;
        RECT 139.900 186.410 140.220 186.470 ;
        RECT 155.540 186.410 155.860 186.470 ;
        RECT 127.570 186.270 136.080 186.410 ;
        RECT 127.035 185.885 127.325 186.115 ;
        RECT 133.000 185.870 133.320 186.130 ;
        RECT 134.010 186.115 134.150 186.270 ;
        RECT 135.760 186.210 136.080 186.270 ;
        RECT 138.150 186.270 140.220 186.410 ;
        RECT 133.935 185.885 134.225 186.115 ;
        RECT 134.380 185.870 134.700 186.130 ;
        RECT 134.840 186.070 135.160 186.130 ;
        RECT 138.150 186.070 138.290 186.270 ;
        RECT 139.900 186.210 140.220 186.270 ;
        RECT 152.410 186.270 155.860 186.410 ;
        RECT 152.410 186.070 152.550 186.270 ;
        RECT 155.540 186.210 155.860 186.270 ;
        RECT 134.840 185.930 138.290 186.070 ;
        RECT 138.610 185.930 152.550 186.070 ;
        RECT 134.840 185.870 135.160 185.930 ;
        RECT 116.915 185.730 117.205 185.775 ;
        RECT 116.070 185.590 117.205 185.730 ;
        RECT 113.680 185.530 114.000 185.590 ;
        RECT 114.600 185.530 114.920 185.590 ;
        RECT 116.915 185.545 117.205 185.590 ;
        RECT 121.040 185.530 121.360 185.790 ;
        RECT 133.090 185.730 133.230 185.870 ;
        RECT 138.610 185.730 138.750 185.930 ;
        RECT 152.780 185.870 153.100 186.130 ;
        RECT 122.050 185.590 124.950 185.730 ;
        RECT 133.090 185.590 138.750 185.730 ;
        RECT 101.720 185.390 102.040 185.450 ;
        RECT 100.430 185.250 102.040 185.390 ;
        RECT 101.720 185.190 102.040 185.250 ;
        RECT 104.480 185.190 104.800 185.450 ;
        RECT 105.840 185.390 106.130 185.435 ;
        RECT 122.050 185.390 122.190 185.590 ;
        RECT 105.840 185.250 122.190 185.390 ;
        RECT 105.840 185.205 106.130 185.250 ;
        RECT 122.420 185.190 122.740 185.450 ;
        RECT 124.810 185.390 124.950 185.590 ;
        RECT 140.360 185.530 140.680 185.790 ;
        RECT 152.320 185.730 152.640 185.790 ;
        RECT 140.910 185.590 152.640 185.730 ;
        RECT 133.920 185.390 134.240 185.450 ;
        RECT 124.810 185.250 134.240 185.390 ;
        RECT 133.920 185.190 134.240 185.250 ;
        RECT 134.380 185.390 134.700 185.450 ;
        RECT 140.910 185.390 141.050 185.590 ;
        RECT 152.320 185.530 152.640 185.590 ;
        RECT 134.380 185.250 141.050 185.390 ;
        RECT 141.425 185.390 141.715 185.435 ;
        RECT 142.200 185.390 142.520 185.450 ;
        RECT 141.425 185.250 142.520 185.390 ;
        RECT 134.380 185.190 134.700 185.250 ;
        RECT 141.425 185.205 141.715 185.250 ;
        RECT 142.200 185.190 142.520 185.250 ;
        RECT 2.750 184.570 159.030 185.050 ;
        RECT 6.040 184.370 6.360 184.430 ;
        RECT 6.975 184.370 7.265 184.415 ;
        RECT 6.040 184.230 7.265 184.370 ;
        RECT 6.040 184.170 6.360 184.230 ;
        RECT 6.975 184.185 7.265 184.230 ;
        RECT 8.355 184.185 8.645 184.415 ;
        RECT 7.895 183.690 8.185 183.735 ;
        RECT 8.430 183.690 8.570 184.185 ;
        RECT 10.640 184.170 10.960 184.430 ;
        RECT 16.175 184.370 16.465 184.415 ;
        RECT 19.840 184.370 20.160 184.430 ;
        RECT 16.175 184.230 20.160 184.370 ;
        RECT 16.175 184.185 16.465 184.230 ;
        RECT 19.840 184.170 20.160 184.230 ;
        RECT 23.520 184.170 23.840 184.430 ;
        RECT 23.980 184.370 24.300 184.430 ;
        RECT 27.215 184.370 27.505 184.415 ;
        RECT 23.980 184.230 27.505 184.370 ;
        RECT 23.980 184.170 24.300 184.230 ;
        RECT 27.215 184.185 27.505 184.230 ;
        RECT 28.120 184.370 28.440 184.430 ;
        RECT 30.420 184.370 30.740 184.430 ;
        RECT 31.355 184.370 31.645 184.415 ;
        RECT 28.120 184.230 31.645 184.370 ;
        RECT 28.120 184.170 28.440 184.230 ;
        RECT 30.420 184.170 30.740 184.230 ;
        RECT 31.355 184.185 31.645 184.230 ;
        RECT 35.035 184.370 35.325 184.415 ;
        RECT 35.480 184.370 35.800 184.430 ;
        RECT 35.035 184.230 35.800 184.370 ;
        RECT 35.035 184.185 35.325 184.230 ;
        RECT 35.480 184.170 35.800 184.230 ;
        RECT 36.875 184.370 37.165 184.415 ;
        RECT 39.620 184.370 39.940 184.430 ;
        RECT 36.875 184.230 39.940 184.370 ;
        RECT 36.875 184.185 37.165 184.230 ;
        RECT 39.620 184.170 39.940 184.230 ;
        RECT 43.300 184.170 43.620 184.430 ;
        RECT 46.060 184.370 46.380 184.430 ;
        RECT 43.850 184.230 46.380 184.370 ;
        RECT 10.730 184.030 10.870 184.170 ;
        RECT 18.575 184.030 18.865 184.075 ;
        RECT 21.815 184.030 22.465 184.075 ;
        RECT 23.610 184.030 23.750 184.170 ;
        RECT 10.730 183.890 11.330 184.030 ;
        RECT 7.895 183.550 8.570 183.690 ;
        RECT 8.800 183.690 9.120 183.750 ;
        RECT 10.195 183.690 10.485 183.735 ;
        RECT 8.800 183.550 10.485 183.690 ;
        RECT 7.895 183.505 8.185 183.550 ;
        RECT 8.800 183.490 9.120 183.550 ;
        RECT 10.195 183.505 10.485 183.550 ;
        RECT 10.270 183.010 10.410 183.505 ;
        RECT 10.640 183.150 10.960 183.410 ;
        RECT 11.190 183.395 11.330 183.890 ;
        RECT 18.575 183.890 23.750 184.030 ;
        RECT 37.780 184.030 38.100 184.090 ;
        RECT 38.715 184.030 39.005 184.075 ;
        RECT 37.780 183.890 39.005 184.030 ;
        RECT 18.575 183.845 19.165 183.890 ;
        RECT 21.815 183.845 22.465 183.890 ;
        RECT 12.940 183.690 13.260 183.750 ;
        RECT 14.335 183.690 14.625 183.735 ;
        RECT 12.940 183.550 14.625 183.690 ;
        RECT 12.940 183.490 13.260 183.550 ;
        RECT 14.335 183.505 14.625 183.550 ;
        RECT 18.875 183.530 19.165 183.845 ;
        RECT 37.780 183.830 38.100 183.890 ;
        RECT 38.715 183.845 39.005 183.890 ;
        RECT 19.955 183.690 20.245 183.735 ;
        RECT 23.535 183.690 23.825 183.735 ;
        RECT 25.370 183.690 25.660 183.735 ;
        RECT 19.955 183.550 25.660 183.690 ;
        RECT 19.955 183.505 20.245 183.550 ;
        RECT 23.535 183.505 23.825 183.550 ;
        RECT 25.370 183.505 25.660 183.550 ;
        RECT 25.835 183.690 26.125 183.735 ;
        RECT 27.660 183.690 27.980 183.750 ;
        RECT 25.835 183.550 27.980 183.690 ;
        RECT 25.835 183.505 26.125 183.550 ;
        RECT 11.115 183.165 11.405 183.395 ;
        RECT 13.030 183.010 13.170 183.490 ;
        RECT 13.415 183.165 13.705 183.395 ;
        RECT 10.270 182.870 13.170 183.010 ;
        RECT 13.490 183.010 13.630 183.165 ;
        RECT 13.860 183.150 14.180 183.410 ;
        RECT 14.410 183.350 14.550 183.505 ;
        RECT 27.660 183.490 27.980 183.550 ;
        RECT 28.135 183.690 28.425 183.735 ;
        RECT 30.895 183.690 31.185 183.735 ;
        RECT 31.340 183.690 31.660 183.750 ;
        RECT 34.575 183.690 34.865 183.735 ;
        RECT 28.135 183.550 29.270 183.690 ;
        RECT 28.135 183.505 28.425 183.550 ;
        RECT 20.760 183.350 21.080 183.410 ;
        RECT 14.410 183.210 21.080 183.350 ;
        RECT 20.760 183.150 21.080 183.210 ;
        RECT 24.440 183.150 24.760 183.410 ;
        RECT 29.130 183.055 29.270 183.550 ;
        RECT 30.895 183.550 34.865 183.690 ;
        RECT 30.895 183.505 31.185 183.550 ;
        RECT 31.340 183.490 31.660 183.550 ;
        RECT 34.575 183.505 34.865 183.550 ;
        RECT 35.480 183.690 35.800 183.750 ;
        RECT 37.320 183.690 37.640 183.750 ;
        RECT 35.480 183.550 37.640 183.690 ;
        RECT 31.815 183.165 32.105 183.395 ;
        RECT 34.115 183.165 34.405 183.395 ;
        RECT 34.650 183.350 34.790 183.505 ;
        RECT 35.480 183.490 35.800 183.550 ;
        RECT 37.320 183.490 37.640 183.550 ;
        RECT 39.175 183.690 39.465 183.735 ;
        RECT 41.920 183.690 42.240 183.750 ;
        RECT 39.175 183.550 42.240 183.690 ;
        RECT 39.175 183.505 39.465 183.550 ;
        RECT 41.920 183.490 42.240 183.550 ;
        RECT 42.380 183.490 42.700 183.750 ;
        RECT 43.850 183.735 43.990 184.230 ;
        RECT 46.060 184.170 46.380 184.230 ;
        RECT 46.520 184.170 46.840 184.430 ;
        RECT 46.995 184.370 47.285 184.415 ;
        RECT 47.440 184.370 47.760 184.430 ;
        RECT 46.995 184.230 47.760 184.370 ;
        RECT 46.995 184.185 47.285 184.230 ;
        RECT 47.440 184.170 47.760 184.230 ;
        RECT 50.200 184.370 50.520 184.430 ;
        RECT 50.675 184.370 50.965 184.415 ;
        RECT 50.200 184.230 50.965 184.370 ;
        RECT 50.200 184.170 50.520 184.230 ;
        RECT 50.675 184.185 50.965 184.230 ;
        RECT 51.580 184.170 51.900 184.430 ;
        RECT 68.140 184.370 68.460 184.430 ;
        RECT 57.190 184.230 68.460 184.370 ;
        RECT 46.610 184.030 46.750 184.170 ;
        RECT 44.770 183.890 46.750 184.030 ;
        RECT 47.900 184.030 48.220 184.090 ;
        RECT 49.295 184.030 49.585 184.075 ;
        RECT 47.900 183.890 49.585 184.030 ;
        RECT 44.770 183.735 44.910 183.890 ;
        RECT 47.900 183.830 48.220 183.890 ;
        RECT 49.295 183.845 49.585 183.890 ;
        RECT 43.775 183.505 44.065 183.735 ;
        RECT 44.515 183.550 44.910 183.735 ;
        RECT 44.515 183.505 44.805 183.550 ;
        RECT 45.140 183.490 45.460 183.750 ;
        RECT 45.615 183.505 45.905 183.735 ;
        RECT 46.305 183.690 46.595 183.735 ;
        RECT 50.200 183.690 50.520 183.750 ;
        RECT 51.670 183.690 51.810 184.170 ;
        RECT 46.305 183.550 51.810 183.690 ;
        RECT 46.305 183.505 46.595 183.550 ;
        RECT 36.400 183.350 36.720 183.410 ;
        RECT 34.650 183.210 36.720 183.350 ;
        RECT 19.955 183.010 20.245 183.055 ;
        RECT 23.075 183.010 23.365 183.055 ;
        RECT 24.965 183.010 25.255 183.055 ;
        RECT 13.490 182.870 19.610 183.010 ;
        RECT 17.095 182.670 17.385 182.715 ;
        RECT 17.540 182.670 17.860 182.730 ;
        RECT 17.095 182.530 17.860 182.670 ;
        RECT 19.470 182.670 19.610 182.870 ;
        RECT 19.955 182.870 25.255 183.010 ;
        RECT 19.955 182.825 20.245 182.870 ;
        RECT 23.075 182.825 23.365 182.870 ;
        RECT 24.965 182.825 25.255 182.870 ;
        RECT 29.055 182.825 29.345 183.055 ;
        RECT 22.600 182.670 22.920 182.730 ;
        RECT 19.470 182.530 22.920 182.670 ;
        RECT 31.890 182.670 32.030 183.165 ;
        RECT 34.190 183.010 34.330 183.165 ;
        RECT 36.400 183.150 36.720 183.210 ;
        RECT 38.240 183.150 38.560 183.410 ;
        RECT 41.460 183.150 41.780 183.410 ;
        RECT 42.010 183.350 42.150 183.490 ;
        RECT 45.690 183.350 45.830 183.505 ;
        RECT 50.200 183.490 50.520 183.550 ;
        RECT 55.720 183.490 56.040 183.750 ;
        RECT 56.180 183.690 56.500 183.750 ;
        RECT 57.190 183.735 57.330 184.230 ;
        RECT 68.140 184.170 68.460 184.230 ;
        RECT 77.340 184.370 77.660 184.430 ;
        RECT 81.035 184.370 81.325 184.415 ;
        RECT 81.480 184.370 81.800 184.430 ;
        RECT 77.340 184.230 78.950 184.370 ;
        RECT 77.340 184.170 77.660 184.230 ;
        RECT 59.860 184.030 60.180 184.090 ;
        RECT 58.110 183.890 60.180 184.030 ;
        RECT 56.655 183.690 56.945 183.735 ;
        RECT 56.180 183.550 56.945 183.690 ;
        RECT 56.180 183.490 56.500 183.550 ;
        RECT 56.655 183.505 56.945 183.550 ;
        RECT 57.115 183.505 57.405 183.735 ;
        RECT 57.575 183.690 57.865 183.735 ;
        RECT 58.110 183.690 58.250 183.890 ;
        RECT 59.860 183.830 60.180 183.890 ;
        RECT 62.620 184.030 62.940 184.090 ;
        RECT 72.740 184.030 73.060 184.090 ;
        RECT 74.120 184.030 74.440 184.090 ;
        RECT 76.880 184.030 77.200 184.090 ;
        RECT 78.810 184.030 78.950 184.230 ;
        RECT 81.035 184.230 81.800 184.370 ;
        RECT 81.035 184.185 81.325 184.230 ;
        RECT 81.480 184.170 81.800 184.230 ;
        RECT 82.415 184.370 82.705 184.415 ;
        RECT 82.860 184.370 83.180 184.430 ;
        RECT 82.415 184.230 83.180 184.370 ;
        RECT 82.415 184.185 82.705 184.230 ;
        RECT 82.860 184.170 83.180 184.230 ;
        RECT 84.715 184.370 85.005 184.415 ;
        RECT 86.080 184.370 86.400 184.430 ;
        RECT 84.715 184.230 86.400 184.370 ;
        RECT 84.715 184.185 85.005 184.230 ;
        RECT 86.080 184.170 86.400 184.230 ;
        RECT 87.000 184.170 87.320 184.430 ;
        RECT 90.220 184.370 90.540 184.430 ;
        RECT 90.695 184.370 90.985 184.415 ;
        RECT 90.220 184.230 90.985 184.370 ;
        RECT 90.220 184.170 90.540 184.230 ;
        RECT 90.695 184.185 90.985 184.230 ;
        RECT 96.660 184.170 96.980 184.430 ;
        RECT 97.135 184.370 97.425 184.415 ;
        RECT 97.580 184.370 97.900 184.430 ;
        RECT 97.135 184.230 97.900 184.370 ;
        RECT 97.135 184.185 97.425 184.230 ;
        RECT 97.580 184.170 97.900 184.230 ;
        RECT 98.975 184.370 99.265 184.415 ;
        RECT 104.940 184.370 105.260 184.430 ;
        RECT 98.975 184.230 105.260 184.370 ;
        RECT 98.975 184.185 99.265 184.230 ;
        RECT 104.940 184.170 105.260 184.230 ;
        RECT 106.320 184.370 106.640 184.430 ;
        RECT 107.255 184.370 107.545 184.415 ;
        RECT 106.320 184.230 107.545 184.370 ;
        RECT 106.320 184.170 106.640 184.230 ;
        RECT 107.255 184.185 107.545 184.230 ;
        RECT 109.540 184.170 109.860 184.430 ;
        RECT 111.840 184.370 112.160 184.430 ;
        RECT 119.215 184.370 119.505 184.415 ;
        RECT 122.895 184.370 123.185 184.415 ;
        RECT 123.340 184.370 123.660 184.430 ;
        RECT 126.115 184.370 126.405 184.415 ;
        RECT 131.160 184.370 131.480 184.430 ;
        RECT 111.840 184.230 119.505 184.370 ;
        RECT 111.840 184.170 112.160 184.230 ;
        RECT 119.215 184.185 119.505 184.230 ;
        RECT 120.670 184.230 126.405 184.370 ;
        RECT 85.160 184.030 85.480 184.090 ;
        RECT 87.090 184.030 87.230 184.170 ;
        RECT 89.775 184.030 90.065 184.075 ;
        RECT 92.075 184.030 92.365 184.075 ;
        RECT 99.880 184.030 100.200 184.090 ;
        RECT 117.360 184.030 117.680 184.090 ;
        RECT 62.620 183.890 73.060 184.030 ;
        RECT 62.620 183.830 62.940 183.890 ;
        RECT 72.740 183.830 73.060 183.890 ;
        RECT 73.750 183.890 78.025 184.030 ;
        RECT 57.575 183.550 58.250 183.690 ;
        RECT 57.575 183.505 57.865 183.550 ;
        RECT 48.820 183.350 49.140 183.410 ;
        RECT 42.010 183.210 45.830 183.350 ;
        RECT 46.150 183.210 49.140 183.350 ;
        RECT 38.330 183.010 38.470 183.150 ;
        RECT 34.190 182.870 38.470 183.010 ;
        RECT 41.015 183.010 41.305 183.055 ;
        RECT 46.150 183.010 46.290 183.210 ;
        RECT 48.820 183.150 49.140 183.210 ;
        RECT 49.280 183.350 49.600 183.410 ;
        RECT 51.580 183.350 51.900 183.410 ;
        RECT 53.435 183.350 53.725 183.395 ;
        RECT 55.260 183.350 55.580 183.410 ;
        RECT 49.280 183.210 51.355 183.350 ;
        RECT 49.280 183.150 49.600 183.210 ;
        RECT 41.015 182.870 46.290 183.010 ;
        RECT 46.980 183.010 47.300 183.070 ;
        RECT 47.455 183.010 47.745 183.055 ;
        RECT 50.660 183.010 50.980 183.070 ;
        RECT 46.980 182.870 47.745 183.010 ;
        RECT 41.015 182.825 41.305 182.870 ;
        RECT 46.980 182.810 47.300 182.870 ;
        RECT 47.455 182.825 47.745 182.870 ;
        RECT 49.370 182.870 50.980 183.010 ;
        RECT 51.215 183.010 51.355 183.210 ;
        RECT 51.580 183.210 55.580 183.350 ;
        RECT 51.580 183.150 51.900 183.210 ;
        RECT 53.435 183.165 53.725 183.210 ;
        RECT 55.260 183.150 55.580 183.210 ;
        RECT 58.110 183.010 58.250 183.550 ;
        RECT 58.480 183.490 58.800 183.750 ;
        RECT 60.795 183.690 61.085 183.735 ;
        RECT 59.950 183.550 61.085 183.690 ;
        RECT 59.400 183.150 59.720 183.410 ;
        RECT 59.950 183.070 60.090 183.550 ;
        RECT 60.795 183.505 61.085 183.550 ;
        RECT 63.095 183.690 63.385 183.735 ;
        RECT 64.000 183.690 64.320 183.750 ;
        RECT 63.095 183.550 64.320 183.690 ;
        RECT 63.095 183.505 63.385 183.550 ;
        RECT 64.000 183.490 64.320 183.550 ;
        RECT 64.935 183.505 65.225 183.735 ;
        RECT 67.695 183.690 67.985 183.735 ;
        RECT 69.520 183.690 69.840 183.750 ;
        RECT 67.695 183.550 69.840 183.690 ;
        RECT 67.695 183.505 67.985 183.550 ;
        RECT 62.175 183.350 62.465 183.395 ;
        RECT 65.010 183.350 65.150 183.505 ;
        RECT 60.870 183.210 65.150 183.350 ;
        RECT 65.395 183.350 65.685 183.395 ;
        RECT 67.220 183.350 67.540 183.410 ;
        RECT 65.395 183.210 67.540 183.350 ;
        RECT 51.215 182.870 58.250 183.010 ;
        RECT 35.020 182.670 35.340 182.730 ;
        RECT 37.320 182.670 37.640 182.730 ;
        RECT 31.890 182.530 37.640 182.670 ;
        RECT 17.095 182.485 17.385 182.530 ;
        RECT 17.540 182.470 17.860 182.530 ;
        RECT 22.600 182.470 22.920 182.530 ;
        RECT 35.020 182.470 35.340 182.530 ;
        RECT 37.320 182.470 37.640 182.530 ;
        RECT 42.380 182.670 42.700 182.730 ;
        RECT 45.600 182.670 45.920 182.730 ;
        RECT 42.380 182.530 45.920 182.670 ;
        RECT 42.380 182.470 42.700 182.530 ;
        RECT 45.600 182.470 45.920 182.530 ;
        RECT 46.060 182.670 46.380 182.730 ;
        RECT 48.360 182.670 48.680 182.730 ;
        RECT 49.370 182.715 49.510 182.870 ;
        RECT 50.660 182.810 50.980 182.870 ;
        RECT 59.860 182.810 60.180 183.070 ;
        RECT 46.060 182.530 48.680 182.670 ;
        RECT 46.060 182.470 46.380 182.530 ;
        RECT 48.360 182.470 48.680 182.530 ;
        RECT 49.295 182.485 49.585 182.715 ;
        RECT 50.215 182.670 50.505 182.715 ;
        RECT 51.120 182.670 51.440 182.730 ;
        RECT 50.215 182.530 51.440 182.670 ;
        RECT 50.215 182.485 50.505 182.530 ;
        RECT 51.120 182.470 51.440 182.530 ;
        RECT 58.020 182.670 58.340 182.730 ;
        RECT 60.870 182.670 61.010 183.210 ;
        RECT 62.175 183.165 62.465 183.210 ;
        RECT 65.395 183.165 65.685 183.210 ;
        RECT 67.220 183.150 67.540 183.210 ;
        RECT 61.255 183.010 61.545 183.055 ;
        RECT 67.770 183.010 67.910 183.505 ;
        RECT 69.520 183.490 69.840 183.550 ;
        RECT 73.200 183.490 73.520 183.750 ;
        RECT 73.750 183.735 73.890 183.890 ;
        RECT 74.120 183.830 74.440 183.890 ;
        RECT 76.880 183.830 77.200 183.890 ;
        RECT 73.675 183.505 73.965 183.735 ;
        RECT 75.040 183.690 75.360 183.750 ;
        RECT 77.340 183.690 77.660 183.750 ;
        RECT 77.885 183.735 78.025 183.890 ;
        RECT 78.810 183.890 85.480 184.030 ;
        RECT 75.040 183.550 77.660 183.690 ;
        RECT 75.040 183.490 75.360 183.550 ;
        RECT 77.340 183.490 77.660 183.550 ;
        RECT 77.810 183.505 78.100 183.735 ;
        RECT 78.260 183.490 78.580 183.750 ;
        RECT 78.810 183.735 78.950 183.890 ;
        RECT 80.650 183.735 80.790 183.890 ;
        RECT 85.160 183.830 85.480 183.890 ;
        RECT 85.710 183.890 86.770 184.030 ;
        RECT 87.090 183.890 89.530 184.030 ;
        RECT 78.735 183.505 79.025 183.735 ;
        RECT 79.655 183.505 79.945 183.735 ;
        RECT 80.575 183.505 80.865 183.735 ;
        RECT 81.495 183.505 81.785 183.735 ;
        RECT 85.710 183.690 85.850 183.890 ;
        RECT 82.950 183.550 85.850 183.690 ;
        RECT 86.630 183.690 86.770 183.890 ;
        RECT 89.390 183.735 89.530 183.890 ;
        RECT 89.775 183.890 97.350 184.030 ;
        RECT 89.775 183.845 90.065 183.890 ;
        RECT 92.075 183.845 92.365 183.890 ;
        RECT 97.210 183.750 97.350 183.890 ;
        RECT 99.880 183.890 117.680 184.030 ;
        RECT 99.880 183.830 100.200 183.890 ;
        RECT 117.360 183.830 117.680 183.890 ;
        RECT 87.015 183.690 87.305 183.735 ;
        RECT 86.630 183.550 87.305 183.690 ;
        RECT 68.615 183.165 68.905 183.395 ;
        RECT 71.820 183.350 72.140 183.410 ;
        RECT 75.515 183.350 75.805 183.395 ;
        RECT 79.730 183.350 79.870 183.505 ;
        RECT 81.570 183.350 81.710 183.505 ;
        RECT 82.950 183.410 83.090 183.550 ;
        RECT 87.015 183.505 87.305 183.550 ;
        RECT 89.315 183.505 89.605 183.735 ;
        RECT 90.220 183.490 90.540 183.750 ;
        RECT 92.980 183.735 93.300 183.750 ;
        RECT 91.615 183.505 91.905 183.735 ;
        RECT 92.535 183.505 92.825 183.735 ;
        RECT 92.980 183.690 93.515 183.735 ;
        RECT 96.200 183.690 96.520 183.750 ;
        RECT 92.980 183.550 96.520 183.690 ;
        RECT 92.980 183.505 93.515 183.550 ;
        RECT 82.860 183.350 83.180 183.410 ;
        RECT 71.820 183.210 83.180 183.350 ;
        RECT 61.255 182.870 67.910 183.010 ;
        RECT 61.255 182.825 61.545 182.870 ;
        RECT 58.020 182.530 61.010 182.670 ;
        RECT 67.220 182.670 67.540 182.730 ;
        RECT 68.690 182.670 68.830 183.165 ;
        RECT 71.820 183.150 72.140 183.210 ;
        RECT 75.515 183.165 75.805 183.210 ;
        RECT 82.860 183.150 83.180 183.210 ;
        RECT 83.320 183.150 83.640 183.410 ;
        RECT 83.780 183.150 84.100 183.410 ;
        RECT 85.175 183.165 85.465 183.395 ;
        RECT 76.435 183.010 76.725 183.055 ;
        RECT 82.400 183.010 82.720 183.070 ;
        RECT 76.435 182.870 82.720 183.010 ;
        RECT 76.435 182.825 76.725 182.870 ;
        RECT 82.400 182.810 82.720 182.870 ;
        RECT 67.220 182.530 68.830 182.670 ;
        RECT 58.020 182.470 58.340 182.530 ;
        RECT 67.220 182.470 67.540 182.530 ;
        RECT 70.440 182.470 70.760 182.730 ;
        RECT 81.940 182.670 82.260 182.730 ;
        RECT 85.250 182.670 85.390 183.165 ;
        RECT 85.620 183.150 85.940 183.410 ;
        RECT 86.095 183.165 86.385 183.395 ;
        RECT 86.540 183.350 86.860 183.410 ;
        RECT 91.140 183.350 91.460 183.410 ;
        RECT 91.690 183.350 91.830 183.505 ;
        RECT 92.060 183.350 92.380 183.410 ;
        RECT 86.540 183.210 92.380 183.350 ;
        RECT 86.170 183.010 86.310 183.165 ;
        RECT 86.540 183.150 86.860 183.210 ;
        RECT 91.140 183.150 91.460 183.210 ;
        RECT 92.060 183.150 92.380 183.210 ;
        RECT 85.710 182.870 86.310 183.010 ;
        RECT 85.710 182.730 85.850 182.870 ;
        RECT 87.935 182.825 88.225 183.055 ;
        RECT 89.760 183.010 90.080 183.070 ;
        RECT 92.610 183.010 92.750 183.505 ;
        RECT 92.980 183.490 93.300 183.505 ;
        RECT 96.200 183.490 96.520 183.550 ;
        RECT 97.120 183.490 97.440 183.750 ;
        RECT 97.595 183.690 97.885 183.735 ;
        RECT 98.960 183.690 99.280 183.750 ;
        RECT 102.180 183.690 102.500 183.750 ;
        RECT 97.595 183.550 99.280 183.690 ;
        RECT 97.595 183.505 97.885 183.550 ;
        RECT 98.960 183.490 99.280 183.550 ;
        RECT 99.470 183.550 102.500 183.690 ;
        RECT 93.900 183.350 94.220 183.410 ;
        RECT 94.820 183.350 95.140 183.410 ;
        RECT 93.900 183.210 95.140 183.350 ;
        RECT 93.900 183.150 94.220 183.210 ;
        RECT 94.820 183.150 95.140 183.210 ;
        RECT 95.280 183.150 95.600 183.410 ;
        RECT 95.755 183.350 96.045 183.395 ;
        RECT 96.660 183.350 96.980 183.410 ;
        RECT 99.470 183.350 99.610 183.550 ;
        RECT 102.180 183.490 102.500 183.550 ;
        RECT 102.655 183.690 102.945 183.735 ;
        RECT 114.600 183.690 114.920 183.750 ;
        RECT 116.900 183.690 117.220 183.750 ;
        RECT 102.655 183.550 117.220 183.690 ;
        RECT 102.655 183.505 102.945 183.550 ;
        RECT 114.600 183.490 114.920 183.550 ;
        RECT 116.900 183.490 117.220 183.550 ;
        RECT 119.200 183.690 119.520 183.750 ;
        RECT 120.670 183.735 120.810 184.230 ;
        RECT 122.895 184.185 123.185 184.230 ;
        RECT 123.340 184.170 123.660 184.230 ;
        RECT 126.115 184.185 126.405 184.230 ;
        RECT 129.870 184.230 131.480 184.370 ;
        RECT 124.260 184.030 124.580 184.090 ;
        RECT 124.735 184.030 125.025 184.075 ;
        RECT 128.860 184.030 129.180 184.090 ;
        RECT 121.130 183.890 124.030 184.030 ;
        RECT 120.595 183.690 120.885 183.735 ;
        RECT 119.200 183.550 120.885 183.690 ;
        RECT 119.200 183.490 119.520 183.550 ;
        RECT 120.595 183.505 120.885 183.550 ;
        RECT 100.800 183.350 101.120 183.410 ;
        RECT 95.755 183.210 99.610 183.350 ;
        RECT 100.430 183.210 101.120 183.350 ;
        RECT 95.755 183.165 96.045 183.210 ;
        RECT 96.660 183.150 96.980 183.210 ;
        RECT 100.430 183.010 100.570 183.210 ;
        RECT 100.800 183.150 101.120 183.210 ;
        RECT 101.720 183.350 102.040 183.410 ;
        RECT 103.115 183.350 103.405 183.395 ;
        RECT 106.780 183.350 107.100 183.410 ;
        RECT 101.720 183.210 107.100 183.350 ;
        RECT 101.720 183.150 102.040 183.210 ;
        RECT 103.115 183.165 103.405 183.210 ;
        RECT 106.780 183.150 107.100 183.210 ;
        RECT 107.700 183.350 108.020 183.410 ;
        RECT 108.175 183.350 108.465 183.395 ;
        RECT 107.700 183.210 108.465 183.350 ;
        RECT 107.700 183.150 108.020 183.210 ;
        RECT 108.175 183.165 108.465 183.210 ;
        RECT 108.620 183.150 108.940 183.410 ;
        RECT 110.015 183.165 110.305 183.395 ;
        RECT 89.760 182.870 100.570 183.010 ;
        RECT 102.180 183.010 102.500 183.070 ;
        RECT 110.090 183.010 110.230 183.165 ;
        RECT 110.460 183.150 110.780 183.410 ;
        RECT 115.060 183.350 115.380 183.410 ;
        RECT 118.755 183.350 119.045 183.395 ;
        RECT 121.130 183.350 121.270 183.890 ;
        RECT 123.890 183.750 124.030 183.890 ;
        RECT 124.260 183.890 129.180 184.030 ;
        RECT 124.260 183.830 124.580 183.890 ;
        RECT 124.735 183.845 125.025 183.890 ;
        RECT 128.860 183.830 129.180 183.890 ;
        RECT 122.435 183.505 122.725 183.735 ;
        RECT 115.060 183.210 121.270 183.350 ;
        RECT 121.515 183.350 121.805 183.395 ;
        RECT 122.510 183.350 122.650 183.505 ;
        RECT 123.800 183.490 124.120 183.750 ;
        RECT 125.655 183.505 125.945 183.735 ;
        RECT 126.100 183.690 126.420 183.750 ;
        RECT 127.035 183.690 127.325 183.735 ;
        RECT 126.100 183.550 127.325 183.690 ;
        RECT 125.730 183.350 125.870 183.505 ;
        RECT 126.100 183.490 126.420 183.550 ;
        RECT 127.035 183.505 127.325 183.550 ;
        RECT 129.320 183.490 129.640 183.750 ;
        RECT 129.870 183.735 130.010 184.230 ;
        RECT 131.160 184.170 131.480 184.230 ;
        RECT 133.015 184.370 133.305 184.415 ;
        RECT 133.460 184.370 133.780 184.430 ;
        RECT 133.015 184.230 133.780 184.370 ;
        RECT 133.015 184.185 133.305 184.230 ;
        RECT 133.460 184.170 133.780 184.230 ;
        RECT 135.760 184.370 136.080 184.430 ;
        RECT 141.280 184.370 141.600 184.430 ;
        RECT 135.760 184.230 141.600 184.370 ;
        RECT 135.760 184.170 136.080 184.230 ;
        RECT 137.140 184.030 137.460 184.090 ;
        RECT 131.250 183.890 138.290 184.030 ;
        RECT 131.250 183.735 131.390 183.890 ;
        RECT 137.140 183.830 137.460 183.890 ;
        RECT 129.795 183.505 130.085 183.735 ;
        RECT 131.175 183.505 131.465 183.735 ;
        RECT 129.870 183.350 130.010 183.505 ;
        RECT 133.000 183.490 133.320 183.750 ;
        RECT 133.920 183.490 134.240 183.750 ;
        RECT 138.150 183.735 138.290 183.890 ;
        RECT 138.610 183.735 138.750 184.230 ;
        RECT 141.280 184.170 141.600 184.230 ;
        RECT 149.100 184.370 149.420 184.430 ;
        RECT 150.035 184.370 150.325 184.415 ;
        RECT 149.100 184.230 150.325 184.370 ;
        RECT 149.100 184.170 149.420 184.230 ;
        RECT 150.035 184.185 150.325 184.230 ;
        RECT 150.480 184.370 150.800 184.430 ;
        RECT 152.320 184.370 152.640 184.430 ;
        RECT 154.620 184.370 154.940 184.430 ;
        RECT 150.480 184.230 154.940 184.370 ;
        RECT 150.480 184.170 150.800 184.230 ;
        RECT 152.320 184.170 152.640 184.230 ;
        RECT 154.620 184.170 154.940 184.230 ;
        RECT 155.095 184.370 155.385 184.415 ;
        RECT 155.540 184.370 155.860 184.430 ;
        RECT 155.095 184.230 155.860 184.370 ;
        RECT 155.095 184.185 155.385 184.230 ;
        RECT 155.540 184.170 155.860 184.230 ;
        RECT 141.370 184.030 141.510 184.170 ;
        RECT 151.860 184.030 152.180 184.090 ;
        RECT 153.715 184.030 154.005 184.075 ;
        RECT 141.370 183.890 154.005 184.030 ;
        RECT 138.075 183.505 138.365 183.735 ;
        RECT 138.535 183.505 138.825 183.735 ;
        RECT 139.455 183.505 139.745 183.735 ;
        RECT 139.915 183.690 140.205 183.735 ;
        RECT 142.660 183.690 142.980 183.750 ;
        RECT 143.210 183.735 143.350 183.890 ;
        RECT 151.860 183.830 152.180 183.890 ;
        RECT 153.715 183.845 154.005 183.890 ;
        RECT 139.915 183.550 142.980 183.690 ;
        RECT 139.915 183.505 140.205 183.550 ;
        RECT 121.515 183.210 125.870 183.350 ;
        RECT 129.410 183.210 130.010 183.350 ;
        RECT 130.255 183.350 130.545 183.395 ;
        RECT 133.090 183.350 133.230 183.490 ;
        RECT 130.255 183.210 133.230 183.350 ;
        RECT 115.060 183.150 115.380 183.210 ;
        RECT 118.755 183.165 119.045 183.210 ;
        RECT 121.515 183.165 121.805 183.210 ;
        RECT 112.300 183.010 112.620 183.070 ;
        RECT 119.660 183.010 119.980 183.070 ;
        RECT 102.180 182.870 119.980 183.010 ;
        RECT 81.940 182.530 85.390 182.670 ;
        RECT 81.940 182.470 82.260 182.530 ;
        RECT 85.620 182.470 85.940 182.730 ;
        RECT 88.010 182.670 88.150 182.825 ;
        RECT 89.760 182.810 90.080 182.870 ;
        RECT 102.180 182.810 102.500 182.870 ;
        RECT 112.300 182.810 112.620 182.870 ;
        RECT 119.660 182.810 119.980 182.870 ;
        RECT 120.120 183.010 120.440 183.070 ;
        RECT 121.590 183.010 121.730 183.165 ;
        RECT 129.410 183.070 129.550 183.210 ;
        RECT 130.255 183.165 130.545 183.210 ;
        RECT 135.315 183.165 135.605 183.395 ;
        RECT 139.530 183.350 139.670 183.505 ;
        RECT 142.660 183.490 142.980 183.550 ;
        RECT 143.135 183.505 143.425 183.735 ;
        RECT 143.580 183.690 143.900 183.750 ;
        RECT 144.055 183.690 144.345 183.735 ;
        RECT 145.420 183.690 145.740 183.750 ;
        RECT 143.580 183.550 145.740 183.690 ;
        RECT 143.580 183.490 143.900 183.550 ;
        RECT 144.055 183.505 144.345 183.550 ;
        RECT 145.420 183.490 145.740 183.550 ;
        RECT 148.180 183.690 148.500 183.750 ;
        RECT 148.655 183.690 148.945 183.735 ;
        RECT 148.180 183.550 148.945 183.690 ;
        RECT 148.180 183.490 148.500 183.550 ;
        RECT 148.655 183.505 148.945 183.550 ;
        RECT 149.575 183.690 149.865 183.735 ;
        RECT 150.020 183.690 150.340 183.750 ;
        RECT 152.335 183.690 152.625 183.735 ;
        RECT 149.575 183.550 152.625 183.690 ;
        RECT 149.575 183.505 149.865 183.550 ;
        RECT 150.020 183.490 150.340 183.550 ;
        RECT 152.335 183.505 152.625 183.550 ;
        RECT 154.160 183.490 154.480 183.750 ;
        RECT 155.080 183.490 155.400 183.750 ;
        RECT 150.480 183.350 150.800 183.410 ;
        RECT 150.955 183.350 151.245 183.395 ;
        RECT 139.530 183.210 140.130 183.350 ;
        RECT 120.120 182.870 121.730 183.010 ;
        RECT 120.120 182.810 120.440 182.870 ;
        RECT 129.320 182.810 129.640 183.070 ;
        RECT 131.175 183.010 131.465 183.055 ;
        RECT 135.390 183.010 135.530 183.165 ;
        RECT 131.175 182.870 135.530 183.010 ;
        RECT 131.175 182.825 131.465 182.870 ;
        RECT 139.990 182.730 140.130 183.210 ;
        RECT 150.480 183.210 151.245 183.350 ;
        RECT 150.480 183.150 150.800 183.210 ;
        RECT 150.955 183.165 151.245 183.210 ;
        RECT 151.415 183.165 151.705 183.395 ;
        RECT 151.875 183.350 152.165 183.395 ;
        RECT 154.250 183.350 154.390 183.490 ;
        RECT 151.875 183.210 154.390 183.350 ;
        RECT 151.875 183.165 152.165 183.210 ;
        RECT 151.490 183.010 151.630 183.165 ;
        RECT 155.170 183.010 155.310 183.490 ;
        RECT 151.490 182.870 155.310 183.010 ;
        RECT 151.950 182.730 152.090 182.870 ;
        RECT 95.740 182.670 96.060 182.730 ;
        RECT 88.010 182.530 96.060 182.670 ;
        RECT 95.740 182.470 96.060 182.530 ;
        RECT 96.200 182.670 96.520 182.730 ;
        RECT 102.655 182.670 102.945 182.715 ;
        RECT 103.100 182.670 103.420 182.730 ;
        RECT 96.200 182.530 103.420 182.670 ;
        RECT 96.200 182.470 96.520 182.530 ;
        RECT 102.655 182.485 102.945 182.530 ;
        RECT 103.100 182.470 103.420 182.530 ;
        RECT 104.495 182.670 104.785 182.715 ;
        RECT 105.860 182.670 106.180 182.730 ;
        RECT 104.495 182.530 106.180 182.670 ;
        RECT 104.495 182.485 104.785 182.530 ;
        RECT 105.860 182.470 106.180 182.530 ;
        RECT 114.140 182.670 114.460 182.730 ;
        RECT 115.980 182.670 116.300 182.730 ;
        RECT 124.260 182.670 124.580 182.730 ;
        RECT 114.140 182.530 124.580 182.670 ;
        RECT 114.140 182.470 114.460 182.530 ;
        RECT 115.980 182.470 116.300 182.530 ;
        RECT 124.260 182.470 124.580 182.530 ;
        RECT 127.035 182.670 127.325 182.715 ;
        RECT 134.380 182.670 134.700 182.730 ;
        RECT 127.035 182.530 134.700 182.670 ;
        RECT 127.035 182.485 127.325 182.530 ;
        RECT 134.380 182.470 134.700 182.530 ;
        RECT 134.855 182.670 135.145 182.715 ;
        RECT 137.155 182.670 137.445 182.715 ;
        RECT 134.855 182.530 137.445 182.670 ;
        RECT 134.855 182.485 135.145 182.530 ;
        RECT 137.155 182.485 137.445 182.530 ;
        RECT 139.900 182.470 140.220 182.730 ;
        RECT 149.100 182.470 149.420 182.730 ;
        RECT 151.860 182.470 152.180 182.730 ;
        RECT 2.750 181.850 158.230 182.330 ;
        RECT 13.860 181.650 14.180 181.710 ;
        RECT 16.405 181.650 16.695 181.695 ;
        RECT 17.080 181.650 17.400 181.710 ;
        RECT 13.860 181.510 17.400 181.650 ;
        RECT 13.860 181.450 14.180 181.510 ;
        RECT 16.405 181.465 16.695 181.510 ;
        RECT 17.080 181.450 17.400 181.510 ;
        RECT 17.540 181.650 17.860 181.710 ;
        RECT 20.760 181.650 21.080 181.710 ;
        RECT 17.540 181.510 21.080 181.650 ;
        RECT 17.540 181.450 17.860 181.510 ;
        RECT 20.760 181.450 21.080 181.510 ;
        RECT 24.440 181.650 24.760 181.710 ;
        RECT 25.835 181.650 26.125 181.695 ;
        RECT 24.440 181.510 26.125 181.650 ;
        RECT 24.440 181.450 24.760 181.510 ;
        RECT 25.835 181.465 26.125 181.510 ;
        RECT 26.740 181.650 27.060 181.710 ;
        RECT 52.055 181.650 52.345 181.695 ;
        RECT 55.720 181.650 56.040 181.710 ;
        RECT 26.740 181.510 50.890 181.650 ;
        RECT 26.740 181.450 27.060 181.510 ;
        RECT 4.680 181.310 4.970 181.355 ;
        RECT 6.540 181.310 6.830 181.355 ;
        RECT 9.320 181.310 9.610 181.355 ;
        RECT 4.680 181.170 9.610 181.310 ;
        RECT 4.680 181.125 4.970 181.170 ;
        RECT 6.540 181.125 6.830 181.170 ;
        RECT 9.320 181.125 9.610 181.170 ;
        RECT 15.255 181.125 15.545 181.355 ;
        RECT 20.270 181.310 20.560 181.355 ;
        RECT 23.050 181.310 23.340 181.355 ;
        RECT 24.910 181.310 25.200 181.355 ;
        RECT 20.270 181.170 25.200 181.310 ;
        RECT 20.270 181.125 20.560 181.170 ;
        RECT 23.050 181.125 23.340 181.170 ;
        RECT 24.910 181.125 25.200 181.170 ;
        RECT 28.545 181.310 28.835 181.355 ;
        RECT 30.435 181.310 30.725 181.355 ;
        RECT 33.555 181.310 33.845 181.355 ;
        RECT 28.545 181.170 33.845 181.310 ;
        RECT 28.545 181.125 28.835 181.170 ;
        RECT 30.435 181.125 30.725 181.170 ;
        RECT 33.555 181.125 33.845 181.170 ;
        RECT 41.460 181.310 41.780 181.370 ;
        RECT 47.440 181.310 47.760 181.370 ;
        RECT 49.280 181.310 49.600 181.370 ;
        RECT 41.460 181.170 49.600 181.310 ;
        RECT 15.330 180.970 15.470 181.125 ;
        RECT 41.460 181.110 41.780 181.170 ;
        RECT 47.440 181.110 47.760 181.170 ;
        RECT 49.280 181.110 49.600 181.170 ;
        RECT 23.535 180.970 23.825 181.015 ;
        RECT 15.330 180.830 23.825 180.970 ;
        RECT 23.535 180.785 23.825 180.830 ;
        RECT 25.375 180.970 25.665 181.015 ;
        RECT 27.660 180.970 27.980 181.030 ;
        RECT 31.800 180.970 32.120 181.030 ;
        RECT 25.375 180.830 32.120 180.970 ;
        RECT 25.375 180.785 25.665 180.830 ;
        RECT 27.660 180.770 27.980 180.830 ;
        RECT 31.800 180.770 32.120 180.830 ;
        RECT 37.320 180.970 37.640 181.030 ;
        RECT 40.095 180.970 40.385 181.015 ;
        RECT 44.680 180.970 45.000 181.030 ;
        RECT 37.320 180.830 40.385 180.970 ;
        RECT 37.320 180.770 37.640 180.830 ;
        RECT 40.095 180.785 40.385 180.830 ;
        RECT 42.010 180.830 48.130 180.970 ;
        RECT 4.215 180.630 4.505 180.675 ;
        RECT 4.660 180.630 4.980 180.690 ;
        RECT 4.215 180.490 4.980 180.630 ;
        RECT 4.215 180.445 4.505 180.490 ;
        RECT 4.660 180.430 4.980 180.490 ;
        RECT 6.040 180.430 6.360 180.690 ;
        RECT 9.320 180.630 9.610 180.675 ;
        RECT 7.075 180.490 9.610 180.630 ;
        RECT 7.075 180.335 7.290 180.490 ;
        RECT 9.320 180.445 9.610 180.490 ;
        RECT 14.320 180.430 14.640 180.690 ;
        RECT 20.270 180.630 20.560 180.675 ;
        RECT 25.820 180.630 26.140 180.690 ;
        RECT 26.755 180.630 27.045 180.675 ;
        RECT 20.270 180.490 22.805 180.630 ;
        RECT 20.270 180.445 20.560 180.490 ;
        RECT 11.100 180.335 11.420 180.350 ;
        RECT 22.590 180.335 22.805 180.490 ;
        RECT 25.820 180.490 27.045 180.630 ;
        RECT 25.820 180.430 26.140 180.490 ;
        RECT 26.755 180.445 27.045 180.490 ;
        RECT 28.140 180.630 28.430 180.675 ;
        RECT 29.975 180.630 30.265 180.675 ;
        RECT 33.555 180.630 33.845 180.675 ;
        RECT 28.140 180.490 33.845 180.630 ;
        RECT 28.140 180.445 28.430 180.490 ;
        RECT 29.975 180.445 30.265 180.490 ;
        RECT 33.555 180.445 33.845 180.490 ;
        RECT 34.560 180.650 34.880 180.690 ;
        RECT 34.560 180.430 34.925 180.650 ;
        RECT 5.140 180.290 5.430 180.335 ;
        RECT 7.000 180.290 7.290 180.335 ;
        RECT 5.140 180.150 7.290 180.290 ;
        RECT 5.140 180.105 5.430 180.150 ;
        RECT 7.000 180.105 7.290 180.150 ;
        RECT 7.920 180.290 8.210 180.335 ;
        RECT 11.100 180.290 11.470 180.335 ;
        RECT 7.920 180.150 11.470 180.290 ;
        RECT 7.920 180.105 8.210 180.150 ;
        RECT 11.100 180.105 11.470 180.150 ;
        RECT 18.410 180.290 18.700 180.335 ;
        RECT 21.670 180.290 21.960 180.335 ;
        RECT 22.590 180.290 22.880 180.335 ;
        RECT 24.450 180.290 24.740 180.335 ;
        RECT 18.410 180.150 22.370 180.290 ;
        RECT 18.410 180.105 18.700 180.150 ;
        RECT 21.670 180.105 21.960 180.150 ;
        RECT 11.100 180.090 11.420 180.105 ;
        RECT 13.185 179.950 13.475 179.995 ;
        RECT 13.860 179.950 14.180 180.010 ;
        RECT 19.380 179.950 19.700 180.010 ;
        RECT 13.185 179.810 19.700 179.950 ;
        RECT 22.230 179.950 22.370 180.150 ;
        RECT 22.590 180.150 24.740 180.290 ;
        RECT 22.590 180.105 22.880 180.150 ;
        RECT 24.450 180.105 24.740 180.150 ;
        RECT 29.040 180.090 29.360 180.350 ;
        RECT 34.635 180.335 34.925 180.430 ;
        RECT 31.335 180.290 31.985 180.335 ;
        RECT 34.635 180.290 35.225 180.335 ;
        RECT 31.335 180.150 35.225 180.290 ;
        RECT 31.335 180.105 31.985 180.150 ;
        RECT 34.935 180.105 35.225 180.150 ;
        RECT 36.490 180.150 38.010 180.290 ;
        RECT 23.520 179.950 23.840 180.010 ;
        RECT 36.490 179.995 36.630 180.150 ;
        RECT 37.870 180.010 38.010 180.150 ;
        RECT 39.175 180.105 39.465 180.335 ;
        RECT 40.170 180.290 40.310 180.785 ;
        RECT 42.010 180.675 42.150 180.830 ;
        RECT 44.680 180.770 45.000 180.830 ;
        RECT 47.990 180.690 48.130 180.830 ;
        RECT 48.360 180.770 48.680 181.030 ;
        RECT 41.935 180.445 42.225 180.675 ;
        RECT 42.840 180.630 43.160 180.690 ;
        RECT 43.775 180.630 44.065 180.675 ;
        RECT 42.840 180.490 44.065 180.630 ;
        RECT 42.840 180.430 43.160 180.490 ;
        RECT 43.775 180.445 44.065 180.490 ;
        RECT 45.600 180.430 45.920 180.690 ;
        RECT 46.075 180.630 46.365 180.675 ;
        RECT 46.980 180.630 47.300 180.690 ;
        RECT 46.075 180.490 47.300 180.630 ;
        RECT 46.075 180.445 46.365 180.490 ;
        RECT 46.980 180.430 47.300 180.490 ;
        RECT 47.440 180.430 47.760 180.690 ;
        RECT 47.900 180.430 48.220 180.690 ;
        RECT 48.450 180.630 48.590 180.770 ;
        RECT 48.835 180.630 49.125 180.675 ;
        RECT 48.450 180.490 49.125 180.630 ;
        RECT 48.835 180.445 49.125 180.490 ;
        RECT 49.300 180.600 49.590 180.675 ;
        RECT 49.740 180.600 50.060 180.690 ;
        RECT 50.750 180.675 50.890 181.510 ;
        RECT 52.055 181.510 56.040 181.650 ;
        RECT 52.055 181.465 52.345 181.510 ;
        RECT 55.720 181.450 56.040 181.510 ;
        RECT 57.510 181.650 57.800 181.695 ;
        RECT 59.400 181.650 59.720 181.710 ;
        RECT 57.510 181.510 59.720 181.650 ;
        RECT 57.510 181.465 57.800 181.510 ;
        RECT 59.400 181.450 59.720 181.510 ;
        RECT 59.860 181.650 60.180 181.710 ;
        RECT 67.220 181.650 67.540 181.710 ;
        RECT 59.860 181.510 67.540 181.650 ;
        RECT 59.860 181.450 60.180 181.510 ;
        RECT 67.220 181.450 67.540 181.510 ;
        RECT 69.075 181.465 69.365 181.695 ;
        RECT 69.995 181.650 70.285 181.695 ;
        RECT 70.900 181.650 71.220 181.710 ;
        RECT 69.995 181.510 71.220 181.650 ;
        RECT 69.995 181.465 70.285 181.510 ;
        RECT 57.065 181.310 57.355 181.355 ;
        RECT 58.955 181.310 59.245 181.355 ;
        RECT 62.075 181.310 62.365 181.355 ;
        RECT 57.065 181.170 62.365 181.310 ;
        RECT 69.150 181.310 69.290 181.465 ;
        RECT 70.900 181.450 71.220 181.510 ;
        RECT 73.200 181.650 73.520 181.710 ;
        RECT 73.675 181.650 73.965 181.695 ;
        RECT 78.260 181.650 78.580 181.710 ;
        RECT 73.200 181.510 78.580 181.650 ;
        RECT 73.200 181.450 73.520 181.510 ;
        RECT 73.675 181.465 73.965 181.510 ;
        RECT 78.260 181.450 78.580 181.510 ;
        RECT 83.320 181.650 83.640 181.710 ;
        RECT 87.920 181.650 88.240 181.710 ;
        RECT 83.320 181.510 88.240 181.650 ;
        RECT 83.320 181.450 83.640 181.510 ;
        RECT 87.920 181.450 88.240 181.510 ;
        RECT 88.840 181.650 89.160 181.710 ;
        RECT 96.660 181.650 96.980 181.710 ;
        RECT 88.840 181.510 96.980 181.650 ;
        RECT 88.840 181.450 89.160 181.510 ;
        RECT 96.660 181.450 96.980 181.510 ;
        RECT 98.975 181.650 99.265 181.695 ;
        RECT 101.720 181.650 102.040 181.710 ;
        RECT 98.975 181.510 102.040 181.650 ;
        RECT 98.975 181.465 99.265 181.510 ;
        RECT 101.720 181.450 102.040 181.510 ;
        RECT 102.180 181.450 102.500 181.710 ;
        RECT 103.100 181.450 103.420 181.710 ;
        RECT 103.560 181.650 103.880 181.710 ;
        RECT 104.035 181.650 104.325 181.695 ;
        RECT 103.560 181.510 104.325 181.650 ;
        RECT 103.560 181.450 103.880 181.510 ;
        RECT 104.035 181.465 104.325 181.510 ;
        RECT 108.620 181.650 108.940 181.710 ;
        RECT 113.235 181.650 113.525 181.695 ;
        RECT 108.620 181.510 113.525 181.650 ;
        RECT 108.620 181.450 108.940 181.510 ;
        RECT 113.235 181.465 113.525 181.510 ;
        RECT 113.680 181.650 114.000 181.710 ;
        RECT 115.535 181.650 115.825 181.695 ;
        RECT 119.200 181.650 119.520 181.710 ;
        RECT 113.680 181.510 119.520 181.650 ;
        RECT 113.680 181.450 114.000 181.510 ;
        RECT 115.535 181.465 115.825 181.510 ;
        RECT 119.200 181.450 119.520 181.510 ;
        RECT 121.960 181.450 122.280 181.710 ;
        RECT 122.970 181.510 129.550 181.650 ;
        RECT 122.970 181.370 123.110 181.510 ;
        RECT 89.300 181.310 89.620 181.370 ;
        RECT 107.700 181.310 108.020 181.370 ;
        RECT 122.420 181.310 122.740 181.370 ;
        RECT 69.150 181.170 71.130 181.310 ;
        RECT 57.065 181.125 57.355 181.170 ;
        RECT 58.955 181.125 59.245 181.170 ;
        RECT 62.075 181.125 62.365 181.170 ;
        RECT 56.195 180.970 56.485 181.015 ;
        RECT 57.560 180.970 57.880 181.030 ;
        RECT 56.195 180.830 57.880 180.970 ;
        RECT 56.195 180.785 56.485 180.830 ;
        RECT 57.560 180.770 57.880 180.830 ;
        RECT 64.920 180.970 65.240 181.030 ;
        RECT 66.315 180.970 66.605 181.015 ;
        RECT 64.920 180.830 66.605 180.970 ;
        RECT 64.920 180.770 65.240 180.830 ;
        RECT 66.315 180.785 66.605 180.830 ;
        RECT 70.990 180.690 71.130 181.170 ;
        RECT 89.300 181.170 122.740 181.310 ;
        RECT 89.300 181.110 89.620 181.170 ;
        RECT 107.700 181.110 108.020 181.170 ;
        RECT 122.420 181.110 122.740 181.170 ;
        RECT 122.880 181.110 123.200 181.370 ;
        RECT 124.260 181.310 124.580 181.370 ;
        RECT 124.260 181.170 127.710 181.310 ;
        RECT 124.260 181.110 124.580 181.170 ;
        RECT 74.135 180.970 74.425 181.015 ;
        RECT 76.880 180.970 77.200 181.030 ;
        RECT 85.620 180.970 85.940 181.030 ;
        RECT 89.775 180.970 90.065 181.015 ;
        RECT 74.135 180.830 85.390 180.970 ;
        RECT 74.135 180.785 74.425 180.830 ;
        RECT 76.880 180.770 77.200 180.830 ;
        RECT 49.300 180.460 50.060 180.600 ;
        RECT 49.300 180.445 49.590 180.460 ;
        RECT 49.740 180.430 50.060 180.460 ;
        RECT 50.675 180.445 50.965 180.675 ;
        RECT 51.365 180.630 51.655 180.675 ;
        RECT 52.040 180.630 52.360 180.690 ;
        RECT 51.365 180.490 52.360 180.630 ;
        RECT 51.365 180.445 51.655 180.490 ;
        RECT 52.040 180.430 52.360 180.490 ;
        RECT 53.435 180.630 53.725 180.675 ;
        RECT 53.880 180.630 54.200 180.690 ;
        RECT 53.435 180.490 54.200 180.630 ;
        RECT 53.435 180.445 53.725 180.490 ;
        RECT 53.880 180.430 54.200 180.490 ;
        RECT 54.815 180.445 55.105 180.675 ;
        RECT 56.660 180.630 56.950 180.675 ;
        RECT 58.495 180.630 58.785 180.675 ;
        RECT 62.075 180.630 62.365 180.675 ;
        RECT 56.660 180.490 62.365 180.630 ;
        RECT 56.660 180.445 56.950 180.490 ;
        RECT 58.495 180.445 58.785 180.490 ;
        RECT 62.075 180.445 62.365 180.490 ;
        RECT 43.315 180.290 43.605 180.335 ;
        RECT 40.170 180.150 43.605 180.290 ;
        RECT 45.690 180.290 45.830 180.430 ;
        RECT 46.535 180.290 46.825 180.335 ;
        RECT 45.690 180.150 46.825 180.290 ;
        RECT 43.315 180.105 43.605 180.150 ;
        RECT 46.535 180.105 46.825 180.150 ;
        RECT 48.375 180.290 48.665 180.335 ;
        RECT 50.215 180.290 50.505 180.335 ;
        RECT 54.890 180.290 55.030 180.445 ;
        RECT 59.860 180.335 60.180 180.350 ;
        RECT 63.155 180.335 63.445 180.650 ;
        RECT 65.840 180.630 66.160 180.690 ;
        RECT 67.695 180.630 67.985 180.675 ;
        RECT 65.840 180.490 67.985 180.630 ;
        RECT 65.840 180.430 66.160 180.490 ;
        RECT 67.695 180.445 67.985 180.490 ;
        RECT 68.615 180.445 68.905 180.675 ;
        RECT 69.075 180.630 69.365 180.675 ;
        RECT 69.980 180.630 70.300 180.690 ;
        RECT 69.075 180.490 70.300 180.630 ;
        RECT 69.075 180.445 69.365 180.490 ;
        RECT 59.855 180.290 60.505 180.335 ;
        RECT 63.155 180.290 63.745 180.335 ;
        RECT 48.375 180.150 50.505 180.290 ;
        RECT 48.375 180.105 48.665 180.150 ;
        RECT 50.215 180.105 50.505 180.150 ;
        RECT 52.130 180.150 55.030 180.290 ;
        RECT 55.350 180.150 63.745 180.290 ;
        RECT 22.230 179.810 23.840 179.950 ;
        RECT 13.185 179.765 13.475 179.810 ;
        RECT 13.860 179.750 14.180 179.810 ;
        RECT 19.380 179.750 19.700 179.810 ;
        RECT 23.520 179.750 23.840 179.810 ;
        RECT 36.415 179.765 36.705 179.995 ;
        RECT 36.860 179.750 37.180 180.010 ;
        RECT 37.780 179.950 38.100 180.010 ;
        RECT 38.715 179.950 39.005 179.995 ;
        RECT 37.780 179.810 39.005 179.950 ;
        RECT 39.250 179.950 39.390 180.105 ;
        RECT 52.130 180.010 52.270 180.150 ;
        RECT 39.620 179.950 39.940 180.010 ;
        RECT 39.250 179.810 39.940 179.950 ;
        RECT 37.780 179.750 38.100 179.810 ;
        RECT 38.715 179.765 39.005 179.810 ;
        RECT 39.620 179.750 39.940 179.810 ;
        RECT 45.600 179.950 45.920 180.010 ;
        RECT 51.580 179.950 51.900 180.010 ;
        RECT 45.600 179.810 51.900 179.950 ;
        RECT 45.600 179.750 45.920 179.810 ;
        RECT 51.580 179.750 51.900 179.810 ;
        RECT 52.040 179.750 52.360 180.010 ;
        RECT 52.500 179.750 52.820 180.010 ;
        RECT 53.880 179.950 54.200 180.010 ;
        RECT 54.355 179.950 54.645 179.995 ;
        RECT 53.880 179.810 54.645 179.950 ;
        RECT 53.880 179.750 54.200 179.810 ;
        RECT 54.355 179.765 54.645 179.810 ;
        RECT 54.800 179.950 55.120 180.010 ;
        RECT 55.350 179.950 55.490 180.150 ;
        RECT 59.855 180.105 60.505 180.150 ;
        RECT 63.455 180.105 63.745 180.150 ;
        RECT 59.860 180.090 60.180 180.105 ;
        RECT 54.800 179.810 55.490 179.950 ;
        RECT 56.180 179.950 56.500 180.010 ;
        RECT 68.690 179.950 68.830 180.445 ;
        RECT 69.980 180.430 70.300 180.490 ;
        RECT 70.900 180.430 71.220 180.690 ;
        RECT 71.825 180.630 72.115 180.675 ;
        RECT 75.040 180.630 75.360 180.690 ;
        RECT 71.825 180.490 75.360 180.630 ;
        RECT 71.825 180.445 72.115 180.490 ;
        RECT 75.040 180.430 75.360 180.490 ;
        RECT 78.260 180.430 78.580 180.690 ;
        RECT 84.700 180.430 85.020 180.690 ;
        RECT 85.250 180.675 85.390 180.830 ;
        RECT 85.620 180.830 90.065 180.970 ;
        RECT 85.620 180.770 85.940 180.830 ;
        RECT 89.775 180.785 90.065 180.830 ;
        RECT 93.440 180.770 93.760 181.030 ;
        RECT 94.820 180.970 95.140 181.030 ;
        RECT 110.000 180.970 110.320 181.030 ;
        RECT 127.570 180.970 127.710 181.170 ;
        RECT 129.410 180.970 129.550 181.510 ;
        RECT 137.140 181.450 137.460 181.710 ;
        RECT 152.780 181.450 153.100 181.710 ;
        RECT 139.915 180.970 140.205 181.015 ;
        RECT 141.280 180.970 141.600 181.030 ;
        RECT 143.120 180.970 143.440 181.030 ;
        RECT 152.870 180.970 153.010 181.450 ;
        RECT 94.820 180.830 110.320 180.970 ;
        RECT 94.820 180.770 95.140 180.830 ;
        RECT 110.000 180.770 110.320 180.830 ;
        RECT 110.550 180.830 121.270 180.970 ;
        RECT 85.175 180.445 85.465 180.675 ;
        RECT 87.935 180.445 88.225 180.675 ;
        RECT 88.380 180.630 88.700 180.690 ;
        RECT 88.855 180.630 89.145 180.675 ;
        RECT 88.380 180.490 89.145 180.630 ;
        RECT 72.280 180.290 72.600 180.350 ;
        RECT 75.960 180.290 76.280 180.350 ;
        RECT 72.280 180.150 76.280 180.290 ;
        RECT 72.280 180.090 72.600 180.150 ;
        RECT 75.960 180.090 76.280 180.150 ;
        RECT 77.340 180.290 77.660 180.350 ;
        RECT 78.350 180.290 78.490 180.430 ;
        RECT 88.010 180.290 88.150 180.445 ;
        RECT 88.380 180.430 88.700 180.490 ;
        RECT 88.855 180.445 89.145 180.490 ;
        RECT 91.140 180.430 91.460 180.690 ;
        RECT 96.660 180.430 96.980 180.690 ;
        RECT 97.120 180.630 97.440 180.690 ;
        RECT 97.595 180.630 97.885 180.675 ;
        RECT 108.160 180.630 108.480 180.690 ;
        RECT 110.550 180.675 110.690 180.830 ;
        RECT 110.475 180.630 110.765 180.675 ;
        RECT 97.120 180.490 97.885 180.630 ;
        RECT 97.120 180.430 97.440 180.490 ;
        RECT 97.595 180.445 97.885 180.490 ;
        RECT 104.570 180.490 110.765 180.630 ;
        RECT 77.340 180.150 88.150 180.290 ;
        RECT 77.340 180.090 77.660 180.150 ;
        RECT 69.060 179.950 69.380 180.010 ;
        RECT 56.180 179.810 69.380 179.950 ;
        RECT 54.800 179.750 55.120 179.810 ;
        RECT 56.180 179.750 56.500 179.810 ;
        RECT 69.060 179.750 69.380 179.810 ;
        RECT 70.440 179.950 70.760 180.010 ;
        RECT 70.915 179.950 71.205 179.995 ;
        RECT 70.440 179.810 71.205 179.950 ;
        RECT 70.440 179.750 70.760 179.810 ;
        RECT 70.915 179.765 71.205 179.810 ;
        RECT 71.820 179.750 72.140 180.010 ;
        RECT 78.260 179.750 78.580 180.010 ;
        RECT 88.010 179.950 88.150 180.150 ;
        RECT 100.800 180.090 101.120 180.350 ;
        RECT 103.955 180.290 104.245 180.335 ;
        RECT 104.570 180.290 104.710 180.490 ;
        RECT 108.160 180.430 108.480 180.490 ;
        RECT 110.475 180.445 110.765 180.490 ;
        RECT 112.575 180.630 112.865 180.675 ;
        RECT 113.220 180.630 113.540 180.690 ;
        RECT 112.575 180.490 113.540 180.630 ;
        RECT 112.575 180.445 112.865 180.490 ;
        RECT 113.220 180.430 113.540 180.490 ;
        RECT 114.155 180.630 114.445 180.675 ;
        RECT 114.600 180.630 114.920 180.690 ;
        RECT 114.155 180.490 114.920 180.630 ;
        RECT 114.155 180.445 114.445 180.490 ;
        RECT 114.600 180.430 114.920 180.490 ;
        RECT 115.150 180.490 117.130 180.630 ;
        RECT 103.955 180.150 104.710 180.290 ;
        RECT 103.955 180.105 104.245 180.150 ;
        RECT 104.940 180.090 105.260 180.350 ;
        RECT 107.700 180.290 108.020 180.350 ;
        RECT 111.395 180.290 111.685 180.335 ;
        RECT 107.700 180.150 111.685 180.290 ;
        RECT 107.700 180.090 108.020 180.150 ;
        RECT 111.395 180.105 111.685 180.150 ;
        RECT 111.855 180.290 112.145 180.335 ;
        RECT 113.680 180.290 114.000 180.350 ;
        RECT 111.855 180.150 114.000 180.290 ;
        RECT 111.855 180.105 112.145 180.150 ;
        RECT 92.520 179.950 92.840 180.010 ;
        RECT 88.010 179.810 92.840 179.950 ;
        RECT 100.890 179.950 101.030 180.090 ;
        RECT 104.480 179.950 104.800 180.010 ;
        RECT 100.890 179.810 104.800 179.950 ;
        RECT 111.470 179.950 111.610 180.105 ;
        RECT 113.680 180.090 114.000 180.150 ;
        RECT 115.150 179.950 115.290 180.490 ;
        RECT 115.980 180.290 116.300 180.350 ;
        RECT 116.455 180.290 116.745 180.335 ;
        RECT 115.980 180.150 116.745 180.290 ;
        RECT 116.990 180.290 117.130 180.490 ;
        RECT 119.200 180.430 119.520 180.690 ;
        RECT 121.130 180.675 121.270 180.830 ;
        RECT 122.970 180.830 127.250 180.970 ;
        RECT 127.570 180.830 129.090 180.970 ;
        RECT 129.410 180.830 143.440 180.970 ;
        RECT 122.970 180.675 123.110 180.830 ;
        RECT 127.110 180.690 127.250 180.830 ;
        RECT 121.055 180.630 121.345 180.675 ;
        RECT 122.895 180.630 123.185 180.675 ;
        RECT 121.055 180.490 123.185 180.630 ;
        RECT 121.055 180.445 121.345 180.490 ;
        RECT 122.895 180.445 123.185 180.490 ;
        RECT 123.800 180.630 124.120 180.690 ;
        RECT 124.275 180.630 124.565 180.675 ;
        RECT 123.800 180.490 124.565 180.630 ;
        RECT 123.800 180.430 124.120 180.490 ;
        RECT 124.275 180.445 124.565 180.490 ;
        RECT 127.020 180.430 127.340 180.690 ;
        RECT 128.950 180.675 129.090 180.830 ;
        RECT 139.915 180.785 140.205 180.830 ;
        RECT 141.280 180.770 141.600 180.830 ;
        RECT 143.120 180.770 143.440 180.830 ;
        RECT 144.820 180.830 153.010 180.970 ;
        RECT 127.955 180.630 128.245 180.675 ;
        RECT 127.570 180.490 128.245 180.630 ;
        RECT 120.595 180.290 120.885 180.335 ;
        RECT 116.990 180.150 120.885 180.290 ;
        RECT 115.980 180.090 116.300 180.150 ;
        RECT 116.455 180.105 116.745 180.150 ;
        RECT 120.595 180.105 120.885 180.150 ;
        RECT 121.960 180.290 122.280 180.350 ;
        RECT 125.195 180.290 125.485 180.335 ;
        RECT 126.100 180.290 126.420 180.350 ;
        RECT 121.960 180.150 126.420 180.290 ;
        RECT 111.470 179.810 115.290 179.950 ;
        RECT 115.535 179.950 115.825 179.995 ;
        RECT 117.820 179.950 118.140 180.010 ;
        RECT 120.120 179.950 120.440 180.010 ;
        RECT 115.535 179.810 120.440 179.950 ;
        RECT 120.670 179.950 120.810 180.105 ;
        RECT 121.960 180.090 122.280 180.150 ;
        RECT 125.195 180.105 125.485 180.150 ;
        RECT 126.100 180.090 126.420 180.150 ;
        RECT 123.355 179.950 123.645 179.995 ;
        RECT 124.260 179.950 124.580 180.010 ;
        RECT 127.570 179.950 127.710 180.490 ;
        RECT 127.955 180.445 128.245 180.490 ;
        RECT 128.875 180.630 129.165 180.675 ;
        RECT 144.820 180.630 144.960 180.830 ;
        RECT 128.875 180.490 144.960 180.630 ;
        RECT 128.875 180.445 129.165 180.490 ;
        RECT 150.940 180.430 151.260 180.690 ;
        RECT 151.860 180.630 152.180 180.690 ;
        RECT 152.335 180.630 152.625 180.675 ;
        RECT 151.860 180.490 152.625 180.630 ;
        RECT 151.860 180.430 152.180 180.490 ;
        RECT 152.335 180.445 152.625 180.490 ;
        RECT 132.540 180.090 132.860 180.350 ;
        RECT 133.460 180.290 133.780 180.350 ;
        RECT 138.995 180.290 139.285 180.335 ;
        RECT 141.740 180.290 142.060 180.350 ;
        RECT 133.460 180.150 142.060 180.290 ;
        RECT 133.460 180.090 133.780 180.150 ;
        RECT 138.995 180.105 139.285 180.150 ;
        RECT 141.740 180.090 142.060 180.150 ;
        RECT 120.670 179.810 127.710 179.950 ;
        RECT 132.630 179.950 132.770 180.090 ;
        RECT 135.300 179.950 135.620 180.010 ;
        RECT 139.455 179.950 139.745 179.995 ;
        RECT 132.630 179.810 139.745 179.950 ;
        RECT 92.520 179.750 92.840 179.810 ;
        RECT 104.480 179.750 104.800 179.810 ;
        RECT 115.535 179.765 115.825 179.810 ;
        RECT 117.820 179.750 118.140 179.810 ;
        RECT 120.120 179.750 120.440 179.810 ;
        RECT 123.355 179.765 123.645 179.810 ;
        RECT 124.260 179.750 124.580 179.810 ;
        RECT 135.300 179.750 135.620 179.810 ;
        RECT 139.455 179.765 139.745 179.810 ;
        RECT 2.750 179.130 159.030 179.610 ;
        RECT 6.040 178.730 6.360 178.990 ;
        RECT 9.275 178.745 9.565 178.975 ;
        RECT 11.115 178.745 11.405 178.975 ;
        RECT 14.320 178.930 14.640 178.990 ;
        RECT 15.255 178.930 15.545 178.975 ;
        RECT 14.320 178.790 15.545 178.930 ;
        RECT 6.975 178.250 7.265 178.295 ;
        RECT 9.350 178.250 9.490 178.745 ;
        RECT 11.190 178.590 11.330 178.745 ;
        RECT 14.320 178.730 14.640 178.790 ;
        RECT 15.255 178.745 15.545 178.790 ;
        RECT 17.080 178.730 17.400 178.990 ;
        RECT 27.660 178.930 27.980 178.990 ;
        RECT 19.470 178.790 27.980 178.930 ;
        RECT 13.860 178.590 14.180 178.650 ;
        RECT 11.190 178.450 14.180 178.590 ;
        RECT 13.860 178.390 14.180 178.450 ;
        RECT 15.330 178.450 17.770 178.590 ;
        RECT 6.975 178.110 9.490 178.250 ;
        RECT 10.640 178.250 10.960 178.310 ;
        RECT 11.575 178.250 11.865 178.295 ;
        RECT 14.780 178.250 15.100 178.310 ;
        RECT 15.330 178.250 15.470 178.450 ;
        RECT 17.630 178.295 17.770 178.450 ;
        RECT 19.470 178.295 19.610 178.790 ;
        RECT 27.660 178.730 27.980 178.790 ;
        RECT 29.040 178.930 29.360 178.990 ;
        RECT 29.975 178.930 30.265 178.975 ;
        RECT 41.920 178.930 42.240 178.990 ;
        RECT 29.040 178.790 30.265 178.930 ;
        RECT 29.040 178.730 29.360 178.790 ;
        RECT 29.975 178.745 30.265 178.790 ;
        RECT 30.415 178.790 42.240 178.930 ;
        RECT 23.520 178.635 23.840 178.650 ;
        RECT 23.055 178.590 23.840 178.635 ;
        RECT 26.655 178.590 26.945 178.635 ;
        RECT 23.055 178.450 26.945 178.590 ;
        RECT 23.055 178.405 23.840 178.450 ;
        RECT 23.520 178.390 23.840 178.405 ;
        RECT 26.355 178.405 26.945 178.450 ;
        RECT 10.640 178.110 15.470 178.250 ;
        RECT 6.975 178.065 7.265 178.110 ;
        RECT 10.640 178.050 10.960 178.110 ;
        RECT 11.575 178.065 11.865 178.110 ;
        RECT 14.780 178.050 15.100 178.110 ;
        RECT 17.555 178.065 17.845 178.295 ;
        RECT 19.395 178.065 19.685 178.295 ;
        RECT 19.860 178.250 20.150 178.295 ;
        RECT 21.695 178.250 21.985 178.295 ;
        RECT 25.275 178.250 25.565 178.295 ;
        RECT 19.860 178.110 25.565 178.250 ;
        RECT 19.860 178.065 20.150 178.110 ;
        RECT 21.695 178.065 21.985 178.110 ;
        RECT 25.275 178.065 25.565 178.110 ;
        RECT 26.355 178.090 26.645 178.405 ;
        RECT 12.495 177.910 12.785 177.955 ;
        RECT 13.400 177.910 13.720 177.970 ;
        RECT 12.495 177.770 13.720 177.910 ;
        RECT 12.495 177.725 12.785 177.770 ;
        RECT 13.400 177.710 13.720 177.770 ;
        RECT 18.460 177.710 18.780 177.970 ;
        RECT 4.660 177.570 4.980 177.630 ;
        RECT 19.470 177.570 19.610 178.065 ;
        RECT 20.760 177.710 21.080 177.970 ;
        RECT 28.120 177.910 28.440 177.970 ;
        RECT 30.415 177.910 30.555 178.790 ;
        RECT 41.920 178.730 42.240 178.790 ;
        RECT 46.455 178.930 46.745 178.975 ;
        RECT 48.820 178.930 49.140 178.990 ;
        RECT 52.040 178.930 52.360 178.990 ;
        RECT 46.455 178.790 52.360 178.930 ;
        RECT 46.455 178.745 46.745 178.790 ;
        RECT 48.820 178.730 49.140 178.790 ;
        RECT 52.040 178.730 52.360 178.790 ;
        RECT 53.420 178.730 53.740 178.990 ;
        RECT 57.575 178.930 57.865 178.975 ;
        RECT 61.700 178.930 62.020 178.990 ;
        RECT 57.575 178.790 62.020 178.930 ;
        RECT 57.575 178.745 57.865 178.790 ;
        RECT 61.700 178.730 62.020 178.790 ;
        RECT 71.830 178.930 72.120 178.975 ;
        RECT 78.270 178.930 78.560 178.975 ;
        RECT 94.820 178.930 95.140 178.990 ;
        RECT 102.640 178.930 102.960 178.990 ;
        RECT 105.860 178.930 106.180 178.990 ;
        RECT 71.830 178.790 78.560 178.930 ;
        RECT 71.830 178.745 72.120 178.790 ;
        RECT 78.270 178.745 78.560 178.790 ;
        RECT 78.810 178.790 92.750 178.930 ;
        RECT 34.560 178.590 34.880 178.650 ;
        RECT 36.395 178.590 37.045 178.635 ;
        RECT 39.995 178.590 40.285 178.635 ;
        RECT 34.560 178.450 40.285 178.590 ;
        RECT 34.560 178.390 34.880 178.450 ;
        RECT 36.395 178.405 37.045 178.450 ;
        RECT 39.695 178.405 40.285 178.450 ;
        RECT 43.315 178.590 43.605 178.635 ;
        RECT 43.760 178.590 44.080 178.650 ;
        RECT 43.315 178.450 44.080 178.590 ;
        RECT 43.315 178.405 43.605 178.450 ;
        RECT 30.895 178.065 31.185 178.295 ;
        RECT 28.120 177.770 30.555 177.910 ;
        RECT 28.120 177.710 28.440 177.770 ;
        RECT 4.660 177.430 19.610 177.570 ;
        RECT 20.265 177.570 20.555 177.615 ;
        RECT 22.155 177.570 22.445 177.615 ;
        RECT 25.275 177.570 25.565 177.615 ;
        RECT 20.265 177.430 25.565 177.570 ;
        RECT 4.660 177.370 4.980 177.430 ;
        RECT 20.265 177.385 20.555 177.430 ;
        RECT 22.155 177.385 22.445 177.430 ;
        RECT 25.275 177.385 25.565 177.430 ;
        RECT 30.970 177.230 31.110 178.065 ;
        RECT 31.340 178.050 31.660 178.310 ;
        RECT 31.800 178.250 32.120 178.310 ;
        RECT 32.735 178.250 33.025 178.295 ;
        RECT 31.800 178.110 33.025 178.250 ;
        RECT 31.800 178.050 32.120 178.110 ;
        RECT 32.735 178.065 33.025 178.110 ;
        RECT 33.200 178.250 33.490 178.295 ;
        RECT 35.035 178.250 35.325 178.295 ;
        RECT 38.615 178.250 38.905 178.295 ;
        RECT 33.200 178.110 38.905 178.250 ;
        RECT 33.200 178.065 33.490 178.110 ;
        RECT 35.035 178.065 35.325 178.110 ;
        RECT 38.615 178.065 38.905 178.110 ;
        RECT 39.695 178.090 39.985 178.405 ;
        RECT 43.760 178.390 44.080 178.450 ;
        RECT 44.235 178.590 44.525 178.635 ;
        RECT 45.600 178.590 45.920 178.650 ;
        RECT 44.235 178.450 45.920 178.590 ;
        RECT 44.235 178.405 44.525 178.450 ;
        RECT 45.600 178.390 45.920 178.450 ;
        RECT 47.440 178.390 47.760 178.650 ;
        RECT 49.295 178.590 49.585 178.635 ;
        RECT 52.500 178.590 52.820 178.650 ;
        RECT 53.510 178.590 53.650 178.730 ;
        RECT 60.320 178.590 60.640 178.650 ;
        RECT 49.295 178.450 52.820 178.590 ;
        RECT 49.295 178.405 49.585 178.450 ;
        RECT 52.500 178.390 52.820 178.450 ;
        RECT 53.075 178.450 53.650 178.590 ;
        RECT 56.730 178.450 60.640 178.590 ;
        RECT 41.935 178.065 42.225 178.295 ;
        RECT 34.115 177.910 34.405 177.955 ;
        RECT 32.350 177.770 34.405 177.910 ;
        RECT 32.350 177.615 32.490 177.770 ;
        RECT 34.115 177.725 34.405 177.770 ;
        RECT 32.275 177.385 32.565 177.615 ;
        RECT 33.605 177.570 33.895 177.615 ;
        RECT 35.495 177.570 35.785 177.615 ;
        RECT 38.615 177.570 38.905 177.615 ;
        RECT 33.605 177.430 38.905 177.570 ;
        RECT 42.010 177.570 42.150 178.065 ;
        RECT 42.840 178.050 43.160 178.310 ;
        RECT 45.140 178.050 45.460 178.310 ;
        RECT 47.900 178.050 48.220 178.310 ;
        RECT 50.200 178.295 50.520 178.310 ;
        RECT 48.605 178.065 48.895 178.295 ;
        RECT 49.755 178.065 50.045 178.295 ;
        RECT 50.200 178.250 50.530 178.295 ;
        RECT 51.120 178.250 51.440 178.310 ;
        RECT 52.055 178.250 52.345 178.295 ;
        RECT 50.200 178.110 50.715 178.250 ;
        RECT 51.120 178.110 52.345 178.250 ;
        RECT 50.200 178.065 50.530 178.110 ;
        RECT 42.395 177.910 42.685 177.955 ;
        RECT 42.395 177.770 48.165 177.910 ;
        RECT 42.395 177.725 42.685 177.770 ;
        RECT 43.300 177.570 43.620 177.630 ;
        RECT 45.140 177.570 45.460 177.630 ;
        RECT 42.010 177.430 45.460 177.570 ;
        RECT 33.605 177.385 33.895 177.430 ;
        RECT 35.495 177.385 35.785 177.430 ;
        RECT 38.615 177.385 38.905 177.430 ;
        RECT 43.300 177.370 43.620 177.430 ;
        RECT 45.140 177.370 45.460 177.430 ;
        RECT 45.615 177.570 45.905 177.615 ;
        RECT 46.060 177.570 46.380 177.630 ;
        RECT 45.615 177.430 46.380 177.570 ;
        RECT 48.025 177.570 48.165 177.770 ;
        RECT 48.680 177.570 48.820 178.065 ;
        RECT 49.830 177.910 49.970 178.065 ;
        RECT 50.200 178.050 50.520 178.065 ;
        RECT 51.120 178.050 51.440 178.110 ;
        RECT 52.055 178.065 52.345 178.110 ;
        RECT 50.660 177.910 50.980 177.970 ;
        RECT 49.830 177.770 50.980 177.910 ;
        RECT 50.660 177.710 50.980 177.770 ;
        RECT 53.075 177.570 53.215 178.450 ;
        RECT 56.730 178.310 56.870 178.450 ;
        RECT 60.320 178.390 60.640 178.450 ;
        RECT 61.240 178.590 61.560 178.650 ;
        RECT 62.155 178.590 62.805 178.635 ;
        RECT 65.755 178.590 66.045 178.635 ;
        RECT 61.240 178.450 66.045 178.590 ;
        RECT 61.240 178.390 61.560 178.450 ;
        RECT 62.155 178.405 62.805 178.450 ;
        RECT 65.455 178.405 66.045 178.450 ;
        RECT 67.220 178.590 67.540 178.650 ;
        RECT 68.615 178.590 68.905 178.635 ;
        RECT 67.220 178.450 68.905 178.590 ;
        RECT 53.420 178.250 53.740 178.310 ;
        RECT 55.275 178.250 55.565 178.295 ;
        RECT 53.420 178.110 55.565 178.250 ;
        RECT 53.420 178.050 53.740 178.110 ;
        RECT 55.275 178.065 55.565 178.110 ;
        RECT 56.180 178.050 56.500 178.310 ;
        RECT 56.640 178.050 56.960 178.310 ;
        RECT 58.960 178.250 59.250 178.295 ;
        RECT 60.795 178.250 61.085 178.295 ;
        RECT 64.375 178.250 64.665 178.295 ;
        RECT 58.960 178.110 64.665 178.250 ;
        RECT 58.960 178.065 59.250 178.110 ;
        RECT 60.795 178.065 61.085 178.110 ;
        RECT 64.375 178.065 64.665 178.110 ;
        RECT 65.455 178.090 65.745 178.405 ;
        RECT 67.220 178.390 67.540 178.450 ;
        RECT 68.615 178.405 68.905 178.450 ;
        RECT 77.800 178.590 78.120 178.650 ;
        RECT 78.810 178.590 78.950 178.790 ;
        RECT 77.800 178.450 78.950 178.590 ;
        RECT 83.335 178.590 83.625 178.635 ;
        RECT 84.240 178.590 84.560 178.650 ;
        RECT 83.335 178.450 84.560 178.590 ;
        RECT 77.800 178.390 78.120 178.450 ;
        RECT 83.335 178.405 83.625 178.450 ;
        RECT 84.240 178.390 84.560 178.450 ;
        RECT 85.160 178.635 85.480 178.650 ;
        RECT 85.160 178.405 85.695 178.635 ;
        RECT 90.220 178.590 90.540 178.650 ;
        RECT 86.630 178.450 90.910 178.590 ;
        RECT 85.160 178.390 85.480 178.405 ;
        RECT 67.680 178.250 68.000 178.310 ;
        RECT 71.820 178.250 72.140 178.310 ;
        RECT 73.215 178.250 73.505 178.295 ;
        RECT 67.680 178.110 69.290 178.250 ;
        RECT 67.680 178.050 68.000 178.110 ;
        RECT 57.560 177.910 57.880 177.970 ;
        RECT 58.495 177.910 58.785 177.955 ;
        RECT 57.560 177.770 58.785 177.910 ;
        RECT 57.560 177.710 57.880 177.770 ;
        RECT 58.495 177.725 58.785 177.770 ;
        RECT 48.025 177.430 48.820 177.570 ;
        RECT 50.755 177.430 57.790 177.570 ;
        RECT 45.615 177.385 45.905 177.430 ;
        RECT 36.860 177.230 37.180 177.290 ;
        RECT 30.970 177.090 37.180 177.230 ;
        RECT 36.860 177.030 37.180 177.090 ;
        RECT 41.460 177.230 41.780 177.290 ;
        RECT 42.380 177.230 42.700 177.290 ;
        RECT 41.460 177.090 42.700 177.230 ;
        RECT 41.460 177.030 41.780 177.090 ;
        RECT 42.380 177.030 42.700 177.090 ;
        RECT 42.840 177.230 43.160 177.290 ;
        RECT 45.690 177.230 45.830 177.385 ;
        RECT 46.060 177.370 46.380 177.430 ;
        RECT 42.840 177.090 45.830 177.230 ;
        RECT 46.535 177.230 46.825 177.275 ;
        RECT 50.755 177.230 50.895 177.430 ;
        RECT 57.650 177.290 57.790 177.430 ;
        RECT 46.535 177.090 50.895 177.230 ;
        RECT 42.840 177.030 43.160 177.090 ;
        RECT 46.535 177.045 46.825 177.090 ;
        RECT 51.120 177.030 51.440 177.290 ;
        RECT 52.500 177.030 52.820 177.290 ;
        RECT 56.655 177.230 56.945 177.275 ;
        RECT 57.100 177.230 57.420 177.290 ;
        RECT 56.655 177.090 57.420 177.230 ;
        RECT 56.655 177.045 56.945 177.090 ;
        RECT 57.100 177.030 57.420 177.090 ;
        RECT 57.560 177.030 57.880 177.290 ;
        RECT 58.570 177.230 58.710 177.725 ;
        RECT 59.860 177.710 60.180 177.970 ;
        RECT 60.320 177.910 60.640 177.970 ;
        RECT 69.150 177.910 69.290 178.110 ;
        RECT 71.820 178.110 73.505 178.250 ;
        RECT 71.820 178.050 72.140 178.110 ;
        RECT 73.215 178.065 73.505 178.110 ;
        RECT 75.040 178.050 75.360 178.310 ;
        RECT 75.500 178.250 75.820 178.310 ;
        RECT 75.975 178.250 76.265 178.295 ;
        RECT 76.880 178.250 77.200 178.310 ;
        RECT 75.500 178.110 77.200 178.250 ;
        RECT 75.500 178.050 75.820 178.110 ;
        RECT 75.975 178.065 76.265 178.110 ;
        RECT 76.880 178.050 77.200 178.110 ;
        RECT 77.340 178.050 77.660 178.310 ;
        RECT 79.180 178.250 79.500 178.310 ;
        RECT 81.495 178.250 81.785 178.295 ;
        RECT 79.180 178.110 81.785 178.250 ;
        RECT 79.180 178.050 79.500 178.110 ;
        RECT 81.495 178.065 81.785 178.110 ;
        RECT 81.955 178.065 82.245 178.295 ;
        RECT 82.860 178.250 83.180 178.310 ;
        RECT 86.630 178.295 86.770 178.450 ;
        RECT 90.220 178.390 90.540 178.450 ;
        RECT 84.715 178.250 85.005 178.295 ;
        RECT 82.860 178.110 85.005 178.250 ;
        RECT 81.020 177.910 81.340 177.970 ;
        RECT 60.320 177.770 65.610 177.910 ;
        RECT 69.150 177.770 81.340 177.910 ;
        RECT 82.030 177.910 82.170 178.065 ;
        RECT 82.860 178.050 83.180 178.110 ;
        RECT 84.715 178.065 85.005 178.110 ;
        RECT 86.095 178.065 86.385 178.295 ;
        RECT 86.555 178.065 86.845 178.295 ;
        RECT 82.030 177.770 83.550 177.910 ;
        RECT 60.320 177.710 60.640 177.770 ;
        RECT 59.365 177.570 59.655 177.615 ;
        RECT 61.255 177.570 61.545 177.615 ;
        RECT 64.375 177.570 64.665 177.615 ;
        RECT 59.365 177.430 64.665 177.570 ;
        RECT 59.365 177.385 59.655 177.430 ;
        RECT 61.255 177.385 61.545 177.430 ;
        RECT 64.375 177.385 64.665 177.430 ;
        RECT 64.920 177.370 65.240 177.630 ;
        RECT 65.470 177.570 65.610 177.770 ;
        RECT 81.020 177.710 81.340 177.770 ;
        RECT 83.410 177.630 83.550 177.770 ;
        RECT 83.780 177.710 84.100 177.970 ;
        RECT 69.980 177.570 70.300 177.630 ;
        RECT 65.470 177.430 70.300 177.570 ;
        RECT 69.980 177.370 70.300 177.430 ;
        RECT 74.580 177.570 74.900 177.630 ;
        RECT 75.515 177.570 75.805 177.615 ;
        RECT 74.580 177.430 75.805 177.570 ;
        RECT 74.580 177.370 74.900 177.430 ;
        RECT 75.515 177.385 75.805 177.430 ;
        RECT 78.720 177.570 79.040 177.630 ;
        RECT 78.720 177.430 83.090 177.570 ;
        RECT 78.720 177.370 79.040 177.430 ;
        RECT 59.860 177.230 60.180 177.290 ;
        RECT 58.570 177.090 60.180 177.230 ;
        RECT 65.010 177.230 65.150 177.370 ;
        RECT 80.575 177.230 80.865 177.275 ;
        RECT 65.010 177.090 80.865 177.230 ;
        RECT 82.950 177.230 83.090 177.430 ;
        RECT 83.320 177.370 83.640 177.630 ;
        RECT 86.170 177.570 86.310 178.065 ;
        RECT 87.000 178.050 87.320 178.310 ;
        RECT 89.760 178.250 90.080 178.310 ;
        RECT 90.770 178.295 90.910 178.450 ;
        RECT 87.550 178.110 90.080 178.250 ;
        RECT 87.550 177.570 87.690 178.110 ;
        RECT 89.760 178.050 90.080 178.110 ;
        RECT 90.695 178.065 90.985 178.295 ;
        RECT 91.155 178.065 91.445 178.295 ;
        RECT 91.615 178.250 91.905 178.295 ;
        RECT 92.610 178.250 92.750 178.790 ;
        RECT 93.530 178.790 95.140 178.930 ;
        RECT 93.530 178.635 93.670 178.790 ;
        RECT 94.820 178.730 95.140 178.790 ;
        RECT 98.590 178.790 106.180 178.930 ;
        RECT 93.455 178.405 93.745 178.635 ;
        RECT 98.590 178.590 98.730 178.790 ;
        RECT 102.640 178.730 102.960 178.790 ;
        RECT 105.860 178.730 106.180 178.790 ;
        RECT 108.160 178.730 108.480 178.990 ;
        RECT 109.080 178.730 109.400 178.990 ;
        RECT 110.920 178.730 111.240 178.990 ;
        RECT 119.215 178.930 119.505 178.975 ;
        RECT 121.055 178.930 121.345 178.975 ;
        RECT 124.720 178.930 125.040 178.990 ;
        RECT 119.215 178.790 120.810 178.930 ;
        RECT 119.215 178.745 119.505 178.790 ;
        RECT 104.020 178.590 104.340 178.650 ;
        RECT 94.450 178.450 98.730 178.590 ;
        RECT 91.615 178.110 92.750 178.250 ;
        RECT 91.615 178.065 91.905 178.110 ;
        RECT 87.920 177.710 88.240 177.970 ;
        RECT 90.770 177.910 90.910 178.065 ;
        RECT 88.470 177.770 90.910 177.910 ;
        RECT 86.170 177.430 87.690 177.570 ;
        RECT 88.470 177.230 88.610 177.770 ;
        RECT 89.760 177.570 90.080 177.630 ;
        RECT 91.230 177.570 91.370 178.065 ;
        RECT 94.450 177.910 94.590 178.450 ;
        RECT 96.675 178.250 96.965 178.295 ;
        RECT 98.040 178.250 98.360 178.310 ;
        RECT 98.590 178.295 98.730 178.450 ;
        RECT 99.510 178.450 107.010 178.590 ;
        RECT 99.510 178.295 99.650 178.450 ;
        RECT 104.020 178.390 104.340 178.450 ;
        RECT 91.690 177.770 94.590 177.910 ;
        RECT 94.910 178.110 98.360 178.250 ;
        RECT 91.690 177.630 91.830 177.770 ;
        RECT 89.760 177.430 91.370 177.570 ;
        RECT 89.760 177.370 90.080 177.430 ;
        RECT 82.950 177.090 88.610 177.230 ;
        RECT 88.855 177.230 89.145 177.275 ;
        RECT 89.300 177.230 89.620 177.290 ;
        RECT 88.855 177.090 89.620 177.230 ;
        RECT 91.230 177.230 91.370 177.430 ;
        RECT 91.600 177.370 91.920 177.630 ;
        RECT 92.520 177.370 92.840 177.630 ;
        RECT 94.910 177.230 95.050 178.110 ;
        RECT 96.675 178.065 96.965 178.110 ;
        RECT 98.040 178.050 98.360 178.110 ;
        RECT 98.515 178.065 98.805 178.295 ;
        RECT 99.435 178.065 99.725 178.295 ;
        RECT 99.895 178.065 100.185 178.295 ;
        RECT 96.200 177.710 96.520 177.970 ;
        RECT 99.970 177.570 100.110 178.065 ;
        RECT 101.260 178.050 101.580 178.310 ;
        RECT 102.180 178.250 102.500 178.310 ;
        RECT 102.180 178.110 102.870 178.250 ;
        RECT 102.180 178.050 102.500 178.110 ;
        RECT 95.370 177.430 100.110 177.570 ;
        RECT 100.355 177.570 100.645 177.615 ;
        RECT 100.800 177.570 101.120 177.630 ;
        RECT 100.355 177.430 101.120 177.570 ;
        RECT 95.370 177.290 95.510 177.430 ;
        RECT 100.355 177.385 100.645 177.430 ;
        RECT 100.800 177.370 101.120 177.430 ;
        RECT 91.230 177.090 95.050 177.230 ;
        RECT 59.860 177.030 60.180 177.090 ;
        RECT 80.575 177.045 80.865 177.090 ;
        RECT 88.855 177.045 89.145 177.090 ;
        RECT 89.300 177.030 89.620 177.090 ;
        RECT 95.280 177.030 95.600 177.290 ;
        RECT 97.120 177.230 97.440 177.290 ;
        RECT 101.350 177.230 101.490 178.050 ;
        RECT 102.730 177.955 102.870 178.110 ;
        RECT 103.560 178.050 103.880 178.310 ;
        RECT 105.860 178.250 106.180 178.310 ;
        RECT 106.870 178.295 107.010 178.450 ;
        RECT 106.335 178.250 106.625 178.295 ;
        RECT 105.860 178.110 106.625 178.250 ;
        RECT 105.860 178.050 106.180 178.110 ;
        RECT 106.335 178.065 106.625 178.110 ;
        RECT 106.795 178.065 107.085 178.295 ;
        RECT 107.700 178.050 108.020 178.310 ;
        RECT 108.250 178.295 108.390 178.730 ;
        RECT 113.220 178.590 113.540 178.650 ;
        RECT 120.670 178.590 120.810 178.790 ;
        RECT 121.055 178.790 125.040 178.930 ;
        RECT 121.055 178.745 121.345 178.790 ;
        RECT 124.720 178.730 125.040 178.790 ;
        RECT 125.180 178.930 125.500 178.990 ;
        RECT 128.860 178.930 129.180 178.990 ;
        RECT 125.180 178.790 129.180 178.930 ;
        RECT 125.180 178.730 125.500 178.790 ;
        RECT 128.860 178.730 129.180 178.790 ;
        RECT 129.320 178.730 129.640 178.990 ;
        RECT 135.315 178.930 135.605 178.975 ;
        RECT 130.330 178.790 135.070 178.930 ;
        RECT 121.500 178.590 121.820 178.650 ;
        RECT 130.330 178.590 130.470 178.790 ;
        RECT 133.935 178.590 134.225 178.635 ;
        RECT 113.220 178.450 118.050 178.590 ;
        RECT 120.670 178.450 121.820 178.590 ;
        RECT 113.220 178.390 113.540 178.450 ;
        RECT 108.175 178.065 108.465 178.295 ;
        RECT 110.460 178.050 110.780 178.310 ;
        RECT 113.680 178.050 114.000 178.310 ;
        RECT 114.690 178.295 114.830 178.450 ;
        RECT 117.910 178.310 118.050 178.450 ;
        RECT 121.500 178.390 121.820 178.450 ;
        RECT 128.030 178.450 130.470 178.590 ;
        RECT 130.790 178.450 134.225 178.590 ;
        RECT 134.930 178.590 135.070 178.790 ;
        RECT 135.315 178.790 142.890 178.930 ;
        RECT 135.315 178.745 135.605 178.790 ;
        RECT 138.520 178.590 138.840 178.650 ;
        RECT 140.360 178.590 140.680 178.650 ;
        RECT 134.930 178.450 138.290 178.590 ;
        RECT 120.135 178.310 120.425 178.345 ;
        RECT 128.030 178.310 128.170 178.450 ;
        RECT 114.615 178.065 114.905 178.295 ;
        RECT 102.655 177.725 102.945 177.955 ;
        RECT 103.650 177.910 103.790 178.050 ;
        RECT 107.790 177.910 107.930 178.050 ;
        RECT 115.535 177.910 115.825 178.125 ;
        RECT 117.820 178.050 118.140 178.310 ;
        RECT 118.280 178.050 118.600 178.310 ;
        RECT 120.120 178.300 120.440 178.310 ;
        RECT 120.120 178.160 120.585 178.300 ;
        RECT 120.120 178.050 120.440 178.160 ;
        RECT 121.040 178.050 121.360 178.310 ;
        RECT 123.340 178.250 123.660 178.310 ;
        RECT 123.815 178.250 124.105 178.295 ;
        RECT 123.340 178.110 124.105 178.250 ;
        RECT 123.340 178.050 123.660 178.110 ;
        RECT 123.815 178.065 124.105 178.110 ;
        RECT 125.195 178.065 125.485 178.295 ;
        RECT 115.980 177.910 116.300 177.970 ;
        RECT 103.650 177.770 107.930 177.910 ;
        RECT 110.320 177.770 116.300 177.910 ;
        RECT 110.320 177.570 110.460 177.770 ;
        RECT 115.980 177.710 116.300 177.770 ;
        RECT 121.960 177.910 122.280 177.970 ;
        RECT 125.270 177.910 125.410 178.065 ;
        RECT 127.940 178.050 128.260 178.310 ;
        RECT 130.790 178.295 130.930 178.450 ;
        RECT 133.935 178.405 134.225 178.450 ;
        RECT 130.715 178.250 131.005 178.295 ;
        RECT 128.950 178.110 131.005 178.250 ;
        RECT 121.960 177.770 125.410 177.910 ;
        RECT 121.960 177.710 122.280 177.770 ;
        RECT 107.330 177.430 110.460 177.570 ;
        RECT 107.330 177.290 107.470 177.430 ;
        RECT 116.440 177.370 116.760 177.630 ;
        RECT 128.950 177.290 129.090 178.110 ;
        RECT 130.715 178.065 131.005 178.110 ;
        RECT 132.080 178.050 132.400 178.310 ;
        RECT 132.555 178.065 132.845 178.295 ;
        RECT 131.620 177.910 131.940 177.970 ;
        RECT 132.630 177.910 132.770 178.065 ;
        RECT 133.460 178.050 133.780 178.310 ;
        RECT 134.395 178.250 134.685 178.295 ;
        RECT 137.140 178.250 137.460 178.310 ;
        RECT 137.615 178.250 137.905 178.295 ;
        RECT 134.395 178.110 135.070 178.250 ;
        RECT 134.395 178.065 134.685 178.110 ;
        RECT 134.930 177.970 135.070 178.110 ;
        RECT 137.140 178.110 137.905 178.250 ;
        RECT 138.150 178.250 138.290 178.450 ;
        RECT 138.520 178.450 140.680 178.590 ;
        RECT 138.520 178.390 138.840 178.450 ;
        RECT 140.360 178.390 140.680 178.450 ;
        RECT 141.740 178.390 142.060 178.650 ;
        RECT 139.455 178.250 139.745 178.295 ;
        RECT 138.150 178.110 139.745 178.250 ;
        RECT 137.140 178.050 137.460 178.110 ;
        RECT 137.615 178.065 137.905 178.110 ;
        RECT 139.455 178.065 139.745 178.110 ;
        RECT 139.915 178.250 140.205 178.295 ;
        RECT 141.830 178.250 141.970 178.390 ;
        RECT 142.750 178.295 142.890 178.790 ;
        RECT 152.320 178.730 152.640 178.990 ;
        RECT 154.160 178.730 154.480 178.990 ;
        RECT 155.080 178.730 155.400 178.990 ;
        RECT 152.410 178.590 152.550 178.730 ;
        RECT 154.250 178.590 154.390 178.730 ;
        RECT 152.410 178.450 153.470 178.590 ;
        RECT 139.915 178.110 141.970 178.250 ;
        RECT 139.915 178.065 140.205 178.110 ;
        RECT 142.675 178.065 142.965 178.295 ;
        RECT 144.975 178.065 145.265 178.295 ;
        RECT 145.420 178.250 145.740 178.310 ;
        RECT 147.275 178.250 147.565 178.295 ;
        RECT 145.420 178.110 147.565 178.250 ;
        RECT 131.620 177.770 132.770 177.910 ;
        RECT 131.620 177.710 131.940 177.770 ;
        RECT 134.840 177.710 135.160 177.970 ;
        RECT 135.300 177.910 135.620 177.970 ;
        RECT 138.520 177.910 138.840 177.970 ;
        RECT 135.300 177.770 138.840 177.910 ;
        RECT 135.300 177.710 135.620 177.770 ;
        RECT 138.520 177.710 138.840 177.770 ;
        RECT 138.995 177.725 139.285 177.955 ;
        RECT 136.220 177.570 136.540 177.630 ;
        RECT 139.070 177.570 139.210 177.725 ;
        RECT 136.220 177.430 139.210 177.570 ;
        RECT 136.220 177.370 136.540 177.430 ;
        RECT 97.120 177.090 101.490 177.230 ;
        RECT 101.720 177.230 102.040 177.290 ;
        RECT 104.940 177.230 105.260 177.290 ;
        RECT 107.240 177.230 107.560 177.290 ;
        RECT 101.720 177.090 107.560 177.230 ;
        RECT 97.120 177.030 97.440 177.090 ;
        RECT 101.720 177.030 102.040 177.090 ;
        RECT 104.940 177.030 105.260 177.090 ;
        RECT 107.240 177.030 107.560 177.090 ;
        RECT 107.700 177.230 108.020 177.290 ;
        RECT 109.540 177.230 109.860 177.290 ;
        RECT 107.700 177.090 109.860 177.230 ;
        RECT 107.700 177.030 108.020 177.090 ;
        RECT 109.540 177.030 109.860 177.090 ;
        RECT 121.500 177.230 121.820 177.290 ;
        RECT 124.735 177.230 125.025 177.275 ;
        RECT 121.500 177.090 125.025 177.230 ;
        RECT 121.500 177.030 121.820 177.090 ;
        RECT 124.735 177.045 125.025 177.090 ;
        RECT 128.860 177.030 129.180 177.290 ;
        RECT 139.530 177.230 139.670 178.065 ;
        RECT 140.835 177.910 141.125 177.955 ;
        RECT 145.050 177.910 145.190 178.065 ;
        RECT 145.420 178.050 145.740 178.110 ;
        RECT 147.275 178.065 147.565 178.110 ;
        RECT 148.655 178.250 148.945 178.295 ;
        RECT 149.100 178.250 149.420 178.310 ;
        RECT 153.330 178.295 153.470 178.450 ;
        RECT 153.790 178.450 154.390 178.590 ;
        RECT 153.790 178.295 153.930 178.450 ;
        RECT 155.170 178.295 155.310 178.730 ;
        RECT 148.655 178.110 149.420 178.250 ;
        RECT 148.655 178.065 148.945 178.110 ;
        RECT 149.100 178.050 149.420 178.110 ;
        RECT 150.035 178.250 150.325 178.295 ;
        RECT 152.335 178.250 152.625 178.295 ;
        RECT 150.035 178.110 152.625 178.250 ;
        RECT 150.035 178.065 150.325 178.110 ;
        RECT 152.335 178.065 152.625 178.110 ;
        RECT 153.255 178.065 153.545 178.295 ;
        RECT 153.715 178.065 154.005 178.295 ;
        RECT 154.635 178.250 154.925 178.295 ;
        RECT 154.250 178.110 154.925 178.250 ;
        RECT 140.835 177.770 145.190 177.910 ;
        RECT 140.835 177.725 141.125 177.770 ;
        RECT 143.120 177.370 143.440 177.630 ;
        RECT 147.260 177.230 147.580 177.290 ;
        RECT 154.250 177.230 154.390 178.110 ;
        RECT 154.635 178.065 154.925 178.110 ;
        RECT 155.095 178.065 155.385 178.295 ;
        RECT 139.530 177.090 154.390 177.230 ;
        RECT 147.260 177.030 147.580 177.090 ;
        RECT 2.750 176.410 158.230 176.890 ;
        RECT 18.475 176.210 18.765 176.255 ;
        RECT 20.760 176.210 21.080 176.270 ;
        RECT 18.475 176.070 21.080 176.210 ;
        RECT 18.475 176.025 18.765 176.070 ;
        RECT 20.760 176.010 21.080 176.070 ;
        RECT 31.340 176.210 31.660 176.270 ;
        RECT 35.955 176.210 36.245 176.255 ;
        RECT 31.340 176.070 36.245 176.210 ;
        RECT 31.340 176.010 31.660 176.070 ;
        RECT 35.955 176.025 36.245 176.070 ;
        RECT 38.240 176.210 38.560 176.270 ;
        RECT 39.620 176.210 39.940 176.270 ;
        RECT 38.240 176.070 39.940 176.210 ;
        RECT 38.240 176.010 38.560 176.070 ;
        RECT 39.620 176.010 39.940 176.070 ;
        RECT 46.060 176.210 46.380 176.270 ;
        RECT 47.440 176.210 47.760 176.270 ;
        RECT 54.800 176.210 55.120 176.270 ;
        RECT 57.100 176.210 57.420 176.270 ;
        RECT 69.075 176.210 69.365 176.255 ;
        RECT 70.915 176.210 71.205 176.255 ;
        RECT 46.060 176.070 52.270 176.210 ;
        RECT 46.060 176.010 46.380 176.070 ;
        RECT 47.440 176.010 47.760 176.070 ;
        RECT 52.130 175.930 52.270 176.070 ;
        RECT 54.800 176.070 63.310 176.210 ;
        RECT 54.800 176.010 55.120 176.070 ;
        RECT 57.100 176.010 57.420 176.070 ;
        RECT 6.005 175.870 6.295 175.915 ;
        RECT 7.895 175.870 8.185 175.915 ;
        RECT 11.015 175.870 11.305 175.915 ;
        RECT 6.005 175.730 11.305 175.870 ;
        RECT 6.005 175.685 6.295 175.730 ;
        RECT 7.895 175.685 8.185 175.730 ;
        RECT 11.015 175.685 11.305 175.730 ;
        RECT 13.860 175.870 14.180 175.930 ;
        RECT 27.200 175.870 27.520 175.930 ;
        RECT 47.900 175.870 48.220 175.930 ;
        RECT 13.860 175.730 27.520 175.870 ;
        RECT 13.860 175.670 14.180 175.730 ;
        RECT 27.200 175.670 27.520 175.730 ;
        RECT 34.650 175.730 41.690 175.870 ;
        RECT 34.650 175.590 34.790 175.730 ;
        RECT 4.660 175.530 4.980 175.590 ;
        RECT 5.135 175.530 5.425 175.575 ;
        RECT 4.660 175.390 5.425 175.530 ;
        RECT 4.660 175.330 4.980 175.390 ;
        RECT 5.135 175.345 5.425 175.390 ;
        RECT 15.700 175.530 16.020 175.590 ;
        RECT 15.700 175.390 21.910 175.530 ;
        RECT 15.700 175.330 16.020 175.390 ;
        RECT 5.600 175.190 5.890 175.235 ;
        RECT 7.435 175.190 7.725 175.235 ;
        RECT 11.015 175.190 11.305 175.235 ;
        RECT 5.600 175.050 11.305 175.190 ;
        RECT 5.600 175.005 5.890 175.050 ;
        RECT 7.435 175.005 7.725 175.050 ;
        RECT 11.015 175.005 11.305 175.050 ;
        RECT 11.560 175.190 11.880 175.250 ;
        RECT 12.095 175.190 12.385 175.210 ;
        RECT 11.560 175.050 12.385 175.190 ;
        RECT 11.560 174.990 11.880 175.050 ;
        RECT 6.500 174.650 6.820 174.910 ;
        RECT 12.095 174.895 12.385 175.050 ;
        RECT 17.080 174.990 17.400 175.250 ;
        RECT 17.555 175.190 17.845 175.235 ;
        RECT 18.000 175.190 18.320 175.250 ;
        RECT 17.555 175.050 18.320 175.190 ;
        RECT 17.555 175.005 17.845 175.050 ;
        RECT 18.000 174.990 18.320 175.050 ;
        RECT 18.935 175.005 19.225 175.235 ;
        RECT 20.315 175.190 20.605 175.235 ;
        RECT 19.470 175.050 20.605 175.190 ;
        RECT 8.795 174.850 9.445 174.895 ;
        RECT 12.095 174.850 12.685 174.895 ;
        RECT 8.795 174.710 12.685 174.850 ;
        RECT 17.170 174.850 17.310 174.990 ;
        RECT 19.010 174.850 19.150 175.005 ;
        RECT 19.470 174.910 19.610 175.050 ;
        RECT 20.315 175.005 20.605 175.050 ;
        RECT 20.775 175.190 21.065 175.235 ;
        RECT 21.220 175.190 21.540 175.250 ;
        RECT 20.775 175.050 21.540 175.190 ;
        RECT 21.770 175.190 21.910 175.390 ;
        RECT 23.060 175.330 23.380 175.590 ;
        RECT 34.560 175.330 34.880 175.590 ;
        RECT 38.240 175.330 38.560 175.590 ;
        RECT 38.700 175.530 39.020 175.590 ;
        RECT 39.175 175.530 39.465 175.575 ;
        RECT 40.540 175.530 40.860 175.590 ;
        RECT 38.700 175.390 40.860 175.530 ;
        RECT 41.550 175.530 41.690 175.730 ;
        RECT 46.610 175.730 48.220 175.870 ;
        RECT 45.155 175.530 45.445 175.575 ;
        RECT 45.600 175.530 45.920 175.590 ;
        RECT 41.550 175.390 42.610 175.530 ;
        RECT 38.700 175.330 39.020 175.390 ;
        RECT 39.175 175.345 39.465 175.390 ;
        RECT 40.540 175.330 40.860 175.390 ;
        RECT 23.535 175.190 23.825 175.235 ;
        RECT 21.770 175.050 23.825 175.190 ;
        RECT 20.775 175.005 21.065 175.050 ;
        RECT 21.220 174.990 21.540 175.050 ;
        RECT 23.535 175.005 23.825 175.050 ;
        RECT 23.995 175.190 24.285 175.235 ;
        RECT 28.120 175.190 28.440 175.250 ;
        RECT 42.470 175.190 42.610 175.390 ;
        RECT 45.155 175.390 45.920 175.530 ;
        RECT 45.155 175.345 45.445 175.390 ;
        RECT 45.600 175.330 45.920 175.390 ;
        RECT 44.220 175.190 44.540 175.250 ;
        RECT 46.610 175.235 46.750 175.730 ;
        RECT 47.900 175.670 48.220 175.730 ;
        RECT 49.755 175.870 50.045 175.915 ;
        RECT 52.040 175.870 52.360 175.930 ;
        RECT 53.880 175.870 54.200 175.930 ;
        RECT 57.525 175.870 57.815 175.915 ;
        RECT 59.415 175.870 59.705 175.915 ;
        RECT 62.535 175.870 62.825 175.915 ;
        RECT 49.755 175.730 51.375 175.870 ;
        RECT 49.755 175.685 50.045 175.730 ;
        RECT 50.215 175.530 50.505 175.575 ;
        RECT 47.990 175.390 50.505 175.530 ;
        RECT 51.235 175.530 51.375 175.730 ;
        RECT 52.040 175.730 54.570 175.870 ;
        RECT 52.040 175.670 52.360 175.730 ;
        RECT 53.880 175.670 54.200 175.730 ;
        RECT 54.430 175.575 54.570 175.730 ;
        RECT 57.525 175.730 62.825 175.870 ;
        RECT 57.525 175.685 57.815 175.730 ;
        RECT 59.415 175.685 59.705 175.730 ;
        RECT 62.535 175.685 62.825 175.730 ;
        RECT 54.355 175.530 54.645 175.575 ;
        RECT 55.720 175.530 56.040 175.590 ;
        RECT 51.235 175.390 52.730 175.530 ;
        RECT 47.440 175.235 47.760 175.250 ;
        RECT 47.990 175.235 48.130 175.390 ;
        RECT 50.215 175.345 50.505 175.390 ;
        RECT 52.590 175.235 52.730 175.390 ;
        RECT 54.355 175.390 56.040 175.530 ;
        RECT 54.355 175.345 54.645 175.390 ;
        RECT 55.720 175.330 56.040 175.390 ;
        RECT 56.655 175.530 56.945 175.575 ;
        RECT 59.860 175.530 60.180 175.590 ;
        RECT 56.655 175.390 60.180 175.530 ;
        RECT 63.170 175.530 63.310 176.070 ;
        RECT 69.075 176.070 71.205 176.210 ;
        RECT 69.075 176.025 69.365 176.070 ;
        RECT 70.915 176.025 71.205 176.070 ;
        RECT 75.500 176.010 75.820 176.270 ;
        RECT 75.960 176.210 76.280 176.270 ;
        RECT 81.940 176.210 82.260 176.270 ;
        RECT 75.960 176.070 82.260 176.210 ;
        RECT 75.960 176.010 76.280 176.070 ;
        RECT 81.940 176.010 82.260 176.070 ;
        RECT 83.780 176.210 84.100 176.270 ;
        RECT 87.475 176.210 87.765 176.255 ;
        RECT 88.840 176.210 89.160 176.270 ;
        RECT 91.600 176.210 91.920 176.270 ;
        RECT 83.780 176.070 88.150 176.210 ;
        RECT 83.780 176.010 84.100 176.070 ;
        RECT 87.475 176.025 87.765 176.070 ;
        RECT 65.380 175.870 65.700 175.930 ;
        RECT 65.380 175.730 72.510 175.870 ;
        RECT 65.380 175.670 65.700 175.730 ;
        RECT 72.370 175.575 72.510 175.730 ;
        RECT 63.170 175.390 71.130 175.530 ;
        RECT 56.655 175.345 56.945 175.390 ;
        RECT 59.860 175.330 60.180 175.390 ;
        RECT 70.990 175.250 71.130 175.390 ;
        RECT 72.295 175.345 72.585 175.575 ;
        RECT 74.595 175.530 74.885 175.575 ;
        RECT 75.590 175.530 75.730 176.010 ;
        RECT 78.275 175.870 78.565 175.915 ;
        RECT 78.720 175.870 79.040 175.930 ;
        RECT 78.275 175.730 79.040 175.870 ;
        RECT 78.275 175.685 78.565 175.730 ;
        RECT 78.720 175.670 79.040 175.730 ;
        RECT 79.605 175.870 79.895 175.915 ;
        RECT 81.495 175.870 81.785 175.915 ;
        RECT 84.615 175.870 84.905 175.915 ;
        RECT 79.605 175.730 84.905 175.870 ;
        RECT 79.605 175.685 79.895 175.730 ;
        RECT 81.495 175.685 81.785 175.730 ;
        RECT 84.615 175.685 84.905 175.730 ;
        RECT 74.595 175.390 75.730 175.530 ;
        RECT 88.010 175.530 88.150 176.070 ;
        RECT 88.840 176.070 91.920 176.210 ;
        RECT 88.840 176.010 89.160 176.070 ;
        RECT 91.600 176.010 91.920 176.070 ;
        RECT 92.060 176.010 92.380 176.270 ;
        RECT 96.200 176.210 96.520 176.270 ;
        RECT 98.055 176.210 98.345 176.255 ;
        RECT 94.450 176.070 98.345 176.210 ;
        RECT 90.695 175.530 90.985 175.575 ;
        RECT 94.450 175.530 94.590 176.070 ;
        RECT 96.200 176.010 96.520 176.070 ;
        RECT 98.055 176.025 98.345 176.070 ;
        RECT 100.800 176.210 101.120 176.270 ;
        RECT 102.195 176.210 102.485 176.255 ;
        RECT 100.800 176.070 102.485 176.210 ;
        RECT 100.800 176.010 101.120 176.070 ;
        RECT 102.195 176.025 102.485 176.070 ;
        RECT 102.640 176.210 102.960 176.270 ;
        RECT 104.020 176.210 104.340 176.270 ;
        RECT 105.415 176.210 105.705 176.255 ;
        RECT 106.320 176.210 106.640 176.270 ;
        RECT 102.640 176.070 103.795 176.210 ;
        RECT 95.740 175.870 96.060 175.930 ;
        RECT 96.675 175.870 96.965 175.915 ;
        RECT 95.740 175.730 96.965 175.870 ;
        RECT 95.740 175.670 96.060 175.730 ;
        RECT 96.675 175.685 96.965 175.730 ;
        RECT 97.580 175.870 97.900 175.930 ;
        RECT 100.340 175.870 100.660 175.930 ;
        RECT 97.580 175.730 100.660 175.870 ;
        RECT 97.580 175.670 97.900 175.730 ;
        RECT 100.340 175.670 100.660 175.730 ;
        RECT 88.010 175.390 90.985 175.530 ;
        RECT 74.595 175.345 74.885 175.390 ;
        RECT 90.695 175.345 90.985 175.390 ;
        RECT 91.230 175.390 94.590 175.530 ;
        RECT 23.995 175.050 28.440 175.190 ;
        RECT 23.995 175.005 24.285 175.050 ;
        RECT 17.170 174.710 19.150 174.850 ;
        RECT 8.795 174.665 9.445 174.710 ;
        RECT 12.395 174.665 12.685 174.710 ;
        RECT 19.380 174.650 19.700 174.910 ;
        RECT 19.840 174.650 20.160 174.910 ;
        RECT 22.600 174.850 22.920 174.910 ;
        RECT 24.070 174.850 24.210 175.005 ;
        RECT 28.120 174.990 28.440 175.050 ;
        RECT 28.670 175.050 42.150 175.190 ;
        RECT 42.470 175.050 44.540 175.190 ;
        RECT 22.600 174.710 24.210 174.850 ;
        RECT 24.440 174.850 24.760 174.910 ;
        RECT 27.200 174.850 27.520 174.910 ;
        RECT 28.670 174.850 28.810 175.050 ;
        RECT 35.035 174.850 35.325 174.895 ;
        RECT 35.480 174.850 35.800 174.910 ;
        RECT 41.460 174.850 41.780 174.910 ;
        RECT 24.440 174.710 26.970 174.850 ;
        RECT 22.600 174.650 22.920 174.710 ;
        RECT 24.440 174.650 24.760 174.710 ;
        RECT 20.760 174.510 21.080 174.570 ;
        RECT 21.695 174.510 21.985 174.555 ;
        RECT 20.760 174.370 21.985 174.510 ;
        RECT 20.760 174.310 21.080 174.370 ;
        RECT 21.695 174.325 21.985 174.370 ;
        RECT 25.820 174.310 26.140 174.570 ;
        RECT 26.830 174.510 26.970 174.710 ;
        RECT 27.200 174.710 28.810 174.850 ;
        RECT 29.590 174.710 35.800 174.850 ;
        RECT 27.200 174.650 27.520 174.710 ;
        RECT 29.590 174.510 29.730 174.710 ;
        RECT 35.035 174.665 35.325 174.710 ;
        RECT 35.480 174.650 35.800 174.710 ;
        RECT 39.250 174.710 41.780 174.850 ;
        RECT 42.010 174.850 42.150 175.050 ;
        RECT 44.220 174.990 44.540 175.050 ;
        RECT 46.535 175.005 46.825 175.235 ;
        RECT 47.275 175.005 47.760 175.235 ;
        RECT 47.915 175.005 48.205 175.235 ;
        RECT 49.065 175.190 49.355 175.235 ;
        RECT 49.065 175.050 50.430 175.190 ;
        RECT 49.065 175.005 49.355 175.050 ;
        RECT 47.440 174.990 47.760 175.005 ;
        RECT 50.290 174.910 50.430 175.050 ;
        RECT 52.515 175.005 52.805 175.235 ;
        RECT 52.960 175.190 53.280 175.250 ;
        RECT 53.435 175.190 53.725 175.235 ;
        RECT 52.960 175.050 53.725 175.190 ;
        RECT 52.960 174.990 53.280 175.050 ;
        RECT 53.435 175.005 53.725 175.050 ;
        RECT 48.375 174.850 48.665 174.895 ;
        RECT 42.010 174.710 48.665 174.850 ;
        RECT 26.830 174.370 29.730 174.510 ;
        RECT 32.720 174.510 33.040 174.570 ;
        RECT 33.655 174.510 33.945 174.555 ;
        RECT 32.720 174.370 33.945 174.510 ;
        RECT 32.720 174.310 33.040 174.370 ;
        RECT 33.655 174.325 33.945 174.370 ;
        RECT 37.795 174.510 38.085 174.555 ;
        RECT 39.250 174.510 39.390 174.710 ;
        RECT 41.460 174.650 41.780 174.710 ;
        RECT 48.375 174.665 48.665 174.710 ;
        RECT 50.200 174.650 50.520 174.910 ;
        RECT 51.135 174.850 51.425 174.895 ;
        RECT 51.580 174.850 51.900 174.910 ;
        RECT 51.135 174.710 51.900 174.850 ;
        RECT 51.135 174.665 51.425 174.710 ;
        RECT 51.580 174.650 51.900 174.710 ;
        RECT 52.055 174.665 52.345 174.895 ;
        RECT 53.510 174.850 53.650 175.005 ;
        RECT 53.880 174.990 54.200 175.250 ;
        RECT 55.275 175.190 55.565 175.235 ;
        RECT 57.120 175.190 57.410 175.235 ;
        RECT 58.955 175.190 59.245 175.235 ;
        RECT 62.535 175.190 62.825 175.235 ;
        RECT 55.275 175.050 55.950 175.190 ;
        RECT 55.275 175.005 55.565 175.050 ;
        RECT 53.510 174.710 55.490 174.850 ;
        RECT 37.795 174.370 39.390 174.510 ;
        RECT 39.620 174.510 39.940 174.570 ;
        RECT 41.935 174.510 42.225 174.555 ;
        RECT 39.620 174.370 42.225 174.510 ;
        RECT 37.795 174.325 38.085 174.370 ;
        RECT 39.620 174.310 39.940 174.370 ;
        RECT 41.935 174.325 42.225 174.370 ;
        RECT 43.760 174.310 44.080 174.570 ;
        RECT 45.140 174.510 45.460 174.570 ;
        RECT 46.520 174.510 46.840 174.570 ;
        RECT 45.140 174.370 46.840 174.510 ;
        RECT 45.140 174.310 45.460 174.370 ;
        RECT 46.520 174.310 46.840 174.370 ;
        RECT 49.740 174.510 50.060 174.570 ;
        RECT 52.130 174.510 52.270 174.665 ;
        RECT 55.350 174.570 55.490 174.710 ;
        RECT 49.740 174.370 52.270 174.510 ;
        RECT 49.740 174.310 50.060 174.370 ;
        RECT 55.260 174.310 55.580 174.570 ;
        RECT 55.810 174.510 55.950 175.050 ;
        RECT 57.120 175.050 62.825 175.190 ;
        RECT 57.120 175.005 57.410 175.050 ;
        RECT 58.955 175.005 59.245 175.050 ;
        RECT 62.535 175.005 62.825 175.050 ;
        RECT 56.195 174.850 56.485 174.895 ;
        RECT 58.035 174.850 58.325 174.895 ;
        RECT 56.195 174.710 58.325 174.850 ;
        RECT 56.195 174.665 56.485 174.710 ;
        RECT 58.035 174.665 58.325 174.710 ;
        RECT 58.480 174.650 58.800 174.910 ;
        RECT 60.315 174.850 60.965 174.895 ;
        RECT 61.700 174.850 62.020 174.910 ;
        RECT 63.615 174.895 63.905 175.210 ;
        RECT 69.980 174.990 70.300 175.250 ;
        RECT 70.900 174.990 71.220 175.250 ;
        RECT 71.375 175.005 71.665 175.235 ;
        RECT 75.960 175.190 76.280 175.250 ;
        RECT 78.735 175.190 79.025 175.235 ;
        RECT 75.960 175.050 79.025 175.190 ;
        RECT 63.615 174.850 64.205 174.895 ;
        RECT 60.315 174.710 64.205 174.850 ;
        RECT 60.315 174.665 60.965 174.710 ;
        RECT 61.700 174.650 62.020 174.710 ;
        RECT 63.915 174.665 64.205 174.710 ;
        RECT 69.060 174.850 69.380 174.910 ;
        RECT 71.450 174.850 71.590 175.005 ;
        RECT 75.960 174.990 76.280 175.050 ;
        RECT 78.735 175.005 79.025 175.050 ;
        RECT 79.200 175.190 79.490 175.235 ;
        RECT 81.035 175.190 81.325 175.235 ;
        RECT 84.615 175.190 84.905 175.235 ;
        RECT 79.200 175.050 84.905 175.190 ;
        RECT 79.200 175.005 79.490 175.050 ;
        RECT 81.035 175.005 81.325 175.050 ;
        RECT 84.615 175.005 84.905 175.050 ;
        RECT 72.280 174.850 72.600 174.910 ;
        RECT 69.060 174.710 72.600 174.850 ;
        RECT 69.060 174.650 69.380 174.710 ;
        RECT 72.280 174.650 72.600 174.710 ;
        RECT 74.580 174.850 74.900 174.910 ;
        RECT 75.515 174.850 75.805 174.895 ;
        RECT 74.580 174.710 75.805 174.850 ;
        RECT 74.580 174.650 74.900 174.710 ;
        RECT 75.515 174.665 75.805 174.710 ;
        RECT 77.340 174.650 77.660 174.910 ;
        RECT 85.695 174.895 85.985 175.210 ;
        RECT 90.220 175.190 90.540 175.250 ;
        RECT 91.230 175.190 91.370 175.390 ;
        RECT 94.450 175.235 94.590 175.390 ;
        RECT 90.220 175.050 91.370 175.190 ;
        RECT 90.220 174.990 90.540 175.050 ;
        RECT 91.615 175.005 91.905 175.235 ;
        RECT 92.535 175.005 92.825 175.235 ;
        RECT 93.455 175.005 93.745 175.235 ;
        RECT 94.375 175.005 94.665 175.235 ;
        RECT 94.835 175.005 95.125 175.235 ;
        RECT 95.465 175.190 95.755 175.235 ;
        RECT 100.890 175.190 101.030 176.010 ;
        RECT 102.270 175.870 102.410 176.025 ;
        RECT 102.640 176.010 102.960 176.070 ;
        RECT 102.270 175.730 103.330 175.870 ;
        RECT 101.720 175.330 102.040 175.590 ;
        RECT 103.190 175.250 103.330 175.730 ;
        RECT 103.655 175.530 103.795 176.070 ;
        RECT 104.020 176.070 106.640 176.210 ;
        RECT 104.020 176.010 104.340 176.070 ;
        RECT 105.415 176.025 105.705 176.070 ;
        RECT 106.320 176.010 106.640 176.070 ;
        RECT 107.255 176.210 107.545 176.255 ;
        RECT 110.460 176.210 110.780 176.270 ;
        RECT 107.255 176.070 110.780 176.210 ;
        RECT 107.255 176.025 107.545 176.070 ;
        RECT 110.460 176.010 110.780 176.070 ;
        RECT 113.680 176.210 114.000 176.270 ;
        RECT 116.455 176.210 116.745 176.255 ;
        RECT 113.680 176.070 116.745 176.210 ;
        RECT 113.680 176.010 114.000 176.070 ;
        RECT 116.455 176.025 116.745 176.070 ;
        RECT 117.375 176.210 117.665 176.255 ;
        RECT 118.280 176.210 118.600 176.270 ;
        RECT 117.375 176.070 118.600 176.210 ;
        RECT 117.375 176.025 117.665 176.070 ;
        RECT 118.280 176.010 118.600 176.070 ;
        RECT 122.435 176.210 122.725 176.255 ;
        RECT 122.880 176.210 123.200 176.270 ;
        RECT 122.435 176.070 123.200 176.210 ;
        RECT 122.435 176.025 122.725 176.070 ;
        RECT 122.880 176.010 123.200 176.070 ;
        RECT 124.260 176.210 124.580 176.270 ;
        RECT 124.735 176.210 125.025 176.255 ;
        RECT 125.180 176.210 125.500 176.270 ;
        RECT 124.260 176.070 125.500 176.210 ;
        RECT 124.260 176.010 124.580 176.070 ;
        RECT 124.735 176.025 125.025 176.070 ;
        RECT 125.180 176.010 125.500 176.070 ;
        RECT 125.655 176.210 125.945 176.255 ;
        RECT 127.940 176.210 128.260 176.270 ;
        RECT 125.655 176.070 128.260 176.210 ;
        RECT 125.655 176.025 125.945 176.070 ;
        RECT 127.940 176.010 128.260 176.070 ;
        RECT 128.860 176.010 129.180 176.270 ;
        RECT 129.320 176.210 129.640 176.270 ;
        RECT 136.680 176.210 137.000 176.270 ;
        RECT 137.155 176.210 137.445 176.255 ;
        RECT 129.320 176.070 136.400 176.210 ;
        RECT 129.320 176.010 129.640 176.070 ;
        RECT 104.480 175.870 104.800 175.930 ;
        RECT 104.955 175.870 105.245 175.915 ;
        RECT 104.480 175.730 105.245 175.870 ;
        RECT 104.480 175.670 104.800 175.730 ;
        RECT 104.955 175.685 105.245 175.730 ;
        RECT 108.635 175.870 108.925 175.915 ;
        RECT 108.635 175.730 135.990 175.870 ;
        RECT 108.635 175.685 108.925 175.730 ;
        RECT 110.000 175.530 110.320 175.590 ;
        RECT 114.600 175.530 114.920 175.590 ;
        RECT 120.580 175.530 120.900 175.590 ;
        RECT 103.655 175.390 108.850 175.530 ;
        RECT 95.465 175.050 101.030 175.190 ;
        RECT 102.195 175.190 102.485 175.235 ;
        RECT 102.655 175.190 102.945 175.235 ;
        RECT 102.195 175.050 102.945 175.190 ;
        RECT 95.465 175.005 95.755 175.050 ;
        RECT 102.195 175.005 102.485 175.050 ;
        RECT 102.655 175.005 102.945 175.050 ;
        RECT 103.100 175.190 103.420 175.250 ;
        RECT 103.575 175.190 103.865 175.235 ;
        RECT 103.100 175.050 103.865 175.190 ;
        RECT 80.115 174.665 80.405 174.895 ;
        RECT 82.395 174.850 83.045 174.895 ;
        RECT 85.695 174.850 86.285 174.895 ;
        RECT 86.540 174.850 86.860 174.910 ;
        RECT 82.395 174.710 86.860 174.850 ;
        RECT 82.395 174.665 83.045 174.710 ;
        RECT 85.995 174.665 86.285 174.710 ;
        RECT 58.570 174.510 58.710 174.650 ;
        RECT 55.810 174.370 58.710 174.510 ;
        RECT 71.360 174.510 71.680 174.570 ;
        RECT 75.960 174.510 76.280 174.570 ;
        RECT 76.435 174.510 76.725 174.555 ;
        RECT 71.360 174.370 76.725 174.510 ;
        RECT 71.360 174.310 71.680 174.370 ;
        RECT 75.960 174.310 76.280 174.370 ;
        RECT 76.435 174.325 76.725 174.370 ;
        RECT 76.895 174.510 77.185 174.555 ;
        RECT 79.180 174.510 79.500 174.570 ;
        RECT 76.895 174.370 79.500 174.510 ;
        RECT 80.190 174.510 80.330 174.665 ;
        RECT 86.540 174.650 86.860 174.710 ;
        RECT 89.300 174.850 89.620 174.910 ;
        RECT 91.690 174.850 91.830 175.005 ;
        RECT 89.300 174.710 91.830 174.850 ;
        RECT 92.060 174.850 92.380 174.910 ;
        RECT 92.610 174.850 92.750 175.005 ;
        RECT 92.060 174.710 92.750 174.850 ;
        RECT 89.300 174.650 89.620 174.710 ;
        RECT 92.060 174.650 92.380 174.710 ;
        RECT 83.780 174.510 84.100 174.570 ;
        RECT 80.190 174.370 84.100 174.510 ;
        RECT 76.895 174.325 77.185 174.370 ;
        RECT 79.180 174.310 79.500 174.370 ;
        RECT 83.780 174.310 84.100 174.370 ;
        RECT 87.920 174.310 88.240 174.570 ;
        RECT 89.760 174.510 90.080 174.570 ;
        RECT 93.530 174.510 93.670 175.005 ;
        RECT 94.910 174.850 95.050 175.005 ;
        RECT 94.910 174.710 95.510 174.850 ;
        RECT 95.370 174.570 95.510 174.710 ;
        RECT 97.120 174.650 97.440 174.910 ;
        RECT 102.270 174.850 102.410 175.005 ;
        RECT 103.100 174.990 103.420 175.050 ;
        RECT 103.575 175.005 103.865 175.050 ;
        RECT 104.020 174.990 104.340 175.250 ;
        RECT 105.490 175.235 105.630 175.390 ;
        RECT 105.415 175.005 105.705 175.235 ;
        RECT 105.875 175.005 106.165 175.235 ;
        RECT 106.320 175.190 106.640 175.250 ;
        RECT 108.710 175.235 108.850 175.390 ;
        RECT 110.000 175.390 114.920 175.530 ;
        RECT 110.000 175.330 110.320 175.390 ;
        RECT 114.600 175.330 114.920 175.390 ;
        RECT 115.150 175.390 120.900 175.530 ;
        RECT 107.715 175.190 108.005 175.235 ;
        RECT 106.320 175.050 108.005 175.190 ;
        RECT 97.670 174.710 102.410 174.850 ;
        RECT 104.480 174.850 104.800 174.910 ;
        RECT 105.950 174.850 106.090 175.005 ;
        RECT 106.320 174.990 106.640 175.050 ;
        RECT 107.715 175.005 108.005 175.050 ;
        RECT 108.635 175.005 108.925 175.235 ;
        RECT 111.380 174.990 111.700 175.250 ;
        RECT 112.300 175.190 112.620 175.250 ;
        RECT 115.150 175.190 115.290 175.390 ;
        RECT 120.580 175.330 120.900 175.390 ;
        RECT 121.055 175.530 121.345 175.575 ;
        RECT 125.640 175.530 125.960 175.590 ;
        RECT 121.055 175.390 128.170 175.530 ;
        RECT 121.055 175.345 121.345 175.390 ;
        RECT 125.640 175.330 125.960 175.390 ;
        RECT 123.355 175.190 123.645 175.235 ;
        RECT 124.260 175.190 124.580 175.250 ;
        RECT 126.575 175.190 126.865 175.235 ;
        RECT 127.020 175.190 127.340 175.250 ;
        RECT 128.030 175.235 128.170 175.390 ;
        RECT 112.300 175.050 115.290 175.190 ;
        RECT 115.610 175.050 122.650 175.190 ;
        RECT 112.300 174.990 112.620 175.050 ;
        RECT 115.610 174.895 115.750 175.050 ;
        RECT 113.235 174.850 113.525 174.895 ;
        RECT 115.535 174.850 115.825 174.895 ;
        RECT 104.480 174.710 115.825 174.850 ;
        RECT 89.760 174.370 93.670 174.510 ;
        RECT 95.280 174.510 95.600 174.570 ;
        RECT 97.670 174.510 97.810 174.710 ;
        RECT 104.480 174.650 104.800 174.710 ;
        RECT 113.235 174.665 113.525 174.710 ;
        RECT 115.535 174.665 115.825 174.710 ;
        RECT 115.980 174.850 116.300 174.910 ;
        RECT 119.675 174.850 119.965 174.895 ;
        RECT 115.980 174.710 119.965 174.850 ;
        RECT 115.980 174.650 116.300 174.710 ;
        RECT 119.675 174.665 119.965 174.710 ;
        RECT 95.280 174.370 97.810 174.510 ;
        RECT 89.760 174.310 90.080 174.370 ;
        RECT 95.280 174.310 95.600 174.370 ;
        RECT 98.040 174.310 98.360 174.570 ;
        RECT 98.975 174.510 99.265 174.555 ;
        RECT 107.700 174.510 108.020 174.570 ;
        RECT 98.975 174.370 108.020 174.510 ;
        RECT 98.975 174.325 99.265 174.370 ;
        RECT 107.700 174.310 108.020 174.370 ;
        RECT 108.160 174.510 108.480 174.570 ;
        RECT 110.475 174.510 110.765 174.555 ;
        RECT 108.160 174.370 110.765 174.510 ;
        RECT 108.160 174.310 108.480 174.370 ;
        RECT 110.475 174.325 110.765 174.370 ;
        RECT 116.585 174.510 116.875 174.555 ;
        RECT 117.820 174.510 118.140 174.570 ;
        RECT 121.960 174.510 122.280 174.570 ;
        RECT 116.585 174.370 122.280 174.510 ;
        RECT 122.510 174.510 122.650 175.050 ;
        RECT 123.355 175.050 124.580 175.190 ;
        RECT 123.355 175.005 123.645 175.050 ;
        RECT 124.260 174.990 124.580 175.050 ;
        RECT 124.810 175.050 127.340 175.190 ;
        RECT 123.800 174.650 124.120 174.910 ;
        RECT 123.340 174.510 123.660 174.570 ;
        RECT 124.810 174.555 124.950 175.050 ;
        RECT 126.575 175.005 126.865 175.050 ;
        RECT 127.020 174.990 127.340 175.050 ;
        RECT 127.955 175.005 128.245 175.235 ;
        RECT 133.475 175.190 133.765 175.235 ;
        RECT 135.300 175.190 135.620 175.250 ;
        RECT 133.475 175.050 135.620 175.190 ;
        RECT 135.850 175.190 135.990 175.730 ;
        RECT 136.260 175.530 136.400 176.070 ;
        RECT 136.680 176.070 137.445 176.210 ;
        RECT 136.680 176.010 137.000 176.070 ;
        RECT 137.155 176.025 137.445 176.070 ;
        RECT 138.535 176.210 138.825 176.255 ;
        RECT 139.900 176.210 140.220 176.270 ;
        RECT 138.535 176.070 140.220 176.210 ;
        RECT 138.535 176.025 138.825 176.070 ;
        RECT 139.900 176.010 140.220 176.070 ;
        RECT 149.100 176.210 149.420 176.270 ;
        RECT 149.575 176.210 149.865 176.255 ;
        RECT 149.100 176.070 149.865 176.210 ;
        RECT 149.100 176.010 149.420 176.070 ;
        RECT 149.575 176.025 149.865 176.070 ;
        RECT 151.400 176.010 151.720 176.270 ;
        RECT 153.240 176.010 153.560 176.270 ;
        RECT 140.820 175.870 141.140 175.930 ;
        RECT 137.690 175.730 141.140 175.870 ;
        RECT 137.690 175.590 137.830 175.730 ;
        RECT 140.820 175.670 141.140 175.730 ;
        RECT 136.695 175.530 136.985 175.575 ;
        RECT 136.260 175.390 136.985 175.530 ;
        RECT 136.695 175.345 136.985 175.390 ;
        RECT 137.600 175.330 137.920 175.590 ;
        RECT 153.330 175.530 153.470 176.010 ;
        RECT 138.150 175.390 153.470 175.530 ;
        RECT 136.235 175.190 136.525 175.235 ;
        RECT 135.850 175.050 136.525 175.190 ;
        RECT 133.475 175.005 133.765 175.050 ;
        RECT 135.300 174.990 135.620 175.050 ;
        RECT 136.235 175.005 136.525 175.050 ;
        RECT 137.140 175.190 137.460 175.250 ;
        RECT 138.150 175.190 138.290 175.390 ;
        RECT 137.140 175.050 138.290 175.190 ;
        RECT 139.915 175.190 140.205 175.235 ;
        RECT 141.280 175.190 141.600 175.250 ;
        RECT 149.650 175.235 149.790 175.390 ;
        RECT 139.915 175.050 141.600 175.190 ;
        RECT 125.180 174.850 125.500 174.910 ;
        RECT 125.180 174.710 127.250 174.850 ;
        RECT 125.180 174.650 125.500 174.710 ;
        RECT 127.110 174.555 127.250 174.710 ;
        RECT 131.620 174.650 131.940 174.910 ;
        RECT 134.380 174.650 134.700 174.910 ;
        RECT 136.310 174.850 136.450 175.005 ;
        RECT 137.140 174.990 137.460 175.050 ;
        RECT 139.915 175.005 140.205 175.050 ;
        RECT 141.280 174.990 141.600 175.050 ;
        RECT 149.575 175.005 149.865 175.235 ;
        RECT 150.035 175.005 150.325 175.235 ;
        RECT 138.535 174.850 138.825 174.895 ;
        RECT 150.110 174.850 150.250 175.005 ;
        RECT 151.860 174.990 152.180 175.250 ;
        RECT 136.310 174.710 138.825 174.850 ;
        RECT 138.535 174.665 138.825 174.710 ;
        RECT 139.070 174.710 150.250 174.850 ;
        RECT 122.510 174.370 123.660 174.510 ;
        RECT 116.585 174.325 116.875 174.370 ;
        RECT 117.820 174.310 118.140 174.370 ;
        RECT 121.960 174.310 122.280 174.370 ;
        RECT 123.340 174.310 123.660 174.370 ;
        RECT 124.735 174.325 125.025 174.555 ;
        RECT 127.035 174.325 127.325 174.555 ;
        RECT 134.840 174.510 135.160 174.570 ;
        RECT 139.070 174.510 139.210 174.710 ;
        RECT 134.840 174.370 139.210 174.510 ;
        RECT 139.455 174.510 139.745 174.555 ;
        RECT 151.950 174.510 152.090 174.990 ;
        RECT 139.455 174.370 152.090 174.510 ;
        RECT 134.840 174.310 135.160 174.370 ;
        RECT 139.455 174.325 139.745 174.370 ;
        RECT 2.750 173.690 159.030 174.170 ;
        RECT 6.500 173.490 6.820 173.550 ;
        RECT 7.435 173.490 7.725 173.535 ;
        RECT 13.860 173.490 14.180 173.550 ;
        RECT 6.500 173.350 7.725 173.490 ;
        RECT 6.500 173.290 6.820 173.350 ;
        RECT 7.435 173.305 7.725 173.350 ;
        RECT 13.720 173.290 14.180 173.490 ;
        RECT 19.380 173.490 19.700 173.550 ;
        RECT 23.995 173.490 24.285 173.535 ;
        RECT 26.740 173.490 27.060 173.550 ;
        RECT 19.380 173.350 27.060 173.490 ;
        RECT 19.380 173.290 19.700 173.350 ;
        RECT 23.995 173.305 24.285 173.350 ;
        RECT 26.740 173.290 27.060 173.350 ;
        RECT 31.340 173.490 31.660 173.550 ;
        RECT 33.195 173.490 33.485 173.535 ;
        RECT 31.340 173.350 33.485 173.490 ;
        RECT 31.340 173.290 31.660 173.350 ;
        RECT 33.195 173.305 33.485 173.350 ;
        RECT 43.760 173.490 44.080 173.550 ;
        RECT 46.075 173.490 46.365 173.535 ;
        RECT 43.760 173.350 46.365 173.490 ;
        RECT 43.760 173.290 44.080 173.350 ;
        RECT 46.075 173.305 46.365 173.350 ;
        RECT 46.980 173.490 47.300 173.550 ;
        RECT 48.360 173.490 48.680 173.550 ;
        RECT 51.120 173.490 51.440 173.550 ;
        RECT 46.980 173.350 48.680 173.490 ;
        RECT 46.980 173.290 47.300 173.350 ;
        RECT 48.360 173.290 48.680 173.350 ;
        RECT 49.375 173.350 50.890 173.490 ;
        RECT 12.035 173.150 12.325 173.195 ;
        RECT 13.720 173.150 13.860 173.290 ;
        RECT 12.035 173.010 13.860 173.150 ;
        RECT 12.035 172.965 12.325 173.010 ;
        RECT 19.840 172.950 20.160 173.210 ;
        RECT 20.300 173.150 20.620 173.210 ;
        RECT 22.600 173.150 22.920 173.210 ;
        RECT 20.300 173.010 22.920 173.150 ;
        RECT 20.300 172.950 20.620 173.010 ;
        RECT 22.600 172.950 22.920 173.010 ;
        RECT 23.060 173.150 23.380 173.210 ;
        RECT 31.800 173.150 32.120 173.210 ;
        RECT 23.060 173.010 32.120 173.150 ;
        RECT 23.060 172.950 23.380 173.010 ;
        RECT 31.800 172.950 32.120 173.010 ;
        RECT 40.995 173.150 41.645 173.195 ;
        RECT 42.380 173.150 42.700 173.210 ;
        RECT 44.595 173.150 44.885 173.195 ;
        RECT 40.995 173.010 44.885 173.150 ;
        RECT 40.995 172.965 41.645 173.010 ;
        RECT 42.380 172.950 42.700 173.010 ;
        RECT 44.295 172.965 44.885 173.010 ;
        RECT 45.600 173.150 45.920 173.210 ;
        RECT 47.900 173.150 48.220 173.210 ;
        RECT 49.375 173.150 49.515 173.350 ;
        RECT 45.600 173.010 47.670 173.150 ;
        RECT 8.355 172.810 8.645 172.855 ;
        RECT 8.355 172.670 10.410 172.810 ;
        RECT 8.355 172.625 8.645 172.670 ;
        RECT 10.270 172.175 10.410 172.670 ;
        RECT 18.920 172.610 19.240 172.870 ;
        RECT 20.775 172.810 21.065 172.855 ;
        RECT 21.220 172.810 21.540 172.870 ;
        RECT 25.360 172.810 25.680 172.870 ;
        RECT 20.775 172.670 25.680 172.810 ;
        RECT 20.775 172.625 21.065 172.670 ;
        RECT 21.220 172.610 21.540 172.670 ;
        RECT 25.360 172.610 25.680 172.670 ;
        RECT 30.435 172.810 30.725 172.855 ;
        RECT 32.735 172.810 33.025 172.855 ;
        RECT 36.860 172.810 37.180 172.870 ;
        RECT 30.435 172.670 31.110 172.810 ;
        RECT 30.435 172.625 30.725 172.670 ;
        RECT 12.480 172.270 12.800 172.530 ;
        RECT 13.400 172.270 13.720 172.530 ;
        RECT 23.060 172.270 23.380 172.530 ;
        RECT 23.535 172.470 23.825 172.515 ;
        RECT 23.980 172.470 24.300 172.530 ;
        RECT 23.535 172.330 24.300 172.470 ;
        RECT 23.535 172.285 23.825 172.330 ;
        RECT 23.980 172.270 24.300 172.330 ;
        RECT 10.195 171.945 10.485 172.175 ;
        RECT 13.490 172.130 13.630 172.270 ;
        RECT 30.970 172.175 31.110 172.670 ;
        RECT 32.735 172.670 37.180 172.810 ;
        RECT 32.735 172.625 33.025 172.670 ;
        RECT 36.860 172.610 37.180 172.670 ;
        RECT 37.800 172.810 38.090 172.855 ;
        RECT 39.635 172.810 39.925 172.855 ;
        RECT 43.215 172.810 43.505 172.855 ;
        RECT 37.800 172.670 43.505 172.810 ;
        RECT 37.800 172.625 38.090 172.670 ;
        RECT 39.635 172.625 39.925 172.670 ;
        RECT 43.215 172.625 43.505 172.670 ;
        RECT 44.295 172.650 44.585 172.965 ;
        RECT 45.600 172.950 45.920 173.010 ;
        RECT 34.115 172.470 34.405 172.515 ;
        RECT 34.115 172.330 34.790 172.470 ;
        RECT 34.115 172.285 34.405 172.330 ;
        RECT 13.490 171.990 30.650 172.130 ;
        RECT 10.640 171.790 10.960 171.850 ;
        RECT 16.620 171.790 16.940 171.850 ;
        RECT 10.640 171.650 16.940 171.790 ;
        RECT 10.640 171.590 10.960 171.650 ;
        RECT 16.620 171.590 16.940 171.650 ;
        RECT 21.695 171.790 21.985 171.835 ;
        RECT 23.060 171.790 23.380 171.850 ;
        RECT 21.695 171.650 23.380 171.790 ;
        RECT 21.695 171.605 21.985 171.650 ;
        RECT 23.060 171.590 23.380 171.650 ;
        RECT 25.835 171.790 26.125 171.835 ;
        RECT 26.740 171.790 27.060 171.850 ;
        RECT 25.835 171.650 27.060 171.790 ;
        RECT 25.835 171.605 26.125 171.650 ;
        RECT 26.740 171.590 27.060 171.650 ;
        RECT 29.515 171.790 29.805 171.835 ;
        RECT 29.960 171.790 30.280 171.850 ;
        RECT 29.515 171.650 30.280 171.790 ;
        RECT 30.510 171.790 30.650 171.990 ;
        RECT 30.895 171.945 31.185 172.175 ;
        RECT 34.650 171.790 34.790 172.330 ;
        RECT 37.320 172.270 37.640 172.530 ;
        RECT 38.700 172.270 39.020 172.530 ;
        RECT 38.205 172.130 38.495 172.175 ;
        RECT 40.095 172.130 40.385 172.175 ;
        RECT 43.215 172.130 43.505 172.175 ;
        RECT 38.205 171.990 43.505 172.130 ;
        RECT 38.205 171.945 38.495 171.990 ;
        RECT 40.095 171.945 40.385 171.990 ;
        RECT 43.215 171.945 43.505 171.990 ;
        RECT 45.690 171.790 45.830 172.950 ;
        RECT 46.520 172.610 46.840 172.870 ;
        RECT 46.980 172.610 47.300 172.870 ;
        RECT 47.530 172.810 47.670 173.010 ;
        RECT 47.900 173.010 49.515 173.150 ;
        RECT 47.900 172.950 48.220 173.010 ;
        RECT 49.740 172.950 50.060 173.210 ;
        RECT 48.820 172.810 49.140 172.870 ;
        RECT 47.530 172.670 49.140 172.810 ;
        RECT 48.820 172.610 49.140 172.670 ;
        RECT 49.295 172.625 49.585 172.855 ;
        RECT 49.830 172.810 49.970 172.950 ;
        RECT 50.750 172.855 50.890 173.350 ;
        RECT 51.120 173.350 53.190 173.490 ;
        RECT 51.120 173.290 51.440 173.350 ;
        RECT 52.515 172.965 52.805 173.195 ;
        RECT 53.050 173.150 53.190 173.350 ;
        RECT 59.400 173.290 59.720 173.550 ;
        RECT 71.375 173.490 71.665 173.535 ;
        RECT 73.200 173.490 73.520 173.550 ;
        RECT 71.375 173.350 73.520 173.490 ;
        RECT 71.375 173.305 71.665 173.350 ;
        RECT 73.200 173.290 73.520 173.350 ;
        RECT 77.340 173.490 77.660 173.550 ;
        RECT 81.020 173.490 81.340 173.550 ;
        RECT 81.955 173.490 82.245 173.535 ;
        RECT 77.340 173.350 80.790 173.490 ;
        RECT 77.340 173.290 77.660 173.350 ;
        RECT 67.220 173.150 67.540 173.210 ;
        RECT 53.050 173.010 55.950 173.150 ;
        RECT 50.215 172.810 50.505 172.855 ;
        RECT 49.830 172.670 50.505 172.810 ;
        RECT 50.215 172.625 50.505 172.670 ;
        RECT 50.675 172.625 50.965 172.855 ;
        RECT 51.140 172.625 51.430 172.855 ;
        RECT 46.610 172.470 46.750 172.610 ;
        RECT 49.370 172.470 49.510 172.625 ;
        RECT 46.610 172.330 49.510 172.470 ;
        RECT 49.755 172.470 50.045 172.515 ;
        RECT 51.215 172.470 51.355 172.625 ;
        RECT 52.040 172.610 52.360 172.870 ;
        RECT 52.590 172.530 52.730 172.965 ;
        RECT 55.810 172.855 55.950 173.010 ;
        RECT 57.190 173.010 67.540 173.150 ;
        RECT 57.190 172.855 57.330 173.010 ;
        RECT 67.220 172.950 67.540 173.010 ;
        RECT 75.040 173.150 75.360 173.210 ;
        RECT 78.720 173.195 79.040 173.210 ;
        RECT 80.650 173.195 80.790 173.350 ;
        RECT 81.020 173.350 82.245 173.490 ;
        RECT 81.020 173.290 81.340 173.350 ;
        RECT 81.955 173.305 82.245 173.350 ;
        RECT 77.815 173.150 78.105 173.195 ;
        RECT 75.040 173.010 78.105 173.150 ;
        RECT 75.040 172.950 75.360 173.010 ;
        RECT 77.815 172.965 78.105 173.010 ;
        RECT 78.720 173.150 79.185 173.195 ;
        RECT 78.720 173.010 80.330 173.150 ;
        RECT 78.720 172.965 79.185 173.010 ;
        RECT 78.720 172.950 79.040 172.965 ;
        RECT 53.000 172.625 53.290 172.855 ;
        RECT 55.735 172.625 56.025 172.855 ;
        RECT 56.655 172.625 56.945 172.855 ;
        RECT 57.115 172.625 57.405 172.855 ;
        RECT 49.755 172.330 51.355 172.470 ;
        RECT 49.755 172.285 50.045 172.330 ;
        RECT 52.500 172.270 52.820 172.530 ;
        RECT 50.200 172.130 50.520 172.190 ;
        RECT 48.910 171.990 50.520 172.130 ;
        RECT 30.510 171.650 45.830 171.790 ;
        RECT 48.375 171.790 48.665 171.835 ;
        RECT 48.910 171.790 49.050 171.990 ;
        RECT 50.200 171.930 50.520 171.990 ;
        RECT 50.660 172.130 50.980 172.190 ;
        RECT 53.075 172.130 53.215 172.625 ;
        RECT 55.260 172.470 55.580 172.530 ;
        RECT 56.730 172.470 56.870 172.625 ;
        RECT 57.560 172.610 57.880 172.870 ;
        RECT 58.480 172.810 58.800 172.870 ;
        RECT 58.480 172.670 67.910 172.810 ;
        RECT 58.480 172.610 58.800 172.670 ;
        RECT 58.940 172.470 59.260 172.530 ;
        RECT 55.260 172.330 59.260 172.470 ;
        RECT 55.260 172.270 55.580 172.330 ;
        RECT 58.940 172.270 59.260 172.330 ;
        RECT 59.400 172.470 59.720 172.530 ;
        RECT 60.795 172.470 61.085 172.515 ;
        RECT 59.400 172.330 61.085 172.470 ;
        RECT 59.400 172.270 59.720 172.330 ;
        RECT 60.795 172.285 61.085 172.330 ;
        RECT 64.920 172.270 65.240 172.530 ;
        RECT 50.660 171.990 53.215 172.130 ;
        RECT 53.420 172.130 53.740 172.190 ;
        RECT 55.720 172.130 56.040 172.190 ;
        RECT 67.770 172.130 67.910 172.670 ;
        RECT 68.140 172.610 68.460 172.870 ;
        RECT 69.060 172.855 69.380 172.870 ;
        RECT 68.890 172.625 69.380 172.855 ;
        RECT 69.060 172.610 69.380 172.625 ;
        RECT 70.440 172.810 70.760 172.870 ;
        RECT 73.215 172.810 73.505 172.855 ;
        RECT 76.420 172.810 76.740 172.870 ;
        RECT 70.440 172.670 76.740 172.810 ;
        RECT 70.440 172.610 70.760 172.670 ;
        RECT 73.215 172.625 73.505 172.670 ;
        RECT 76.420 172.610 76.740 172.670 ;
        RECT 76.895 172.810 77.185 172.855 ;
        RECT 79.640 172.810 79.960 172.870 ;
        RECT 76.895 172.670 79.960 172.810 ;
        RECT 80.190 172.810 80.330 173.010 ;
        RECT 80.575 172.965 80.865 173.195 ;
        RECT 82.030 173.150 82.170 173.305 ;
        RECT 83.780 173.290 84.100 173.550 ;
        RECT 84.700 173.490 85.020 173.550 ;
        RECT 90.680 173.490 91.000 173.550 ;
        RECT 84.700 173.350 91.000 173.490 ;
        RECT 84.700 173.290 85.020 173.350 ;
        RECT 90.680 173.290 91.000 173.350 ;
        RECT 91.140 173.490 91.460 173.550 ;
        RECT 91.615 173.490 91.905 173.535 ;
        RECT 91.140 173.350 91.905 173.490 ;
        RECT 91.140 173.290 91.460 173.350 ;
        RECT 91.615 173.305 91.905 173.350 ;
        RECT 92.520 173.490 92.840 173.550 ;
        RECT 92.520 173.350 94.130 173.490 ;
        RECT 92.520 173.290 92.840 173.350 ;
        RECT 83.335 173.150 83.625 173.195 ;
        RECT 85.160 173.150 85.480 173.210 ;
        RECT 90.770 173.150 90.910 173.290 ;
        RECT 93.455 173.150 93.745 173.195 ;
        RECT 82.030 173.010 83.090 173.150 ;
        RECT 81.020 172.855 81.340 172.870 ;
        RECT 81.020 172.810 81.585 172.855 ;
        RECT 80.190 172.670 81.585 172.810 ;
        RECT 76.895 172.625 77.185 172.670 ;
        RECT 79.640 172.610 79.960 172.670 ;
        RECT 81.020 172.625 81.585 172.670 ;
        RECT 81.940 172.810 82.260 172.870 ;
        RECT 82.415 172.810 82.705 172.855 ;
        RECT 81.940 172.670 82.705 172.810 ;
        RECT 82.950 172.810 83.090 173.010 ;
        RECT 83.335 173.010 85.480 173.150 ;
        RECT 83.335 172.965 83.625 173.010 ;
        RECT 85.160 172.950 85.480 173.010 ;
        RECT 85.710 173.010 89.530 173.150 ;
        RECT 90.770 173.010 93.745 173.150 ;
        RECT 93.990 173.150 94.130 173.350 ;
        RECT 95.280 173.290 95.600 173.550 ;
        RECT 95.740 173.490 96.060 173.550 ;
        RECT 100.800 173.490 101.120 173.550 ;
        RECT 104.940 173.490 105.260 173.550 ;
        RECT 109.540 173.490 109.860 173.550 ;
        RECT 95.740 173.350 100.570 173.490 ;
        RECT 95.740 173.290 96.060 173.350 ;
        RECT 93.990 173.010 99.190 173.150 ;
        RECT 84.240 172.810 84.560 172.870 ;
        RECT 85.710 172.855 85.850 173.010 ;
        RECT 89.390 172.870 89.530 173.010 ;
        RECT 93.455 172.965 93.745 173.010 ;
        RECT 82.950 172.670 84.560 172.810 ;
        RECT 81.020 172.610 81.340 172.625 ;
        RECT 81.940 172.610 82.260 172.670 ;
        RECT 82.415 172.625 82.705 172.670 ;
        RECT 84.240 172.610 84.560 172.670 ;
        RECT 84.715 172.625 85.005 172.855 ;
        RECT 85.635 172.625 85.925 172.855 ;
        RECT 86.095 172.625 86.385 172.855 ;
        RECT 69.980 172.470 70.300 172.530 ;
        RECT 84.790 172.470 84.930 172.625 ;
        RECT 69.980 172.330 75.960 172.470 ;
        RECT 69.980 172.270 70.300 172.330 ;
        RECT 53.420 171.990 65.610 172.130 ;
        RECT 67.770 171.990 73.430 172.130 ;
        RECT 50.660 171.930 50.980 171.990 ;
        RECT 53.420 171.930 53.740 171.990 ;
        RECT 55.720 171.930 56.040 171.990 ;
        RECT 65.470 171.850 65.610 171.990 ;
        RECT 48.375 171.650 49.050 171.790 ;
        RECT 29.515 171.605 29.805 171.650 ;
        RECT 29.960 171.590 30.280 171.650 ;
        RECT 48.375 171.605 48.665 171.650 ;
        RECT 53.880 171.590 54.200 171.850 ;
        RECT 62.620 171.790 62.940 171.850 ;
        RECT 64.015 171.790 64.305 171.835 ;
        RECT 62.620 171.650 64.305 171.790 ;
        RECT 62.620 171.590 62.940 171.650 ;
        RECT 64.015 171.605 64.305 171.650 ;
        RECT 65.380 171.590 65.700 171.850 ;
        RECT 67.680 171.590 68.000 171.850 ;
        RECT 69.535 171.790 69.825 171.835 ;
        RECT 70.900 171.790 71.220 171.850 ;
        RECT 69.535 171.650 71.220 171.790 ;
        RECT 73.290 171.790 73.430 171.990 ;
        RECT 73.660 171.930 73.980 172.190 ;
        RECT 75.820 172.130 75.960 172.330 ;
        RECT 79.730 172.330 84.930 172.470 ;
        RECT 86.170 172.470 86.310 172.625 ;
        RECT 87.000 172.610 87.320 172.870 ;
        RECT 89.300 172.610 89.620 172.870 ;
        RECT 89.760 172.810 90.080 172.870 ;
        RECT 90.235 172.810 90.525 172.855 ;
        RECT 89.760 172.670 90.525 172.810 ;
        RECT 89.760 172.610 90.080 172.670 ;
        RECT 90.235 172.625 90.525 172.670 ;
        RECT 88.380 172.470 88.700 172.530 ;
        RECT 88.855 172.470 89.145 172.515 ;
        RECT 86.170 172.330 89.145 172.470 ;
        RECT 90.310 172.470 90.450 172.625 ;
        RECT 91.140 172.610 91.460 172.870 ;
        RECT 92.060 172.610 92.380 172.870 ;
        RECT 92.150 172.470 92.290 172.610 ;
        RECT 92.980 172.470 93.300 172.530 ;
        RECT 90.310 172.330 93.300 172.470 ;
        RECT 93.530 172.470 93.670 172.965 ;
        RECT 93.900 172.610 94.220 172.870 ;
        RECT 94.360 172.610 94.680 172.870 ;
        RECT 98.055 172.810 98.345 172.855 ;
        RECT 95.370 172.670 98.345 172.810 ;
        RECT 94.820 172.470 95.140 172.530 ;
        RECT 95.370 172.470 95.510 172.670 ;
        RECT 98.055 172.625 98.345 172.670 ;
        RECT 93.530 172.330 95.510 172.470 ;
        RECT 95.740 172.470 96.060 172.530 ;
        RECT 97.135 172.470 97.425 172.515 ;
        RECT 95.740 172.330 97.425 172.470 ;
        RECT 79.730 172.175 79.870 172.330 ;
        RECT 88.380 172.270 88.700 172.330 ;
        RECT 88.855 172.285 89.145 172.330 ;
        RECT 92.980 172.270 93.300 172.330 ;
        RECT 94.820 172.270 95.140 172.330 ;
        RECT 95.740 172.270 96.060 172.330 ;
        RECT 97.135 172.285 97.425 172.330 ;
        RECT 97.595 172.285 97.885 172.515 ;
        RECT 98.515 172.285 98.805 172.515 ;
        RECT 99.050 172.470 99.190 173.010 ;
        RECT 100.430 172.855 100.570 173.350 ;
        RECT 100.800 173.350 109.860 173.490 ;
        RECT 100.800 173.290 101.120 173.350 ;
        RECT 104.940 173.290 105.260 173.350 ;
        RECT 109.540 173.290 109.860 173.350 ;
        RECT 110.475 173.490 110.765 173.535 ;
        RECT 111.380 173.490 111.700 173.550 ;
        RECT 110.475 173.350 111.700 173.490 ;
        RECT 110.475 173.305 110.765 173.350 ;
        RECT 111.380 173.290 111.700 173.350 ;
        RECT 112.850 173.350 118.970 173.490 ;
        RECT 100.890 173.150 101.030 173.290 ;
        RECT 102.655 173.150 102.945 173.195 ;
        RECT 103.100 173.150 103.420 173.210 ;
        RECT 110.920 173.150 111.240 173.210 ;
        RECT 100.890 173.010 101.950 173.150 ;
        RECT 100.355 172.625 100.645 172.855 ;
        RECT 100.800 172.610 101.120 172.870 ;
        RECT 101.810 172.855 101.950 173.010 ;
        RECT 102.655 173.010 103.420 173.150 ;
        RECT 102.655 172.965 102.945 173.010 ;
        RECT 103.100 172.950 103.420 173.010 ;
        RECT 109.170 173.010 111.240 173.150 ;
        RECT 101.735 172.625 102.025 172.855 ;
        RECT 102.270 172.670 105.170 172.810 ;
        RECT 102.270 172.470 102.410 172.670 ;
        RECT 99.050 172.330 102.410 172.470 ;
        RECT 102.640 172.470 102.960 172.530 ;
        RECT 104.480 172.470 104.800 172.530 ;
        RECT 102.640 172.330 104.800 172.470 ;
        RECT 105.030 172.470 105.170 172.670 ;
        RECT 105.400 172.610 105.720 172.870 ;
        RECT 109.170 172.855 109.310 173.010 ;
        RECT 110.920 172.950 111.240 173.010 ;
        RECT 106.795 172.625 107.085 172.855 ;
        RECT 109.095 172.625 109.385 172.855 ;
        RECT 109.540 172.810 109.860 172.870 ;
        RECT 111.395 172.810 111.685 172.855 ;
        RECT 112.850 172.810 112.990 173.350 ;
        RECT 118.830 173.150 118.970 173.350 ;
        RECT 120.580 173.290 120.900 173.550 ;
        RECT 121.960 173.290 122.280 173.550 ;
        RECT 125.655 173.490 125.945 173.535 ;
        RECT 127.825 173.490 128.115 173.535 ;
        RECT 122.510 173.350 128.115 173.490 ;
        RECT 120.670 173.150 120.810 173.290 ;
        RECT 122.510 173.150 122.650 173.350 ;
        RECT 125.655 173.305 125.945 173.350 ;
        RECT 127.825 173.305 128.115 173.350 ;
        RECT 136.220 173.290 136.540 173.550 ;
        RECT 126.100 173.150 126.420 173.210 ;
        RECT 126.575 173.150 126.865 173.195 ;
        RECT 118.830 173.010 119.430 173.150 ;
        RECT 120.670 173.010 122.650 173.150 ;
        RECT 122.970 173.010 126.865 173.150 ;
        RECT 109.540 172.670 112.990 172.810 ;
        RECT 113.220 172.810 113.540 172.870 ;
        RECT 113.695 172.810 113.985 172.855 ;
        RECT 117.835 172.810 118.125 172.855 ;
        RECT 118.740 172.810 119.060 172.870 ;
        RECT 119.290 172.855 119.430 173.010 ;
        RECT 113.220 172.670 118.125 172.810 ;
        RECT 106.870 172.470 107.010 172.625 ;
        RECT 109.540 172.610 109.860 172.670 ;
        RECT 111.395 172.625 111.685 172.670 ;
        RECT 113.220 172.610 113.540 172.670 ;
        RECT 113.695 172.625 113.985 172.670 ;
        RECT 117.835 172.625 118.125 172.670 ;
        RECT 118.370 172.670 119.060 172.810 ;
        RECT 105.030 172.330 107.010 172.470 ;
        RECT 108.620 172.470 108.940 172.530 ;
        RECT 112.315 172.470 112.605 172.515 ;
        RECT 108.620 172.330 115.290 172.470 ;
        RECT 75.820 171.990 79.410 172.130 ;
        RECT 78.720 171.790 79.040 171.850 ;
        RECT 73.290 171.650 79.040 171.790 ;
        RECT 79.270 171.790 79.410 171.990 ;
        RECT 79.655 171.945 79.945 172.175 ;
        RECT 80.560 172.130 80.880 172.190 ;
        RECT 81.940 172.130 82.260 172.190 ;
        RECT 84.240 172.130 84.560 172.190 ;
        RECT 90.220 172.130 90.540 172.190 ;
        RECT 92.535 172.130 92.825 172.175 ;
        RECT 93.440 172.130 93.760 172.190 ;
        RECT 97.670 172.130 97.810 172.285 ;
        RECT 80.560 171.990 84.560 172.130 ;
        RECT 80.560 171.930 80.880 171.990 ;
        RECT 81.940 171.930 82.260 171.990 ;
        RECT 84.240 171.930 84.560 171.990 ;
        RECT 87.550 171.990 89.990 172.130 ;
        RECT 87.550 171.790 87.690 171.990 ;
        RECT 79.270 171.650 87.690 171.790 ;
        RECT 69.535 171.605 69.825 171.650 ;
        RECT 70.900 171.590 71.220 171.650 ;
        RECT 78.720 171.590 79.040 171.650 ;
        RECT 87.920 171.590 88.240 171.850 ;
        RECT 89.850 171.790 89.990 171.990 ;
        RECT 90.220 171.990 97.810 172.130 ;
        RECT 98.590 172.130 98.730 172.285 ;
        RECT 102.640 172.270 102.960 172.330 ;
        RECT 104.480 172.270 104.800 172.330 ;
        RECT 108.620 172.270 108.940 172.330 ;
        RECT 112.315 172.285 112.605 172.330 ;
        RECT 100.800 172.130 101.120 172.190 ;
        RECT 98.590 171.990 101.120 172.130 ;
        RECT 90.220 171.930 90.540 171.990 ;
        RECT 92.535 171.945 92.825 171.990 ;
        RECT 93.440 171.930 93.760 171.990 ;
        RECT 100.800 171.930 101.120 171.990 ;
        RECT 101.260 171.930 101.580 172.190 ;
        RECT 103.100 172.130 103.420 172.190 ;
        RECT 104.955 172.130 105.245 172.175 ;
        RECT 105.400 172.130 105.720 172.190 ;
        RECT 103.100 171.990 105.720 172.130 ;
        RECT 103.100 171.930 103.420 171.990 ;
        RECT 104.955 171.945 105.245 171.990 ;
        RECT 105.400 171.930 105.720 171.990 ;
        RECT 110.015 172.130 110.305 172.175 ;
        RECT 112.760 172.130 113.080 172.190 ;
        RECT 115.150 172.130 115.290 172.330 ;
        RECT 116.900 172.270 117.220 172.530 ;
        RECT 118.370 172.130 118.510 172.670 ;
        RECT 118.740 172.610 119.060 172.670 ;
        RECT 119.215 172.810 119.505 172.855 ;
        RECT 120.120 172.810 120.440 172.870 ;
        RECT 119.215 172.670 120.440 172.810 ;
        RECT 119.215 172.625 119.505 172.670 ;
        RECT 120.120 172.610 120.440 172.670 ;
        RECT 122.420 172.610 122.740 172.870 ;
        RECT 122.970 172.855 123.110 173.010 ;
        RECT 126.100 172.950 126.420 173.010 ;
        RECT 126.575 172.965 126.865 173.010 ;
        RECT 128.400 173.150 128.720 173.210 ;
        RECT 128.875 173.150 129.165 173.195 ;
        RECT 128.400 173.010 129.165 173.150 ;
        RECT 128.400 172.950 128.720 173.010 ;
        RECT 128.875 172.965 129.165 173.010 ;
        RECT 122.895 172.625 123.185 172.855 ;
        RECT 124.275 172.810 124.565 172.855 ;
        RECT 136.310 172.810 136.450 173.290 ;
        RECT 124.275 172.670 136.450 172.810 ;
        RECT 124.275 172.625 124.565 172.670 ;
        RECT 120.580 172.470 120.900 172.530 ;
        RECT 118.830 172.330 120.900 172.470 ;
        RECT 118.830 172.190 118.970 172.330 ;
        RECT 120.580 172.270 120.900 172.330 ;
        RECT 121.040 172.270 121.360 172.530 ;
        RECT 123.815 172.470 124.105 172.515 ;
        RECT 132.080 172.470 132.400 172.530 ;
        RECT 123.815 172.330 132.400 172.470 ;
        RECT 123.815 172.285 124.105 172.330 ;
        RECT 132.080 172.270 132.400 172.330 ;
        RECT 134.380 172.470 134.700 172.530 ;
        RECT 137.615 172.470 137.905 172.515 ;
        RECT 134.380 172.330 137.905 172.470 ;
        RECT 134.380 172.270 134.700 172.330 ;
        RECT 137.615 172.285 137.905 172.330 ;
        RECT 110.015 171.990 113.080 172.130 ;
        RECT 110.015 171.945 110.305 171.990 ;
        RECT 112.760 171.930 113.080 171.990 ;
        RECT 113.770 171.990 114.830 172.130 ;
        RECT 115.150 171.990 118.510 172.130 ;
        RECT 98.960 171.790 99.280 171.850 ;
        RECT 89.850 171.650 99.280 171.790 ;
        RECT 98.960 171.590 99.280 171.650 ;
        RECT 99.435 171.790 99.725 171.835 ;
        RECT 108.620 171.790 108.940 171.850 ;
        RECT 99.435 171.650 108.940 171.790 ;
        RECT 99.435 171.605 99.725 171.650 ;
        RECT 108.620 171.590 108.940 171.650 ;
        RECT 109.095 171.790 109.385 171.835 ;
        RECT 110.460 171.790 110.780 171.850 ;
        RECT 109.095 171.650 110.780 171.790 ;
        RECT 109.095 171.605 109.385 171.650 ;
        RECT 110.460 171.590 110.780 171.650 ;
        RECT 111.380 171.790 111.700 171.850 ;
        RECT 113.770 171.790 113.910 171.990 ;
        RECT 111.380 171.650 113.910 171.790 ;
        RECT 111.380 171.590 111.700 171.650 ;
        RECT 114.140 171.590 114.460 171.850 ;
        RECT 114.690 171.790 114.830 171.990 ;
        RECT 118.740 171.930 119.060 172.190 ;
        RECT 120.135 172.130 120.425 172.175 ;
        RECT 121.130 172.130 121.270 172.270 ;
        RECT 120.135 171.990 121.270 172.130 ;
        RECT 120.135 171.945 120.425 171.990 ;
        RECT 117.820 171.790 118.140 171.850 ;
        RECT 114.690 171.650 118.140 171.790 ;
        RECT 121.130 171.790 121.270 171.990 ;
        RECT 125.180 172.130 125.500 172.190 ;
        RECT 127.035 172.130 127.325 172.175 ;
        RECT 125.180 171.990 127.325 172.130 ;
        RECT 125.180 171.930 125.500 171.990 ;
        RECT 127.035 171.945 127.325 171.990 ;
        RECT 125.655 171.790 125.945 171.835 ;
        RECT 127.955 171.790 128.245 171.835 ;
        RECT 121.130 171.650 128.245 171.790 ;
        RECT 117.820 171.590 118.140 171.650 ;
        RECT 125.655 171.605 125.945 171.650 ;
        RECT 127.955 171.605 128.245 171.650 ;
        RECT 134.840 171.590 135.160 171.850 ;
        RECT 2.750 170.970 158.230 171.450 ;
        RECT 14.780 170.770 15.100 170.830 ;
        RECT 17.080 170.770 17.400 170.830 ;
        RECT 14.780 170.630 17.400 170.770 ;
        RECT 14.780 170.570 15.100 170.630 ;
        RECT 17.080 170.570 17.400 170.630 ;
        RECT 18.000 170.770 18.320 170.830 ;
        RECT 22.600 170.770 22.920 170.830 ;
        RECT 18.000 170.630 22.920 170.770 ;
        RECT 18.000 170.570 18.320 170.630 ;
        RECT 22.600 170.570 22.920 170.630 ;
        RECT 23.980 170.770 24.300 170.830 ;
        RECT 25.145 170.770 25.435 170.815 ;
        RECT 23.980 170.630 25.435 170.770 ;
        RECT 23.980 170.570 24.300 170.630 ;
        RECT 25.145 170.585 25.435 170.630 ;
        RECT 38.700 170.570 39.020 170.830 ;
        RECT 45.600 170.570 45.920 170.830 ;
        RECT 47.440 170.570 47.760 170.830 ;
        RECT 47.990 170.630 53.190 170.770 ;
        RECT 5.085 170.430 5.375 170.475 ;
        RECT 6.975 170.430 7.265 170.475 ;
        RECT 10.095 170.430 10.385 170.475 ;
        RECT 5.085 170.290 10.385 170.430 ;
        RECT 5.085 170.245 5.375 170.290 ;
        RECT 6.975 170.245 7.265 170.290 ;
        RECT 10.095 170.245 10.385 170.290 ;
        RECT 15.255 170.245 15.545 170.475 ;
        RECT 16.640 170.430 16.930 170.475 ;
        RECT 18.500 170.430 18.790 170.475 ;
        RECT 21.280 170.430 21.570 170.475 ;
        RECT 16.640 170.290 21.570 170.430 ;
        RECT 16.640 170.245 16.930 170.290 ;
        RECT 18.500 170.245 18.790 170.290 ;
        RECT 21.280 170.245 21.570 170.290 ;
        RECT 22.140 170.430 22.460 170.490 ;
        RECT 24.070 170.430 24.210 170.570 ;
        RECT 22.140 170.290 24.210 170.430 ;
        RECT 29.465 170.430 29.755 170.475 ;
        RECT 31.355 170.430 31.645 170.475 ;
        RECT 34.475 170.430 34.765 170.475 ;
        RECT 29.465 170.290 34.765 170.430 ;
        RECT 4.200 169.550 4.520 169.810 ;
        RECT 4.680 169.750 4.970 169.795 ;
        RECT 6.515 169.750 6.805 169.795 ;
        RECT 10.095 169.750 10.385 169.795 ;
        RECT 4.680 169.610 10.385 169.750 ;
        RECT 4.680 169.565 4.970 169.610 ;
        RECT 6.515 169.565 6.805 169.610 ;
        RECT 10.095 169.565 10.385 169.610 ;
        RECT 5.580 169.210 5.900 169.470 ;
        RECT 7.875 169.410 8.525 169.455 ;
        RECT 8.800 169.410 9.120 169.470 ;
        RECT 11.175 169.455 11.465 169.770 ;
        RECT 14.320 169.550 14.640 169.810 ;
        RECT 15.330 169.750 15.470 170.245 ;
        RECT 22.140 170.230 22.460 170.290 ;
        RECT 29.465 170.245 29.755 170.290 ;
        RECT 31.355 170.245 31.645 170.290 ;
        RECT 34.475 170.245 34.765 170.290 ;
        RECT 36.860 170.430 37.180 170.490 ;
        RECT 37.335 170.430 37.625 170.475 ;
        RECT 47.990 170.430 48.130 170.630 ;
        RECT 53.050 170.490 53.190 170.630 ;
        RECT 53.880 170.570 54.200 170.830 ;
        RECT 54.800 170.570 55.120 170.830 ;
        RECT 56.655 170.770 56.945 170.815 ;
        RECT 58.020 170.770 58.340 170.830 ;
        RECT 56.655 170.630 58.340 170.770 ;
        RECT 56.655 170.585 56.945 170.630 ;
        RECT 58.020 170.570 58.340 170.630 ;
        RECT 59.400 170.770 59.720 170.830 ;
        RECT 61.255 170.770 61.545 170.815 ;
        RECT 59.400 170.630 61.545 170.770 ;
        RECT 59.400 170.570 59.720 170.630 ;
        RECT 61.255 170.585 61.545 170.630 ;
        RECT 64.920 170.770 65.240 170.830 ;
        RECT 66.775 170.770 67.065 170.815 ;
        RECT 74.580 170.770 74.900 170.830 ;
        RECT 76.435 170.770 76.725 170.815 ;
        RECT 64.920 170.630 67.065 170.770 ;
        RECT 64.920 170.570 65.240 170.630 ;
        RECT 66.775 170.585 67.065 170.630 ;
        RECT 67.310 170.630 76.725 170.770 ;
        RECT 36.860 170.290 48.130 170.430 ;
        RECT 36.860 170.230 37.180 170.290 ;
        RECT 37.335 170.245 37.625 170.290 ;
        RECT 50.660 170.230 50.980 170.490 ;
        RECT 52.515 170.245 52.805 170.475 ;
        RECT 16.175 170.090 16.465 170.135 ;
        RECT 17.540 170.090 17.860 170.150 ;
        RECT 16.175 169.950 28.810 170.090 ;
        RECT 16.175 169.905 16.465 169.950 ;
        RECT 17.540 169.890 17.860 169.950 ;
        RECT 28.670 169.795 28.810 169.950 ;
        RECT 29.960 169.890 30.280 170.150 ;
        RECT 31.800 170.090 32.120 170.150 ;
        RECT 42.395 170.090 42.685 170.135 ;
        RECT 45.140 170.090 45.460 170.150 ;
        RECT 31.800 169.950 45.460 170.090 ;
        RECT 31.800 169.890 32.120 169.950 ;
        RECT 42.395 169.905 42.685 169.950 ;
        RECT 45.140 169.890 45.460 169.950 ;
        RECT 45.690 169.950 49.510 170.090 ;
        RECT 18.015 169.750 18.305 169.795 ;
        RECT 21.280 169.750 21.570 169.795 ;
        RECT 15.330 169.610 18.305 169.750 ;
        RECT 18.015 169.565 18.305 169.610 ;
        RECT 19.035 169.610 21.570 169.750 ;
        RECT 11.175 169.410 11.765 169.455 ;
        RECT 7.875 169.270 11.765 169.410 ;
        RECT 7.875 169.225 8.525 169.270 ;
        RECT 8.800 169.210 9.120 169.270 ;
        RECT 11.475 169.225 11.765 169.270 ;
        RECT 14.780 169.210 15.100 169.470 ;
        RECT 19.035 169.455 19.250 169.610 ;
        RECT 21.280 169.565 21.570 169.610 ;
        RECT 28.595 169.565 28.885 169.795 ;
        RECT 29.060 169.750 29.350 169.795 ;
        RECT 30.895 169.750 31.185 169.795 ;
        RECT 34.475 169.750 34.765 169.795 ;
        RECT 29.060 169.610 34.765 169.750 ;
        RECT 29.060 169.565 29.350 169.610 ;
        RECT 30.895 169.565 31.185 169.610 ;
        RECT 34.475 169.565 34.765 169.610 ;
        RECT 17.100 169.410 17.390 169.455 ;
        RECT 18.960 169.410 19.250 169.455 ;
        RECT 19.880 169.410 20.170 169.455 ;
        RECT 23.140 169.410 23.430 169.455 ;
        RECT 17.100 169.270 19.250 169.410 ;
        RECT 17.100 169.225 17.390 169.270 ;
        RECT 18.960 169.225 19.250 169.270 ;
        RECT 19.470 169.270 23.430 169.410 ;
        RECT 28.670 169.410 28.810 169.565 ;
        RECT 32.720 169.455 33.040 169.470 ;
        RECT 32.255 169.410 33.040 169.455 ;
        RECT 35.555 169.455 35.845 169.770 ;
        RECT 39.620 169.550 39.940 169.810 ;
        RECT 40.095 169.750 40.385 169.795 ;
        RECT 44.220 169.750 44.540 169.810 ;
        RECT 40.095 169.610 44.540 169.750 ;
        RECT 40.095 169.565 40.385 169.610 ;
        RECT 44.220 169.550 44.540 169.610 ;
        RECT 35.555 169.410 36.145 169.455 ;
        RECT 43.315 169.410 43.605 169.455 ;
        RECT 28.670 169.270 29.270 169.410 ;
        RECT 12.940 168.870 13.260 169.130 ;
        RECT 14.870 169.070 15.010 169.210 ;
        RECT 19.470 169.070 19.610 169.270 ;
        RECT 19.880 169.225 20.170 169.270 ;
        RECT 23.140 169.225 23.430 169.270 ;
        RECT 29.130 169.130 29.270 169.270 ;
        RECT 32.255 169.270 36.145 169.410 ;
        RECT 32.255 169.225 33.040 169.270 ;
        RECT 35.855 169.225 36.145 169.270 ;
        RECT 37.870 169.270 43.605 169.410 ;
        RECT 32.720 169.210 33.040 169.225 ;
        RECT 24.440 169.070 24.760 169.130 ;
        RECT 14.870 168.930 24.760 169.070 ;
        RECT 24.440 168.870 24.760 168.930 ;
        RECT 29.040 168.870 29.360 169.130 ;
        RECT 34.100 169.070 34.420 169.130 ;
        RECT 37.870 169.070 38.010 169.270 ;
        RECT 43.315 169.225 43.605 169.270 ;
        RECT 43.760 169.410 44.080 169.470 ;
        RECT 45.690 169.410 45.830 169.950 ;
        RECT 49.370 169.810 49.510 169.950 ;
        RECT 46.075 169.565 46.365 169.795 ;
        RECT 46.520 169.750 46.840 169.810 ;
        RECT 47.455 169.750 47.745 169.795 ;
        RECT 46.520 169.610 47.745 169.750 ;
        RECT 43.760 169.270 45.830 169.410 ;
        RECT 46.150 169.410 46.290 169.565 ;
        RECT 46.520 169.550 46.840 169.610 ;
        RECT 47.455 169.565 47.745 169.610 ;
        RECT 47.900 169.550 48.220 169.810 ;
        RECT 48.375 169.565 48.665 169.795 ;
        RECT 48.450 169.410 48.590 169.565 ;
        RECT 49.280 169.550 49.600 169.810 ;
        RECT 49.755 169.750 50.045 169.795 ;
        RECT 50.750 169.750 50.890 170.230 ;
        RECT 52.590 170.090 52.730 170.245 ;
        RECT 52.960 170.230 53.280 170.490 ;
        RECT 53.970 170.430 54.110 170.570 ;
        RECT 65.380 170.430 65.700 170.490 ;
        RECT 67.310 170.430 67.450 170.630 ;
        RECT 74.580 170.570 74.900 170.630 ;
        RECT 76.435 170.585 76.725 170.630 ;
        RECT 77.355 170.770 77.645 170.815 ;
        RECT 77.800 170.770 78.120 170.830 ;
        RECT 87.935 170.770 88.225 170.815 ;
        RECT 88.840 170.770 89.160 170.830 ;
        RECT 77.355 170.630 78.120 170.770 ;
        RECT 77.355 170.585 77.645 170.630 ;
        RECT 77.800 170.570 78.120 170.630 ;
        RECT 78.350 170.630 87.690 170.770 ;
        RECT 53.970 170.290 57.790 170.430 ;
        RECT 55.275 170.090 55.565 170.135 ;
        RECT 56.180 170.090 56.500 170.150 ;
        RECT 52.130 169.950 52.730 170.090 ;
        RECT 53.970 169.950 55.030 170.090 ;
        RECT 49.755 169.610 50.890 169.750 ;
        RECT 49.755 169.565 50.045 169.610 ;
        RECT 51.120 169.550 51.440 169.810 ;
        RECT 52.130 169.795 52.270 169.950 ;
        RECT 52.055 169.565 52.345 169.795 ;
        RECT 52.515 169.750 52.805 169.795 ;
        RECT 53.420 169.750 53.740 169.810 ;
        RECT 53.970 169.795 54.110 169.950 ;
        RECT 54.890 169.810 55.030 169.950 ;
        RECT 55.275 169.950 56.500 170.090 ;
        RECT 55.275 169.905 55.565 169.950 ;
        RECT 56.180 169.890 56.500 169.950 ;
        RECT 52.515 169.610 53.740 169.750 ;
        RECT 52.515 169.565 52.805 169.610 ;
        RECT 53.420 169.550 53.740 169.610 ;
        RECT 53.895 169.565 54.185 169.795 ;
        RECT 54.340 169.550 54.660 169.810 ;
        RECT 54.800 169.550 55.120 169.810 ;
        RECT 55.735 169.750 56.025 169.795 ;
        RECT 56.640 169.750 56.960 169.810 ;
        RECT 57.650 169.795 57.790 170.290 ;
        RECT 59.490 170.290 64.690 170.430 ;
        RECT 58.940 170.090 59.260 170.150 ;
        RECT 59.490 170.090 59.630 170.290 ;
        RECT 64.550 170.150 64.690 170.290 ;
        RECT 65.010 170.290 67.450 170.430 ;
        RECT 63.540 170.090 63.860 170.150 ;
        RECT 58.940 169.950 59.630 170.090 ;
        RECT 60.410 169.950 63.860 170.090 ;
        RECT 58.940 169.890 59.260 169.950 ;
        RECT 55.735 169.610 56.960 169.750 ;
        RECT 55.735 169.565 56.025 169.610 ;
        RECT 56.640 169.550 56.960 169.610 ;
        RECT 57.575 169.565 57.865 169.795 ;
        RECT 58.480 169.550 58.800 169.810 ;
        RECT 59.400 169.550 59.720 169.810 ;
        RECT 60.410 169.795 60.550 169.950 ;
        RECT 63.540 169.890 63.860 169.950 ;
        RECT 64.460 169.890 64.780 170.150 ;
        RECT 60.335 169.565 60.625 169.795 ;
        RECT 63.095 169.565 63.385 169.795 ;
        RECT 51.595 169.410 51.885 169.455 ;
        RECT 63.170 169.410 63.310 169.565 ;
        RECT 46.150 169.270 47.210 169.410 ;
        RECT 48.450 169.270 51.885 169.410 ;
        RECT 43.760 169.210 44.080 169.270 ;
        RECT 34.100 168.930 38.010 169.070 ;
        RECT 41.015 169.070 41.305 169.115 ;
        RECT 45.140 169.070 45.460 169.130 ;
        RECT 41.015 168.930 45.460 169.070 ;
        RECT 34.100 168.870 34.420 168.930 ;
        RECT 41.015 168.885 41.305 168.930 ;
        RECT 45.140 168.870 45.460 168.930 ;
        RECT 46.060 169.070 46.380 169.130 ;
        RECT 46.535 169.070 46.825 169.115 ;
        RECT 46.060 168.930 46.825 169.070 ;
        RECT 47.070 169.070 47.210 169.270 ;
        RECT 51.595 169.225 51.885 169.270 ;
        RECT 53.050 169.270 63.310 169.410 ;
        RECT 63.645 169.410 63.785 169.890 ;
        RECT 64.000 169.550 64.320 169.810 ;
        RECT 65.010 169.795 65.150 170.290 ;
        RECT 65.380 170.230 65.700 170.290 ;
        RECT 67.680 170.230 68.000 170.490 ;
        RECT 68.565 170.430 68.855 170.475 ;
        RECT 70.455 170.430 70.745 170.475 ;
        RECT 73.575 170.430 73.865 170.475 ;
        RECT 68.565 170.290 73.865 170.430 ;
        RECT 68.565 170.245 68.855 170.290 ;
        RECT 70.455 170.245 70.745 170.290 ;
        RECT 73.575 170.245 73.865 170.290 ;
        RECT 67.770 170.090 67.910 170.230 ;
        RECT 69.075 170.090 69.365 170.135 ;
        RECT 67.770 169.950 69.365 170.090 ;
        RECT 69.075 169.905 69.365 169.950 ;
        RECT 70.900 170.090 71.220 170.150 ;
        RECT 78.350 170.090 78.490 170.630 ;
        RECT 81.020 170.430 81.340 170.490 ;
        RECT 83.795 170.430 84.085 170.475 ;
        RECT 87.550 170.430 87.690 170.630 ;
        RECT 87.935 170.630 89.160 170.770 ;
        RECT 87.935 170.585 88.225 170.630 ;
        RECT 88.840 170.570 89.160 170.630 ;
        RECT 89.300 170.570 89.620 170.830 ;
        RECT 90.680 170.770 91.000 170.830 ;
        RECT 91.615 170.770 91.905 170.815 ;
        RECT 101.260 170.770 101.580 170.830 ;
        RECT 105.875 170.770 106.165 170.815 ;
        RECT 106.780 170.770 107.100 170.830 ;
        RECT 90.680 170.630 91.905 170.770 ;
        RECT 90.680 170.570 91.000 170.630 ;
        RECT 91.615 170.585 91.905 170.630 ;
        RECT 92.150 170.630 105.170 170.770 ;
        RECT 92.150 170.430 92.290 170.630 ;
        RECT 101.260 170.570 101.580 170.630 ;
        RECT 100.800 170.430 101.120 170.490 ;
        RECT 81.020 170.290 87.230 170.430 ;
        RECT 87.550 170.290 92.290 170.430 ;
        RECT 93.990 170.290 101.120 170.430 ;
        RECT 81.020 170.230 81.340 170.290 ;
        RECT 83.795 170.245 84.085 170.290 ;
        RECT 70.900 169.950 78.490 170.090 ;
        RECT 70.900 169.890 71.220 169.950 ;
        RECT 64.935 169.565 65.225 169.795 ;
        RECT 65.855 169.565 66.145 169.795 ;
        RECT 65.930 169.410 66.070 169.565 ;
        RECT 67.680 169.550 68.000 169.810 ;
        RECT 68.160 169.750 68.450 169.795 ;
        RECT 69.995 169.750 70.285 169.795 ;
        RECT 73.575 169.750 73.865 169.795 ;
        RECT 68.160 169.610 73.865 169.750 ;
        RECT 68.160 169.565 68.450 169.610 ;
        RECT 69.995 169.565 70.285 169.610 ;
        RECT 73.575 169.565 73.865 169.610 ;
        RECT 63.645 169.270 66.070 169.410 ;
        RECT 49.740 169.070 50.060 169.130 ;
        RECT 47.070 168.930 50.060 169.070 ;
        RECT 46.060 168.870 46.380 168.930 ;
        RECT 46.535 168.885 46.825 168.930 ;
        RECT 49.740 168.870 50.060 168.930 ;
        RECT 50.675 169.070 50.965 169.115 ;
        RECT 53.050 169.070 53.190 169.270 ;
        RECT 50.675 168.930 53.190 169.070 ;
        RECT 53.435 169.070 53.725 169.115 ;
        RECT 57.560 169.070 57.880 169.130 ;
        RECT 53.435 168.930 57.880 169.070 ;
        RECT 65.930 169.070 66.070 169.270 ;
        RECT 69.060 169.410 69.380 169.470 ;
        RECT 74.655 169.455 74.945 169.770 ;
        RECT 76.420 169.750 76.740 169.810 ;
        RECT 80.560 169.750 80.880 169.810 ;
        RECT 76.420 169.610 80.880 169.750 ;
        RECT 81.110 169.750 81.250 170.230 ;
        RECT 82.415 170.090 82.705 170.135 ;
        RECT 83.320 170.090 83.640 170.150 ;
        RECT 82.415 169.950 83.640 170.090 ;
        RECT 82.415 169.905 82.705 169.950 ;
        RECT 83.320 169.890 83.640 169.950 ;
        RECT 84.240 170.090 84.560 170.150 ;
        RECT 87.090 170.090 87.230 170.290 ;
        RECT 93.990 170.150 94.130 170.290 ;
        RECT 100.800 170.230 101.120 170.290 ;
        RECT 102.180 170.230 102.500 170.490 ;
        RECT 102.655 170.430 102.945 170.475 ;
        RECT 103.560 170.430 103.880 170.490 ;
        RECT 102.655 170.290 103.880 170.430 ;
        RECT 102.655 170.245 102.945 170.290 ;
        RECT 103.560 170.230 103.880 170.290 ;
        RECT 104.020 170.230 104.340 170.490 ;
        RECT 104.495 170.430 104.785 170.475 ;
        RECT 105.030 170.430 105.170 170.630 ;
        RECT 105.875 170.630 107.100 170.770 ;
        RECT 105.875 170.585 106.165 170.630 ;
        RECT 106.780 170.570 107.100 170.630 ;
        RECT 107.240 170.570 107.560 170.830 ;
        RECT 112.760 170.770 113.080 170.830 ;
        RECT 117.360 170.770 117.680 170.830 ;
        RECT 112.760 170.630 117.680 170.770 ;
        RECT 112.760 170.570 113.080 170.630 ;
        RECT 117.360 170.570 117.680 170.630 ;
        RECT 117.820 170.770 118.140 170.830 ;
        RECT 119.675 170.770 119.965 170.815 ;
        RECT 117.820 170.630 119.965 170.770 ;
        RECT 117.820 170.570 118.140 170.630 ;
        RECT 119.675 170.585 119.965 170.630 ;
        RECT 120.120 170.770 120.440 170.830 ;
        RECT 122.895 170.770 123.185 170.815 ;
        RECT 120.120 170.630 123.185 170.770 ;
        RECT 120.120 170.570 120.440 170.630 ;
        RECT 122.895 170.585 123.185 170.630 ;
        RECT 133.705 170.770 133.995 170.815 ;
        RECT 134.380 170.770 134.700 170.830 ;
        RECT 133.705 170.630 134.700 170.770 ;
        RECT 133.705 170.585 133.995 170.630 ;
        RECT 134.380 170.570 134.700 170.630 ;
        RECT 134.840 170.570 135.160 170.830 ;
        RECT 111.380 170.430 111.700 170.490 ;
        RECT 104.495 170.290 111.700 170.430 ;
        RECT 104.495 170.245 104.785 170.290 ;
        RECT 111.380 170.230 111.700 170.290 ;
        RECT 125.200 170.430 125.490 170.475 ;
        RECT 127.060 170.430 127.350 170.475 ;
        RECT 129.840 170.430 130.130 170.475 ;
        RECT 125.200 170.290 130.130 170.430 ;
        RECT 125.200 170.245 125.490 170.290 ;
        RECT 127.060 170.245 127.350 170.290 ;
        RECT 129.840 170.245 130.130 170.290 ;
        RECT 90.220 170.090 90.540 170.150 ;
        RECT 93.455 170.090 93.745 170.135 ;
        RECT 93.900 170.090 94.220 170.150 ;
        RECT 97.580 170.090 97.900 170.150 ;
        RECT 99.435 170.090 99.725 170.135 ;
        RECT 102.270 170.090 102.410 170.230 ;
        RECT 84.240 169.950 86.770 170.090 ;
        RECT 87.090 169.950 90.540 170.090 ;
        RECT 84.240 169.890 84.560 169.950 ;
        RECT 81.495 169.750 81.785 169.795 ;
        RECT 81.110 169.610 81.785 169.750 ;
        RECT 76.420 169.550 76.740 169.610 ;
        RECT 71.355 169.410 72.005 169.455 ;
        RECT 74.655 169.410 75.245 169.455 ;
        RECT 77.800 169.410 78.120 169.470 ;
        RECT 78.810 169.455 78.950 169.610 ;
        RECT 80.560 169.550 80.880 169.610 ;
        RECT 81.495 169.565 81.785 169.610 ;
        RECT 82.875 169.750 83.165 169.795 ;
        RECT 83.780 169.750 84.100 169.810 ;
        RECT 86.630 169.795 86.770 169.950 ;
        RECT 88.930 169.795 89.070 169.950 ;
        RECT 90.220 169.890 90.540 169.950 ;
        RECT 92.150 169.950 94.220 170.090 ;
        RECT 85.175 169.750 85.465 169.795 ;
        RECT 82.875 169.610 85.465 169.750 ;
        RECT 82.875 169.565 83.165 169.610 ;
        RECT 69.060 169.270 75.245 169.410 ;
        RECT 69.060 169.210 69.380 169.270 ;
        RECT 71.355 169.225 72.005 169.270 ;
        RECT 74.955 169.225 75.245 169.270 ;
        RECT 75.590 169.270 78.120 169.410 ;
        RECT 75.590 169.070 75.730 169.270 ;
        RECT 77.800 169.210 78.120 169.270 ;
        RECT 78.735 169.225 79.025 169.455 ;
        RECT 80.115 169.410 80.405 169.455 ;
        RECT 82.950 169.410 83.090 169.565 ;
        RECT 83.780 169.550 84.100 169.610 ;
        RECT 85.175 169.565 85.465 169.610 ;
        RECT 86.555 169.750 86.845 169.795 ;
        RECT 86.555 169.610 88.610 169.750 ;
        RECT 86.555 169.565 86.845 169.610 ;
        RECT 80.115 169.270 83.090 169.410 ;
        RECT 84.240 169.410 84.560 169.470 ;
        RECT 88.470 169.410 88.610 169.610 ;
        RECT 88.855 169.565 89.145 169.795 ;
        RECT 89.775 169.750 90.065 169.795 ;
        RECT 91.600 169.750 91.920 169.810 ;
        RECT 89.775 169.610 91.920 169.750 ;
        RECT 89.775 169.565 90.065 169.610 ;
        RECT 91.600 169.550 91.920 169.610 ;
        RECT 92.150 169.410 92.290 169.950 ;
        RECT 93.455 169.905 93.745 169.950 ;
        RECT 93.900 169.890 94.220 169.950 ;
        RECT 94.450 169.950 95.510 170.090 ;
        RECT 94.450 169.810 94.590 169.950 ;
        RECT 92.520 169.550 92.840 169.810 ;
        RECT 94.360 169.550 94.680 169.810 ;
        RECT 95.370 169.795 95.510 169.950 ;
        RECT 97.580 169.950 98.270 170.090 ;
        RECT 97.580 169.890 97.900 169.950 ;
        RECT 94.835 169.565 95.125 169.795 ;
        RECT 95.295 169.750 95.585 169.795 ;
        RECT 98.130 169.750 98.270 169.950 ;
        RECT 99.435 169.950 102.410 170.090 ;
        RECT 99.435 169.905 99.725 169.950 ;
        RECT 99.895 169.750 100.185 169.795 ;
        RECT 95.295 169.610 97.810 169.750 ;
        RECT 98.130 169.610 100.185 169.750 ;
        RECT 95.295 169.565 95.585 169.610 ;
        RECT 84.240 169.270 87.230 169.410 ;
        RECT 88.470 169.270 92.290 169.410 ;
        RECT 93.440 169.410 93.760 169.470 ;
        RECT 94.910 169.410 95.050 169.565 ;
        RECT 93.440 169.270 95.050 169.410 ;
        RECT 80.115 169.225 80.405 169.270 ;
        RECT 84.240 169.210 84.560 169.270 ;
        RECT 65.930 168.930 75.730 169.070 ;
        RECT 76.880 169.070 77.200 169.130 ;
        RECT 78.275 169.070 78.565 169.115 ;
        RECT 76.880 168.930 78.565 169.070 ;
        RECT 50.675 168.885 50.965 168.930 ;
        RECT 53.435 168.885 53.725 168.930 ;
        RECT 57.560 168.870 57.880 168.930 ;
        RECT 76.880 168.870 77.200 168.930 ;
        RECT 78.275 168.885 78.565 168.930 ;
        RECT 79.180 168.870 79.500 169.130 ;
        RECT 79.640 169.070 79.960 169.130 ;
        RECT 80.575 169.070 80.865 169.115 ;
        RECT 82.400 169.070 82.720 169.130 ;
        RECT 79.640 168.930 82.720 169.070 ;
        RECT 79.640 168.870 79.960 168.930 ;
        RECT 80.575 168.885 80.865 168.930 ;
        RECT 82.400 168.870 82.720 168.930 ;
        RECT 84.700 169.070 85.020 169.130 ;
        RECT 87.090 169.115 87.230 169.270 ;
        RECT 93.440 169.210 93.760 169.270 ;
        RECT 86.095 169.070 86.385 169.115 ;
        RECT 84.700 168.930 86.385 169.070 ;
        RECT 84.700 168.870 85.020 168.930 ;
        RECT 86.095 168.885 86.385 168.930 ;
        RECT 87.015 169.070 87.305 169.115 ;
        RECT 92.060 169.070 92.380 169.130 ;
        RECT 87.015 168.930 92.380 169.070 ;
        RECT 94.910 169.070 95.050 169.270 ;
        RECT 96.660 169.410 96.980 169.470 ;
        RECT 97.135 169.410 97.425 169.455 ;
        RECT 96.660 169.270 97.425 169.410 ;
        RECT 97.670 169.410 97.810 169.610 ;
        RECT 99.895 169.565 100.185 169.610 ;
        RECT 101.720 169.550 102.040 169.810 ;
        RECT 102.180 169.750 102.500 169.810 ;
        RECT 104.110 169.795 104.250 170.230 ;
        RECT 110.920 170.090 111.240 170.150 ;
        RECT 124.735 170.090 125.025 170.135 ;
        RECT 134.930 170.090 135.070 170.570 ;
        RECT 135.265 170.430 135.555 170.475 ;
        RECT 137.155 170.430 137.445 170.475 ;
        RECT 140.275 170.430 140.565 170.475 ;
        RECT 135.265 170.290 140.565 170.430 ;
        RECT 135.265 170.245 135.555 170.290 ;
        RECT 137.155 170.245 137.445 170.290 ;
        RECT 140.275 170.245 140.565 170.290 ;
        RECT 135.775 170.090 136.065 170.135 ;
        RECT 110.920 169.950 122.650 170.090 ;
        RECT 110.920 169.890 111.240 169.950 ;
        RECT 104.940 169.795 105.260 169.810 ;
        RECT 103.575 169.750 103.865 169.795 ;
        RECT 102.180 169.610 103.865 169.750 ;
        RECT 102.180 169.550 102.500 169.610 ;
        RECT 103.575 169.565 103.865 169.610 ;
        RECT 104.035 169.565 104.325 169.795 ;
        RECT 104.895 169.565 105.260 169.795 ;
        RECT 104.940 169.550 105.260 169.565 ;
        RECT 105.400 169.750 105.720 169.810 ;
        RECT 106.795 169.750 107.085 169.795 ;
        RECT 105.400 169.610 107.085 169.750 ;
        RECT 105.400 169.550 105.720 169.610 ;
        RECT 106.795 169.565 107.085 169.610 ;
        RECT 107.240 169.750 107.560 169.810 ;
        RECT 109.095 169.750 109.385 169.795 ;
        RECT 107.240 169.610 109.385 169.750 ;
        RECT 107.240 169.550 107.560 169.610 ;
        RECT 109.095 169.565 109.385 169.610 ;
        RECT 111.380 169.550 111.700 169.810 ;
        RECT 122.510 169.795 122.650 169.950 ;
        RECT 124.735 169.950 134.150 170.090 ;
        RECT 134.930 169.950 136.065 170.090 ;
        RECT 124.735 169.905 125.025 169.950 ;
        RECT 134.010 169.810 134.150 169.950 ;
        RECT 135.775 169.905 136.065 169.950 ;
        RECT 113.235 169.565 113.525 169.795 ;
        RECT 115.995 169.565 116.285 169.795 ;
        RECT 122.435 169.565 122.725 169.795 ;
        RECT 124.260 169.750 124.580 169.810 ;
        RECT 126.575 169.750 126.865 169.795 ;
        RECT 129.840 169.750 130.130 169.795 ;
        RECT 124.260 169.610 126.865 169.750 ;
        RECT 105.030 169.410 105.170 169.550 ;
        RECT 113.310 169.410 113.450 169.565 ;
        RECT 97.670 169.270 101.490 169.410 ;
        RECT 105.030 169.270 113.450 169.410 ;
        RECT 116.070 169.410 116.210 169.565 ;
        RECT 124.260 169.550 124.580 169.610 ;
        RECT 126.575 169.565 126.865 169.610 ;
        RECT 127.595 169.610 130.130 169.750 ;
        RECT 116.440 169.410 116.760 169.470 ;
        RECT 116.070 169.270 116.760 169.410 ;
        RECT 96.660 169.210 96.980 169.270 ;
        RECT 97.135 169.225 97.425 169.270 ;
        RECT 101.350 169.115 101.490 169.270 ;
        RECT 116.440 169.210 116.760 169.270 ;
        RECT 121.055 169.410 121.345 169.455 ;
        RECT 121.500 169.410 121.820 169.470 ;
        RECT 127.595 169.455 127.810 169.610 ;
        RECT 129.840 169.565 130.130 169.610 ;
        RECT 133.920 169.750 134.240 169.810 ;
        RECT 134.395 169.750 134.685 169.795 ;
        RECT 133.920 169.610 134.685 169.750 ;
        RECT 133.920 169.550 134.240 169.610 ;
        RECT 134.395 169.565 134.685 169.610 ;
        RECT 134.860 169.750 135.150 169.795 ;
        RECT 136.695 169.750 136.985 169.795 ;
        RECT 140.275 169.750 140.565 169.795 ;
        RECT 134.860 169.610 140.565 169.750 ;
        RECT 134.860 169.565 135.150 169.610 ;
        RECT 136.695 169.565 136.985 169.610 ;
        RECT 140.275 169.565 140.565 169.610 ;
        RECT 131.620 169.455 131.940 169.470 ;
        RECT 141.355 169.455 141.645 169.770 ;
        RECT 121.055 169.270 121.820 169.410 ;
        RECT 121.055 169.225 121.345 169.270 ;
        RECT 121.500 169.210 121.820 169.270 ;
        RECT 125.660 169.410 125.950 169.455 ;
        RECT 127.520 169.410 127.810 169.455 ;
        RECT 125.660 169.270 127.810 169.410 ;
        RECT 125.660 169.225 125.950 169.270 ;
        RECT 127.520 169.225 127.810 169.270 ;
        RECT 128.440 169.410 128.730 169.455 ;
        RECT 131.620 169.410 131.990 169.455 ;
        RECT 138.055 169.410 138.705 169.455 ;
        RECT 141.355 169.410 141.945 169.455 ;
        RECT 128.440 169.270 141.945 169.410 ;
        RECT 128.440 169.225 128.730 169.270 ;
        RECT 131.620 169.225 131.990 169.270 ;
        RECT 131.620 169.210 131.940 169.225 ;
        RECT 137.690 169.130 137.830 169.270 ;
        RECT 138.055 169.225 138.705 169.270 ;
        RECT 141.655 169.225 141.945 169.270 ;
        RECT 100.815 169.070 101.105 169.115 ;
        RECT 94.910 168.930 101.105 169.070 ;
        RECT 87.015 168.885 87.305 168.930 ;
        RECT 92.060 168.870 92.380 168.930 ;
        RECT 100.815 168.885 101.105 168.930 ;
        RECT 101.275 168.885 101.565 169.115 ;
        RECT 104.480 169.070 104.800 169.130 ;
        RECT 116.900 169.070 117.220 169.130 ;
        RECT 123.800 169.070 124.120 169.130 ;
        RECT 104.480 168.930 124.120 169.070 ;
        RECT 104.480 168.870 104.800 168.930 ;
        RECT 116.900 168.870 117.220 168.930 ;
        RECT 123.800 168.870 124.120 168.930 ;
        RECT 137.600 168.870 137.920 169.130 ;
        RECT 143.120 168.870 143.440 169.130 ;
        RECT 2.750 168.250 159.030 168.730 ;
        RECT 5.580 168.050 5.900 168.110 ;
        RECT 6.055 168.050 6.345 168.095 ;
        RECT 5.580 167.910 6.345 168.050 ;
        RECT 5.580 167.850 5.900 167.910 ;
        RECT 6.055 167.865 6.345 167.910 ;
        RECT 14.320 168.050 14.640 168.110 ;
        RECT 16.175 168.050 16.465 168.095 ;
        RECT 22.140 168.050 22.460 168.110 ;
        RECT 14.320 167.910 16.465 168.050 ;
        RECT 14.320 167.850 14.640 167.910 ;
        RECT 16.175 167.865 16.465 167.910 ;
        RECT 18.090 167.910 22.460 168.050 ;
        RECT 18.090 167.755 18.230 167.910 ;
        RECT 22.140 167.850 22.460 167.910 ;
        RECT 23.060 168.050 23.380 168.110 ;
        RECT 23.060 167.910 23.750 168.050 ;
        RECT 23.060 167.850 23.380 167.910 ;
        RECT 18.015 167.525 18.305 167.755 ;
        RECT 6.975 167.370 7.265 167.415 ;
        RECT 6.975 167.230 8.570 167.370 ;
        RECT 6.975 167.185 7.265 167.230 ;
        RECT 8.430 166.735 8.570 167.230 ;
        RECT 10.180 167.170 10.500 167.430 ;
        RECT 10.655 167.370 10.945 167.415 ;
        RECT 12.495 167.370 12.785 167.415 ;
        RECT 10.655 167.230 12.785 167.370 ;
        RECT 10.655 167.185 10.945 167.230 ;
        RECT 12.495 167.185 12.785 167.230 ;
        RECT 12.940 167.170 13.260 167.430 ;
        RECT 23.610 167.370 23.750 167.910 ;
        RECT 25.450 167.910 26.970 168.050 ;
        RECT 25.450 167.755 25.590 167.910 ;
        RECT 26.830 167.770 26.970 167.910 ;
        RECT 40.655 167.910 47.210 168.050 ;
        RECT 25.375 167.525 25.665 167.755 ;
        RECT 25.820 167.510 26.140 167.770 ;
        RECT 26.740 167.510 27.060 167.770 ;
        RECT 32.720 167.755 33.040 167.770 ;
        RECT 32.715 167.710 33.365 167.755 ;
        RECT 36.315 167.710 36.605 167.755 ;
        RECT 40.655 167.710 40.795 167.910 ;
        RECT 28.210 167.570 36.605 167.710 ;
        RECT 28.210 167.430 28.350 167.570 ;
        RECT 32.715 167.525 33.365 167.570 ;
        RECT 36.015 167.525 36.605 167.570 ;
        RECT 37.410 167.570 40.795 167.710 ;
        RECT 44.235 167.710 44.525 167.755 ;
        RECT 46.535 167.710 46.825 167.755 ;
        RECT 32.720 167.510 33.040 167.525 ;
        RECT 23.995 167.370 24.285 167.415 ;
        RECT 23.610 167.230 24.285 167.370 ;
        RECT 23.995 167.185 24.285 167.230 ;
        RECT 24.440 167.370 24.760 167.430 ;
        RECT 26.320 167.370 26.610 167.415 ;
        RECT 24.440 167.230 24.955 167.370 ;
        RECT 25.220 167.230 26.610 167.370 ;
        RECT 24.440 167.170 24.760 167.230 ;
        RECT 11.560 166.830 11.880 167.090 ;
        RECT 13.030 167.030 13.170 167.170 ;
        RECT 15.255 167.030 15.545 167.075 ;
        RECT 13.030 166.890 15.545 167.030 ;
        RECT 15.255 166.845 15.545 166.890 ;
        RECT 17.080 167.030 17.400 167.090 ;
        RECT 18.475 167.030 18.765 167.075 ;
        RECT 17.080 166.890 18.765 167.030 ;
        RECT 8.355 166.505 8.645 166.735 ;
        RECT 15.330 166.690 15.470 166.845 ;
        RECT 17.080 166.830 17.400 166.890 ;
        RECT 18.475 166.845 18.765 166.890 ;
        RECT 19.380 166.830 19.700 167.090 ;
        RECT 24.440 166.690 24.760 166.750 ;
        RECT 15.330 166.550 24.760 166.690 ;
        RECT 24.440 166.490 24.760 166.550 ;
        RECT 19.840 166.350 20.160 166.410 ;
        RECT 25.220 166.350 25.360 167.230 ;
        RECT 26.320 167.185 26.610 167.230 ;
        RECT 28.120 167.170 28.440 167.430 ;
        RECT 29.040 167.170 29.360 167.430 ;
        RECT 29.520 167.370 29.810 167.415 ;
        RECT 31.355 167.370 31.645 167.415 ;
        RECT 34.935 167.370 35.225 167.415 ;
        RECT 29.520 167.230 35.225 167.370 ;
        RECT 29.520 167.185 29.810 167.230 ;
        RECT 31.355 167.185 31.645 167.230 ;
        RECT 34.935 167.185 35.225 167.230 ;
        RECT 36.015 167.210 36.305 167.525 ;
        RECT 30.880 167.030 31.200 167.090 ;
        RECT 37.410 167.030 37.550 167.570 ;
        RECT 38.240 167.170 38.560 167.430 ;
        RECT 39.160 167.415 39.480 167.430 ;
        RECT 38.995 167.185 39.480 167.415 ;
        RECT 39.160 167.170 39.480 167.185 ;
        RECT 39.620 167.170 39.940 167.430 ;
        RECT 40.655 167.415 40.795 167.570 ;
        RECT 40.095 167.185 40.385 167.415 ;
        RECT 40.580 167.185 40.870 167.415 ;
        RECT 43.085 167.370 43.375 167.585 ;
        RECT 44.235 167.570 46.825 167.710 ;
        RECT 47.070 167.710 47.210 167.910 ;
        RECT 47.440 167.850 47.760 168.110 ;
        RECT 64.920 168.050 65.240 168.110 ;
        RECT 66.300 168.050 66.620 168.110 ;
        RECT 48.455 167.910 52.730 168.050 ;
        RECT 48.455 167.710 48.595 167.910 ;
        RECT 49.740 167.710 50.060 167.770 ;
        RECT 51.595 167.710 51.885 167.755 ;
        RECT 47.070 167.570 48.595 167.710 ;
        RECT 48.910 167.570 51.885 167.710 ;
        RECT 44.235 167.525 44.525 167.570 ;
        RECT 46.535 167.525 46.825 167.570 ;
        RECT 44.680 167.370 45.000 167.430 ;
        RECT 45.600 167.370 45.920 167.430 ;
        RECT 43.085 167.355 45.920 167.370 ;
        RECT 43.210 167.230 45.920 167.355 ;
        RECT 46.610 167.370 46.750 167.525 ;
        RECT 47.900 167.370 48.220 167.430 ;
        RECT 48.910 167.415 49.050 167.570 ;
        RECT 49.740 167.510 50.060 167.570 ;
        RECT 51.595 167.525 51.885 167.570 ;
        RECT 46.610 167.230 48.220 167.370 ;
        RECT 40.170 167.030 40.310 167.185 ;
        RECT 44.680 167.170 45.000 167.230 ;
        RECT 45.600 167.170 45.920 167.230 ;
        RECT 47.900 167.170 48.220 167.230 ;
        RECT 48.835 167.185 49.125 167.415 ;
        RECT 50.215 167.185 50.505 167.415 ;
        RECT 50.660 167.370 50.980 167.430 ;
        RECT 52.590 167.415 52.730 167.910 ;
        RECT 53.970 167.910 66.620 168.050 ;
        RECT 50.660 167.230 51.175 167.370 ;
        RECT 30.880 166.890 37.550 167.030 ;
        RECT 37.870 166.890 40.310 167.030 ;
        RECT 49.280 167.030 49.600 167.090 ;
        RECT 49.755 167.030 50.045 167.075 ;
        RECT 49.280 166.890 50.045 167.030 ;
        RECT 30.880 166.830 31.200 166.890 ;
        RECT 27.215 166.690 27.505 166.735 ;
        RECT 29.040 166.690 29.360 166.750 ;
        RECT 27.215 166.550 29.360 166.690 ;
        RECT 27.215 166.505 27.505 166.550 ;
        RECT 29.040 166.490 29.360 166.550 ;
        RECT 29.925 166.690 30.215 166.735 ;
        RECT 31.815 166.690 32.105 166.735 ;
        RECT 34.935 166.690 35.225 166.735 ;
        RECT 29.925 166.550 35.225 166.690 ;
        RECT 29.925 166.505 30.215 166.550 ;
        RECT 31.815 166.505 32.105 166.550 ;
        RECT 34.935 166.505 35.225 166.550 ;
        RECT 35.940 166.690 36.260 166.750 ;
        RECT 36.860 166.690 37.180 166.750 ;
        RECT 35.940 166.550 37.180 166.690 ;
        RECT 35.940 166.490 36.260 166.550 ;
        RECT 36.860 166.490 37.180 166.550 ;
        RECT 19.840 166.210 25.360 166.350 ;
        RECT 27.660 166.350 27.980 166.410 ;
        RECT 30.340 166.350 30.630 166.395 ;
        RECT 27.660 166.210 30.630 166.350 ;
        RECT 19.840 166.150 20.160 166.210 ;
        RECT 27.660 166.150 27.980 166.210 ;
        RECT 30.340 166.165 30.630 166.210 ;
        RECT 34.100 166.350 34.420 166.410 ;
        RECT 37.870 166.395 38.010 166.890 ;
        RECT 49.280 166.830 49.600 166.890 ;
        RECT 49.755 166.845 50.045 166.890 ;
        RECT 42.395 166.690 42.685 166.735 ;
        RECT 42.840 166.690 43.160 166.750 ;
        RECT 42.395 166.550 43.160 166.690 ;
        RECT 42.395 166.505 42.685 166.550 ;
        RECT 42.840 166.490 43.160 166.550 ;
        RECT 44.680 166.490 45.000 166.750 ;
        RECT 46.060 166.690 46.380 166.750 ;
        RECT 47.915 166.690 48.205 166.735 ;
        RECT 46.060 166.550 48.205 166.690 ;
        RECT 46.060 166.490 46.380 166.550 ;
        RECT 47.915 166.505 48.205 166.550 ;
        RECT 48.360 166.690 48.680 166.750 ;
        RECT 50.290 166.690 50.430 167.185 ;
        RECT 50.660 167.170 50.980 167.230 ;
        RECT 52.055 167.185 52.345 167.415 ;
        RECT 52.540 167.370 52.830 167.415 ;
        RECT 53.420 167.370 53.740 167.430 ;
        RECT 52.540 167.230 53.740 167.370 ;
        RECT 52.540 167.185 52.830 167.230 ;
        RECT 52.130 167.030 52.270 167.185 ;
        RECT 53.420 167.170 53.740 167.230 ;
        RECT 53.970 167.030 54.110 167.910 ;
        RECT 64.920 167.850 65.240 167.910 ;
        RECT 66.300 167.850 66.620 167.910 ;
        RECT 68.615 167.865 68.905 168.095 ;
        RECT 54.815 167.710 55.105 167.755 ;
        RECT 55.260 167.710 55.580 167.770 ;
        RECT 54.815 167.570 55.580 167.710 ;
        RECT 54.815 167.525 55.105 167.570 ;
        RECT 55.260 167.510 55.580 167.570 ;
        RECT 56.180 167.510 56.500 167.770 ;
        RECT 56.640 167.510 56.960 167.770 ;
        RECT 59.400 167.710 59.720 167.770 ;
        RECT 60.780 167.710 61.100 167.770 ;
        RECT 57.235 167.570 61.100 167.710 ;
        RECT 57.235 167.430 57.375 167.570 ;
        RECT 59.400 167.510 59.720 167.570 ;
        RECT 60.780 167.510 61.100 167.570 ;
        RECT 61.255 167.710 61.545 167.755 ;
        RECT 62.620 167.710 62.940 167.770 ;
        RECT 63.540 167.755 63.860 167.770 ;
        RECT 61.255 167.570 62.940 167.710 ;
        RECT 61.255 167.525 61.545 167.570 ;
        RECT 62.620 167.510 62.940 167.570 ;
        RECT 63.535 167.710 64.185 167.755 ;
        RECT 67.135 167.710 67.425 167.755 ;
        RECT 63.535 167.570 67.425 167.710 ;
        RECT 63.535 167.525 64.185 167.570 ;
        RECT 66.835 167.525 67.425 167.570 ;
        RECT 68.690 167.710 68.830 167.865 ;
        RECT 69.520 167.850 69.840 168.110 ;
        RECT 77.340 168.050 77.660 168.110 ;
        RECT 70.070 167.910 77.660 168.050 ;
        RECT 70.070 167.710 70.210 167.910 ;
        RECT 77.340 167.850 77.660 167.910 ;
        RECT 77.800 168.050 78.120 168.110 ;
        RECT 88.840 168.050 89.160 168.110 ;
        RECT 92.520 168.050 92.840 168.110 ;
        RECT 98.515 168.050 98.805 168.095 ;
        RECT 77.800 167.910 88.610 168.050 ;
        RECT 77.800 167.850 78.120 167.910 ;
        RECT 70.440 167.755 70.760 167.770 ;
        RECT 68.690 167.570 70.210 167.710 ;
        RECT 63.540 167.510 63.860 167.525 ;
        RECT 55.735 167.360 56.025 167.415 ;
        RECT 57.100 167.370 57.420 167.430 ;
        RECT 56.270 167.360 57.420 167.370 ;
        RECT 55.735 167.230 57.420 167.360 ;
        RECT 55.735 167.220 56.410 167.230 ;
        RECT 55.735 167.185 56.025 167.220 ;
        RECT 57.100 167.170 57.420 167.230 ;
        RECT 57.560 167.170 57.880 167.430 ;
        RECT 58.480 167.170 58.800 167.430 ;
        RECT 60.340 167.370 60.630 167.415 ;
        RECT 62.175 167.370 62.465 167.415 ;
        RECT 65.755 167.370 66.045 167.415 ;
        RECT 60.340 167.230 66.045 167.370 ;
        RECT 60.340 167.185 60.630 167.230 ;
        RECT 62.175 167.185 62.465 167.230 ;
        RECT 65.755 167.185 66.045 167.230 ;
        RECT 66.835 167.210 67.125 167.525 ;
        RECT 52.130 166.890 54.110 167.030 ;
        RECT 54.800 167.030 55.120 167.090 ;
        RECT 56.640 167.030 56.960 167.090 ;
        RECT 54.800 166.890 56.960 167.030 ;
        RECT 54.800 166.830 55.120 166.890 ;
        RECT 56.640 166.830 56.960 166.890 ;
        RECT 59.860 166.830 60.180 167.090 ;
        RECT 61.240 167.030 61.560 167.090 ;
        RECT 68.690 167.030 68.830 167.570 ;
        RECT 70.375 167.525 70.760 167.755 ;
        RECT 70.440 167.510 70.760 167.525 ;
        RECT 71.360 167.510 71.680 167.770 ;
        RECT 73.215 167.185 73.505 167.415 ;
        RECT 73.675 167.370 73.965 167.415 ;
        RECT 74.120 167.370 74.440 167.430 ;
        RECT 73.675 167.230 74.440 167.370 ;
        RECT 73.675 167.185 73.965 167.230 ;
        RECT 61.240 166.890 68.830 167.030 ;
        RECT 61.240 166.830 61.560 166.890 ;
        RECT 72.280 166.830 72.600 167.090 ;
        RECT 48.360 166.550 50.430 166.690 ;
        RECT 52.960 166.690 53.280 166.750 ;
        RECT 53.435 166.690 53.725 166.735 ;
        RECT 52.960 166.550 53.725 166.690 ;
        RECT 48.360 166.490 48.680 166.550 ;
        RECT 52.960 166.490 53.280 166.550 ;
        RECT 53.435 166.505 53.725 166.550 ;
        RECT 58.020 166.690 58.340 166.750 ;
        RECT 59.950 166.690 60.090 166.830 ;
        RECT 73.290 166.750 73.430 167.185 ;
        RECT 74.120 167.170 74.440 167.230 ;
        RECT 77.800 167.170 78.120 167.430 ;
        RECT 81.570 167.415 81.710 167.910 ;
        RECT 88.470 167.770 88.610 167.910 ;
        RECT 88.840 167.910 92.290 168.050 ;
        RECT 88.840 167.850 89.160 167.910 ;
        RECT 82.860 167.710 83.180 167.770 ;
        RECT 86.555 167.710 86.845 167.755 ;
        RECT 82.860 167.570 84.010 167.710 ;
        RECT 82.860 167.510 83.180 167.570 ;
        RECT 81.495 167.185 81.785 167.415 ;
        RECT 81.940 167.370 82.260 167.430 ;
        RECT 82.415 167.370 82.705 167.415 ;
        RECT 81.940 167.230 82.705 167.370 ;
        RECT 81.940 167.170 82.260 167.230 ;
        RECT 82.415 167.185 82.705 167.230 ;
        RECT 83.335 167.185 83.625 167.415 ;
        RECT 74.580 167.030 74.900 167.090 ;
        RECT 77.355 167.030 77.645 167.075 ;
        RECT 74.580 166.890 77.645 167.030 ;
        RECT 77.890 167.030 78.030 167.170 ;
        RECT 82.030 167.030 82.170 167.170 ;
        RECT 77.890 166.890 82.170 167.030 ;
        RECT 74.580 166.830 74.900 166.890 ;
        RECT 58.020 166.550 60.090 166.690 ;
        RECT 58.020 166.490 58.340 166.550 ;
        RECT 37.795 166.350 38.085 166.395 ;
        RECT 34.100 166.210 38.085 166.350 ;
        RECT 34.100 166.150 34.420 166.210 ;
        RECT 37.795 166.165 38.085 166.210 ;
        RECT 39.160 166.350 39.480 166.410 ;
        RECT 41.475 166.350 41.765 166.395 ;
        RECT 39.160 166.210 41.765 166.350 ;
        RECT 39.160 166.150 39.480 166.210 ;
        RECT 41.475 166.165 41.765 166.210 ;
        RECT 43.315 166.350 43.605 166.395 ;
        RECT 44.770 166.350 44.910 166.490 ;
        RECT 43.315 166.210 44.910 166.350 ;
        RECT 45.600 166.350 45.920 166.410 ;
        RECT 46.535 166.350 46.825 166.395 ;
        RECT 53.880 166.350 54.200 166.410 ;
        RECT 45.600 166.210 54.200 166.350 ;
        RECT 43.315 166.165 43.605 166.210 ;
        RECT 45.600 166.150 45.920 166.210 ;
        RECT 46.535 166.165 46.825 166.210 ;
        RECT 53.880 166.150 54.200 166.210 ;
        RECT 59.400 166.150 59.720 166.410 ;
        RECT 59.950 166.350 60.090 166.550 ;
        RECT 60.745 166.690 61.035 166.735 ;
        RECT 62.635 166.690 62.925 166.735 ;
        RECT 65.755 166.690 66.045 166.735 ;
        RECT 60.745 166.550 66.045 166.690 ;
        RECT 60.745 166.505 61.035 166.550 ;
        RECT 62.635 166.505 62.925 166.550 ;
        RECT 65.755 166.505 66.045 166.550 ;
        RECT 66.300 166.690 66.620 166.750 ;
        RECT 73.200 166.690 73.520 166.750 ;
        RECT 66.300 166.550 73.520 166.690 ;
        RECT 66.300 166.490 66.620 166.550 ;
        RECT 73.200 166.490 73.520 166.550 ;
        RECT 75.040 166.690 75.360 166.750 ;
        RECT 75.515 166.690 75.805 166.735 ;
        RECT 75.040 166.550 75.805 166.690 ;
        RECT 75.040 166.490 75.360 166.550 ;
        RECT 75.515 166.505 75.805 166.550 ;
        RECT 75.960 166.490 76.280 166.750 ;
        RECT 76.970 166.690 77.110 166.890 ;
        RECT 77.355 166.845 77.645 166.890 ;
        RECT 82.860 166.830 83.180 167.090 ;
        RECT 76.970 166.550 79.870 166.690 ;
        RECT 67.680 166.350 68.000 166.410 ;
        RECT 59.950 166.210 68.000 166.350 ;
        RECT 67.680 166.150 68.000 166.210 ;
        RECT 70.455 166.350 70.745 166.395 ;
        RECT 79.180 166.350 79.500 166.410 ;
        RECT 70.455 166.210 79.500 166.350 ;
        RECT 79.730 166.350 79.870 166.550 ;
        RECT 80.560 166.490 80.880 166.750 ;
        RECT 83.410 166.690 83.550 167.185 ;
        RECT 83.870 167.030 84.010 167.570 ;
        RECT 84.330 167.570 86.845 167.710 ;
        RECT 84.330 167.415 84.470 167.570 ;
        RECT 86.555 167.525 86.845 167.570 ;
        RECT 88.380 167.710 88.700 167.770 ;
        RECT 92.150 167.710 92.290 167.910 ;
        RECT 92.520 167.910 98.805 168.050 ;
        RECT 92.520 167.850 92.840 167.910 ;
        RECT 98.515 167.865 98.805 167.910 ;
        RECT 101.735 168.050 102.025 168.095 ;
        RECT 102.640 168.050 102.960 168.110 ;
        RECT 101.735 167.910 102.960 168.050 ;
        RECT 101.735 167.865 102.025 167.910 ;
        RECT 102.640 167.850 102.960 167.910 ;
        RECT 104.020 168.050 104.340 168.110 ;
        RECT 107.240 168.050 107.560 168.110 ;
        RECT 104.020 167.910 107.560 168.050 ;
        RECT 104.020 167.850 104.340 167.910 ;
        RECT 107.240 167.850 107.560 167.910 ;
        RECT 148.640 167.850 148.960 168.110 ;
        RECT 98.960 167.710 99.280 167.770 ;
        RECT 88.380 167.570 89.530 167.710 ;
        RECT 92.150 167.570 99.280 167.710 ;
        RECT 88.380 167.510 88.700 167.570 ;
        RECT 84.255 167.185 84.545 167.415 ;
        RECT 84.700 167.170 85.020 167.430 ;
        RECT 85.635 167.185 85.925 167.415 ;
        RECT 85.710 167.030 85.850 167.185 ;
        RECT 88.840 167.170 89.160 167.430 ;
        RECT 89.390 167.415 89.530 167.570 ;
        RECT 98.960 167.510 99.280 167.570 ;
        RECT 99.435 167.710 99.725 167.755 ;
        RECT 104.480 167.710 104.800 167.770 ;
        RECT 99.435 167.570 104.800 167.710 ;
        RECT 99.435 167.525 99.725 167.570 ;
        RECT 104.480 167.510 104.800 167.570 ;
        RECT 106.780 167.710 107.100 167.770 ;
        RECT 123.340 167.755 123.660 167.770 ;
        RECT 119.775 167.710 120.065 167.755 ;
        RECT 123.015 167.710 123.665 167.755 ;
        RECT 131.620 167.710 131.940 167.770 ;
        RECT 106.780 167.570 110.230 167.710 ;
        RECT 106.780 167.510 107.100 167.570 ;
        RECT 89.315 167.185 89.605 167.415 ;
        RECT 89.775 167.370 90.065 167.415 ;
        RECT 91.140 167.370 91.460 167.430 ;
        RECT 92.535 167.370 92.825 167.415 ;
        RECT 89.775 167.230 91.460 167.370 ;
        RECT 89.775 167.185 90.065 167.230 ;
        RECT 91.140 167.170 91.460 167.230 ;
        RECT 91.690 167.230 92.825 167.370 ;
        RECT 86.080 167.030 86.400 167.090 ;
        RECT 83.870 166.890 86.400 167.030 ;
        RECT 86.080 166.830 86.400 166.890 ;
        RECT 88.395 166.845 88.685 167.075 ;
        RECT 90.220 167.030 90.540 167.090 ;
        RECT 91.690 167.030 91.830 167.230 ;
        RECT 92.535 167.185 92.825 167.230 ;
        RECT 92.980 167.170 93.300 167.430 ;
        RECT 94.820 167.170 95.140 167.430 ;
        RECT 100.355 167.370 100.645 167.415 ;
        RECT 101.720 167.370 102.040 167.430 ;
        RECT 96.520 167.230 102.040 167.370 ;
        RECT 90.220 166.890 91.830 167.030 ;
        RECT 85.620 166.690 85.940 166.750 ;
        RECT 83.410 166.550 85.940 166.690 ;
        RECT 88.470 166.690 88.610 166.845 ;
        RECT 90.220 166.830 90.540 166.890 ;
        RECT 92.060 166.830 92.380 167.090 ;
        RECT 93.440 166.830 93.760 167.090 ;
        RECT 96.520 167.030 96.660 167.230 ;
        RECT 100.355 167.185 100.645 167.230 ;
        RECT 101.720 167.170 102.040 167.230 ;
        RECT 103.100 167.170 103.420 167.430 ;
        RECT 107.330 167.415 107.470 167.570 ;
        RECT 105.415 167.400 105.705 167.415 ;
        RECT 105.030 167.370 105.705 167.400 ;
        RECT 103.650 167.260 105.705 167.370 ;
        RECT 103.650 167.230 105.170 167.260 ;
        RECT 93.990 166.890 96.660 167.030 ;
        RECT 98.055 167.030 98.345 167.075 ;
        RECT 98.500 167.030 98.820 167.090 ;
        RECT 98.055 166.890 98.820 167.030 ;
        RECT 91.155 166.690 91.445 166.735 ;
        RECT 88.470 166.550 91.445 166.690 ;
        RECT 85.620 166.490 85.940 166.550 ;
        RECT 91.155 166.505 91.445 166.550 ;
        RECT 91.600 166.690 91.920 166.750 ;
        RECT 93.990 166.690 94.130 166.890 ;
        RECT 98.055 166.845 98.345 166.890 ;
        RECT 98.500 166.830 98.820 166.890 ;
        RECT 102.640 167.030 102.960 167.090 ;
        RECT 103.650 167.030 103.790 167.230 ;
        RECT 105.415 167.185 105.705 167.260 ;
        RECT 107.255 167.185 107.545 167.415 ;
        RECT 107.715 167.370 108.005 167.415 ;
        RECT 109.540 167.370 109.860 167.430 ;
        RECT 107.715 167.230 109.860 167.370 ;
        RECT 110.090 167.370 110.230 167.570 ;
        RECT 119.775 167.570 131.940 167.710 ;
        RECT 119.775 167.525 120.365 167.570 ;
        RECT 123.015 167.525 123.665 167.570 ;
        RECT 110.090 167.230 117.130 167.370 ;
        RECT 107.715 167.185 108.005 167.230 ;
        RECT 109.540 167.170 109.860 167.230 ;
        RECT 102.640 166.890 103.790 167.030 ;
        RECT 104.035 167.030 104.325 167.075 ;
        RECT 110.460 167.030 110.780 167.090 ;
        RECT 104.035 166.890 110.780 167.030 ;
        RECT 102.640 166.830 102.960 166.890 ;
        RECT 104.035 166.845 104.325 166.890 ;
        RECT 110.320 166.830 110.780 166.890 ;
        RECT 115.060 167.030 115.380 167.090 ;
        RECT 116.990 167.075 117.130 167.230 ;
        RECT 120.075 167.210 120.365 167.525 ;
        RECT 123.340 167.510 123.660 167.525 ;
        RECT 131.620 167.510 131.940 167.570 ;
        RECT 133.000 167.510 133.320 167.770 ;
        RECT 148.730 167.710 148.870 167.850 ;
        RECT 135.390 167.570 142.430 167.710 ;
        RECT 148.730 167.570 150.250 167.710 ;
        RECT 135.390 167.430 135.530 167.570 ;
        RECT 121.155 167.370 121.445 167.415 ;
        RECT 124.735 167.370 125.025 167.415 ;
        RECT 126.570 167.370 126.860 167.415 ;
        RECT 121.155 167.230 126.860 167.370 ;
        RECT 121.155 167.185 121.445 167.230 ;
        RECT 124.735 167.185 125.025 167.230 ;
        RECT 126.570 167.185 126.860 167.230 ;
        RECT 133.935 167.185 134.225 167.415 ;
        RECT 134.380 167.370 134.700 167.430 ;
        RECT 134.380 167.230 135.070 167.370 ;
        RECT 115.535 167.030 115.825 167.075 ;
        RECT 115.060 166.890 115.825 167.030 ;
        RECT 115.060 166.830 115.380 166.890 ;
        RECT 115.535 166.845 115.825 166.890 ;
        RECT 116.915 166.845 117.205 167.075 ;
        RECT 120.580 166.830 120.900 167.090 ;
        RECT 127.035 166.845 127.325 167.075 ;
        RECT 133.000 167.030 133.320 167.090 ;
        RECT 134.010 167.030 134.150 167.185 ;
        RECT 134.380 167.170 134.700 167.230 ;
        RECT 134.930 167.030 135.070 167.230 ;
        RECT 135.300 167.170 135.620 167.430 ;
        RECT 142.290 167.415 142.430 167.570 ;
        RECT 137.155 167.185 137.445 167.415 ;
        RECT 142.215 167.370 142.505 167.415 ;
        RECT 143.120 167.370 143.440 167.430 ;
        RECT 144.515 167.370 144.805 167.415 ;
        RECT 142.215 167.230 144.805 167.370 ;
        RECT 142.215 167.185 142.505 167.230 ;
        RECT 137.230 167.030 137.370 167.185 ;
        RECT 143.120 167.170 143.440 167.230 ;
        RECT 144.515 167.185 144.805 167.230 ;
        RECT 149.560 167.170 149.880 167.430 ;
        RECT 150.110 167.415 150.250 167.570 ;
        RECT 150.035 167.185 150.325 167.415 ;
        RECT 133.000 166.890 134.610 167.030 ;
        RECT 134.930 166.890 137.370 167.030 ;
        RECT 104.495 166.690 104.785 166.735 ;
        RECT 108.620 166.690 108.940 166.750 ;
        RECT 110.320 166.690 110.460 166.830 ;
        RECT 120.670 166.690 120.810 166.830 ;
        RECT 91.600 166.550 94.130 166.690 ;
        RECT 96.750 166.550 104.250 166.690 ;
        RECT 91.600 166.490 91.920 166.550 ;
        RECT 96.750 166.410 96.890 166.550 ;
        RECT 90.220 166.350 90.540 166.410 ;
        RECT 79.730 166.210 90.540 166.350 ;
        RECT 70.455 166.165 70.745 166.210 ;
        RECT 79.180 166.150 79.500 166.210 ;
        RECT 90.220 166.150 90.540 166.210 ;
        RECT 90.695 166.350 90.985 166.395 ;
        RECT 95.740 166.350 96.060 166.410 ;
        RECT 90.695 166.210 96.060 166.350 ;
        RECT 90.695 166.165 90.985 166.210 ;
        RECT 95.740 166.150 96.060 166.210 ;
        RECT 96.660 166.150 96.980 166.410 ;
        RECT 102.180 166.350 102.500 166.410 ;
        RECT 103.560 166.350 103.880 166.410 ;
        RECT 102.180 166.210 103.880 166.350 ;
        RECT 104.110 166.350 104.250 166.550 ;
        RECT 104.495 166.550 109.770 166.690 ;
        RECT 110.320 166.550 120.810 166.690 ;
        RECT 121.155 166.690 121.445 166.735 ;
        RECT 124.275 166.690 124.565 166.735 ;
        RECT 126.165 166.690 126.455 166.735 ;
        RECT 121.155 166.550 126.455 166.690 ;
        RECT 127.110 166.690 127.250 166.845 ;
        RECT 133.000 166.830 133.320 166.890 ;
        RECT 133.920 166.690 134.240 166.750 ;
        RECT 127.110 166.550 134.240 166.690 ;
        RECT 134.470 166.690 134.610 166.890 ;
        RECT 138.075 166.845 138.365 167.075 ;
        RECT 138.150 166.690 138.290 166.845 ;
        RECT 140.820 166.830 141.140 167.090 ;
        RECT 134.470 166.550 138.290 166.690 ;
        RECT 104.495 166.505 104.785 166.550 ;
        RECT 108.620 166.490 108.940 166.550 ;
        RECT 106.795 166.350 107.085 166.395 ;
        RECT 104.110 166.210 107.085 166.350 ;
        RECT 109.630 166.350 109.770 166.550 ;
        RECT 121.155 166.505 121.445 166.550 ;
        RECT 124.275 166.505 124.565 166.550 ;
        RECT 126.165 166.505 126.455 166.550 ;
        RECT 133.920 166.490 134.240 166.550 ;
        RECT 110.920 166.350 111.240 166.410 ;
        RECT 109.630 166.210 111.240 166.350 ;
        RECT 102.180 166.150 102.500 166.210 ;
        RECT 103.560 166.150 103.880 166.210 ;
        RECT 106.795 166.165 107.085 166.210 ;
        RECT 110.920 166.150 111.240 166.210 ;
        RECT 114.600 166.350 114.920 166.410 ;
        RECT 123.340 166.350 123.660 166.410 ;
        RECT 114.600 166.210 123.660 166.350 ;
        RECT 114.600 166.150 114.920 166.210 ;
        RECT 123.340 166.150 123.660 166.210 ;
        RECT 124.720 166.350 125.040 166.410 ;
        RECT 125.715 166.350 126.005 166.395 ;
        RECT 124.720 166.210 126.005 166.350 ;
        RECT 124.720 166.150 125.040 166.210 ;
        RECT 125.715 166.165 126.005 166.210 ;
        RECT 147.720 166.150 148.040 166.410 ;
        RECT 150.940 166.150 151.260 166.410 ;
        RECT 2.750 165.530 158.230 166.010 ;
        RECT 12.940 165.375 13.260 165.390 ;
        RECT 12.940 165.330 13.475 165.375 ;
        RECT 20.300 165.330 20.620 165.390 ;
        RECT 24.440 165.330 24.760 165.390 ;
        RECT 12.940 165.190 19.610 165.330 ;
        RECT 12.940 165.145 13.475 165.190 ;
        RECT 12.940 165.130 13.260 165.145 ;
        RECT 4.680 164.990 4.970 165.035 ;
        RECT 6.540 164.990 6.830 165.035 ;
        RECT 9.320 164.990 9.610 165.035 ;
        RECT 4.680 164.850 9.610 164.990 ;
        RECT 4.680 164.805 4.970 164.850 ;
        RECT 6.540 164.805 6.830 164.850 ;
        RECT 9.320 164.805 9.610 164.850 ;
        RECT 10.640 164.990 10.960 165.050 ;
        RECT 17.540 164.990 17.860 165.050 ;
        RECT 10.640 164.850 17.860 164.990 ;
        RECT 10.640 164.790 10.960 164.850 ;
        RECT 17.540 164.790 17.860 164.850 ;
        RECT 4.200 164.650 4.520 164.710 ;
        RECT 10.730 164.650 10.870 164.790 ;
        RECT 4.200 164.510 10.870 164.650 ;
        RECT 11.560 164.650 11.880 164.710 ;
        RECT 18.935 164.650 19.225 164.695 ;
        RECT 11.560 164.510 19.225 164.650 ;
        RECT 19.470 164.650 19.610 165.190 ;
        RECT 20.300 165.190 24.760 165.330 ;
        RECT 20.300 165.130 20.620 165.190 ;
        RECT 24.440 165.130 24.760 165.190 ;
        RECT 27.660 165.130 27.980 165.390 ;
        RECT 29.500 165.330 29.820 165.390 ;
        RECT 34.575 165.330 34.865 165.375 ;
        RECT 37.320 165.330 37.640 165.390 ;
        RECT 50.200 165.330 50.520 165.390 ;
        RECT 29.500 165.190 37.640 165.330 ;
        RECT 29.500 165.130 29.820 165.190 ;
        RECT 34.575 165.145 34.865 165.190 ;
        RECT 37.320 165.130 37.640 165.190 ;
        RECT 37.870 165.190 50.520 165.330 ;
        RECT 37.870 164.990 38.010 165.190 ;
        RECT 50.200 165.130 50.520 165.190 ;
        RECT 50.660 165.330 50.980 165.390 ;
        RECT 50.660 165.190 61.930 165.330 ;
        RECT 50.660 165.130 50.980 165.190 ;
        RECT 31.430 164.850 38.010 164.990 ;
        RECT 38.700 164.990 39.020 165.050 ;
        RECT 46.995 164.990 47.285 165.035 ;
        RECT 38.700 164.850 47.285 164.990 ;
        RECT 31.430 164.710 31.570 164.850 ;
        RECT 38.700 164.790 39.020 164.850 ;
        RECT 46.995 164.805 47.285 164.850 ;
        RECT 48.820 164.990 49.140 165.050 ;
        RECT 53.845 164.990 54.135 165.035 ;
        RECT 55.735 164.990 56.025 165.035 ;
        RECT 58.855 164.990 59.145 165.035 ;
        RECT 48.820 164.850 51.810 164.990 ;
        RECT 48.820 164.790 49.140 164.850 ;
        RECT 30.880 164.650 31.200 164.710 ;
        RECT 19.470 164.510 22.835 164.650 ;
        RECT 4.200 164.450 4.520 164.510 ;
        RECT 11.560 164.450 11.880 164.510 ;
        RECT 18.935 164.465 19.225 164.510 ;
        RECT 6.055 164.310 6.345 164.355 ;
        RECT 9.320 164.310 9.610 164.355 ;
        RECT 2.910 164.170 6.345 164.310 ;
        RECT 2.910 163.970 3.050 164.170 ;
        RECT 6.055 164.125 6.345 164.170 ;
        RECT 7.075 164.170 9.610 164.310 ;
        RECT 7.075 164.015 7.290 164.170 ;
        RECT 9.320 164.125 9.610 164.170 ;
        RECT 14.795 164.310 15.085 164.355 ;
        RECT 19.010 164.310 19.150 164.465 ;
        RECT 20.300 164.310 20.620 164.370 ;
        RECT 14.795 164.170 16.390 164.310 ;
        RECT 19.010 164.170 20.620 164.310 ;
        RECT 14.795 164.125 15.085 164.170 ;
        RECT 2.450 163.830 3.050 163.970 ;
        RECT 5.140 163.970 5.430 164.015 ;
        RECT 7.000 163.970 7.290 164.015 ;
        RECT 5.140 163.830 7.290 163.970 ;
        RECT 2.450 162.610 2.590 163.830 ;
        RECT 5.140 163.785 5.430 163.830 ;
        RECT 7.000 163.785 7.290 163.830 ;
        RECT 7.920 163.970 8.210 164.015 ;
        RECT 8.800 163.970 9.120 164.030 ;
        RECT 11.180 163.970 11.470 164.015 ;
        RECT 7.920 163.830 11.470 163.970 ;
        RECT 7.920 163.785 8.210 163.830 ;
        RECT 8.800 163.770 9.120 163.830 ;
        RECT 11.180 163.785 11.470 163.830 ;
        RECT 13.860 163.430 14.180 163.690 ;
        RECT 16.250 163.675 16.390 164.170 ;
        RECT 20.300 164.110 20.620 164.170 ;
        RECT 20.760 164.310 21.080 164.370 ;
        RECT 22.695 164.355 22.835 164.510 ;
        RECT 23.150 164.510 31.200 164.650 ;
        RECT 22.155 164.310 22.445 164.355 ;
        RECT 20.760 164.170 22.445 164.310 ;
        RECT 20.760 164.110 21.080 164.170 ;
        RECT 22.155 164.125 22.445 164.170 ;
        RECT 22.620 164.125 22.910 164.355 ;
        RECT 16.620 163.970 16.940 164.030 ;
        RECT 18.015 163.970 18.305 164.015 ;
        RECT 16.620 163.830 18.305 163.970 ;
        RECT 16.620 163.770 16.940 163.830 ;
        RECT 18.015 163.785 18.305 163.830 ;
        RECT 16.175 163.445 16.465 163.675 ;
        RECT 18.460 163.430 18.780 163.690 ;
        RECT 23.150 163.630 23.290 164.510 ;
        RECT 23.980 164.110 24.300 164.370 ;
        RECT 24.555 164.355 24.695 164.510 ;
        RECT 30.880 164.450 31.200 164.510 ;
        RECT 31.340 164.450 31.660 164.710 ;
        RECT 34.560 164.450 34.880 164.710 ;
        RECT 46.520 164.650 46.840 164.710 ;
        RECT 51.670 164.695 51.810 164.850 ;
        RECT 53.845 164.850 59.145 164.990 ;
        RECT 53.845 164.805 54.135 164.850 ;
        RECT 55.735 164.805 56.025 164.850 ;
        RECT 58.855 164.805 59.145 164.850 ;
        RECT 46.520 164.510 51.355 164.650 ;
        RECT 46.520 164.450 46.840 164.510 ;
        RECT 24.480 164.125 24.770 164.355 ;
        RECT 26.755 164.310 27.045 164.355 ;
        RECT 29.975 164.310 30.265 164.355 ;
        RECT 34.100 164.310 34.420 164.370 ;
        RECT 26.755 164.170 28.350 164.310 ;
        RECT 26.755 164.125 27.045 164.170 ;
        RECT 23.535 163.970 23.825 164.015 ;
        RECT 23.535 163.830 26.970 163.970 ;
        RECT 23.535 163.785 23.825 163.830 ;
        RECT 26.830 163.690 26.970 163.830 ;
        RECT 23.980 163.630 24.300 163.690 ;
        RECT 23.150 163.490 24.300 163.630 ;
        RECT 23.980 163.430 24.300 163.490 ;
        RECT 25.360 163.430 25.680 163.690 ;
        RECT 26.740 163.430 27.060 163.690 ;
        RECT 28.210 163.675 28.350 164.170 ;
        RECT 29.975 164.170 34.420 164.310 ;
        RECT 29.975 164.125 30.265 164.170 ;
        RECT 34.100 164.110 34.420 164.170 ;
        RECT 30.435 163.970 30.725 164.015 ;
        RECT 34.650 163.970 34.790 164.450 ;
        RECT 38.240 164.310 38.560 164.370 ;
        RECT 41.935 164.310 42.225 164.355 ;
        RECT 38.240 164.170 42.225 164.310 ;
        RECT 38.240 164.110 38.560 164.170 ;
        RECT 41.935 164.125 42.225 164.170 ;
        RECT 42.400 164.125 42.690 164.355 ;
        RECT 30.435 163.830 34.790 163.970 ;
        RECT 40.080 163.970 40.400 164.030 ;
        RECT 41.015 163.970 41.305 164.015 ;
        RECT 40.080 163.830 41.305 163.970 ;
        RECT 30.435 163.785 30.725 163.830 ;
        RECT 40.080 163.770 40.400 163.830 ;
        RECT 41.015 163.785 41.305 163.830 ;
        RECT 28.135 163.445 28.425 163.675 ;
        RECT 37.780 163.630 38.100 163.690 ;
        RECT 42.470 163.630 42.610 164.125 ;
        RECT 43.760 164.110 44.080 164.370 ;
        RECT 44.680 164.355 45.000 164.370 ;
        RECT 44.465 164.125 45.000 164.355 ;
        RECT 44.680 164.110 45.000 164.125 ;
        RECT 50.660 164.110 50.980 164.370 ;
        RECT 43.315 163.970 43.605 164.015 ;
        RECT 43.315 163.830 43.990 163.970 ;
        RECT 43.315 163.785 43.605 163.830 ;
        RECT 43.850 163.690 43.990 163.830 ;
        RECT 47.900 163.770 48.220 164.030 ;
        RECT 51.215 163.970 51.355 164.510 ;
        RECT 51.595 164.465 51.885 164.695 ;
        RECT 52.500 164.650 52.820 164.710 ;
        RECT 52.975 164.650 53.265 164.695 ;
        RECT 58.020 164.650 58.340 164.710 ;
        RECT 61.790 164.695 61.930 165.190 ;
        RECT 65.840 165.130 66.160 165.390 ;
        RECT 67.680 165.330 68.000 165.390 ;
        RECT 68.600 165.330 68.920 165.390 ;
        RECT 75.055 165.330 75.345 165.375 ;
        RECT 75.500 165.330 75.820 165.390 ;
        RECT 67.680 165.190 75.820 165.330 ;
        RECT 67.680 165.130 68.000 165.190 ;
        RECT 68.600 165.130 68.920 165.190 ;
        RECT 75.055 165.145 75.345 165.190 ;
        RECT 75.500 165.130 75.820 165.190 ;
        RECT 82.415 165.330 82.705 165.375 ;
        RECT 84.700 165.330 85.020 165.390 ;
        RECT 82.415 165.190 85.020 165.330 ;
        RECT 82.415 165.145 82.705 165.190 ;
        RECT 84.700 165.130 85.020 165.190 ;
        RECT 88.855 165.330 89.145 165.375 ;
        RECT 91.140 165.330 91.460 165.390 ;
        RECT 88.855 165.190 91.460 165.330 ;
        RECT 88.855 165.145 89.145 165.190 ;
        RECT 91.140 165.130 91.460 165.190 ;
        RECT 92.535 165.330 92.825 165.375 ;
        RECT 93.440 165.330 93.760 165.390 ;
        RECT 92.535 165.190 93.760 165.330 ;
        RECT 92.535 165.145 92.825 165.190 ;
        RECT 93.440 165.130 93.760 165.190 ;
        RECT 95.740 165.330 96.060 165.390 ;
        RECT 101.720 165.330 102.040 165.390 ;
        RECT 107.240 165.330 107.560 165.390 ;
        RECT 95.740 165.190 97.350 165.330 ;
        RECT 95.740 165.130 96.060 165.190 ;
        RECT 72.280 164.990 72.600 165.050 ;
        RECT 86.095 164.990 86.385 165.035 ;
        RECT 96.660 164.990 96.980 165.050 ;
        RECT 62.710 164.850 72.600 164.990 ;
        RECT 52.500 164.510 58.340 164.650 ;
        RECT 52.500 164.450 52.820 164.510 ;
        RECT 52.975 164.465 53.265 164.510 ;
        RECT 58.020 164.450 58.340 164.510 ;
        RECT 61.715 164.465 62.005 164.695 ;
        RECT 62.160 164.650 62.480 164.710 ;
        RECT 62.710 164.695 62.850 164.850 ;
        RECT 72.280 164.790 72.600 164.850 ;
        RECT 79.270 164.850 86.385 164.990 ;
        RECT 62.635 164.650 62.925 164.695 ;
        RECT 62.160 164.510 62.925 164.650 ;
        RECT 53.440 164.310 53.730 164.355 ;
        RECT 55.275 164.310 55.565 164.355 ;
        RECT 58.855 164.310 59.145 164.355 ;
        RECT 53.440 164.170 59.145 164.310 ;
        RECT 53.440 164.125 53.730 164.170 ;
        RECT 55.275 164.125 55.565 164.170 ;
        RECT 58.855 164.125 59.145 164.170 ;
        RECT 56.640 164.015 56.960 164.030 ;
        RECT 59.935 164.015 60.225 164.330 ;
        RECT 61.790 164.310 61.930 164.465 ;
        RECT 62.160 164.450 62.480 164.510 ;
        RECT 62.635 164.465 62.925 164.510 ;
        RECT 63.555 164.650 63.845 164.695 ;
        RECT 66.300 164.650 66.620 164.710 ;
        RECT 63.555 164.510 66.620 164.650 ;
        RECT 63.555 164.465 63.845 164.510 ;
        RECT 66.300 164.450 66.620 164.510 ;
        RECT 73.660 164.650 73.980 164.710 ;
        RECT 79.270 164.695 79.410 164.850 ;
        RECT 86.095 164.805 86.385 164.850 ;
        RECT 88.930 164.850 96.980 164.990 ;
        RECT 79.195 164.650 79.485 164.695 ;
        RECT 88.930 164.650 89.070 164.850 ;
        RECT 96.660 164.790 96.980 164.850 ;
        RECT 89.760 164.650 90.080 164.710 ;
        RECT 73.660 164.510 79.485 164.650 ;
        RECT 73.660 164.450 73.980 164.510 ;
        RECT 79.195 164.465 79.485 164.510 ;
        RECT 80.650 164.510 89.070 164.650 ;
        RECT 89.390 164.510 90.080 164.650 ;
        RECT 74.120 164.310 74.440 164.370 ;
        RECT 80.650 164.355 80.790 164.510 ;
        RECT 61.790 164.170 74.440 164.310 ;
        RECT 74.120 164.110 74.440 164.170 ;
        RECT 80.575 164.125 80.865 164.355 ;
        RECT 87.000 164.110 87.320 164.370 ;
        RECT 89.390 164.355 89.530 164.510 ;
        RECT 89.760 164.450 90.080 164.510 ;
        RECT 90.695 164.650 90.985 164.695 ;
        RECT 97.210 164.650 97.350 165.190 ;
        RECT 101.720 165.190 107.560 165.330 ;
        RECT 101.720 165.130 102.040 165.190 ;
        RECT 107.240 165.130 107.560 165.190 ;
        RECT 121.055 165.330 121.345 165.375 ;
        RECT 121.960 165.330 122.280 165.390 ;
        RECT 121.055 165.190 122.280 165.330 ;
        RECT 121.055 165.145 121.345 165.190 ;
        RECT 121.960 165.130 122.280 165.190 ;
        RECT 122.880 165.130 123.200 165.390 ;
        RECT 97.695 164.990 97.985 165.035 ;
        RECT 100.815 164.990 101.105 165.035 ;
        RECT 102.705 164.990 102.995 165.035 ;
        RECT 97.695 164.850 102.995 164.990 ;
        RECT 97.695 164.805 97.985 164.850 ;
        RECT 100.815 164.805 101.105 164.850 ;
        RECT 102.705 164.805 102.995 164.850 ;
        RECT 112.415 164.990 112.705 165.035 ;
        RECT 115.535 164.990 115.825 165.035 ;
        RECT 117.425 164.990 117.715 165.035 ;
        RECT 112.415 164.850 117.715 164.990 ;
        RECT 112.415 164.805 112.705 164.850 ;
        RECT 115.535 164.805 115.825 164.850 ;
        RECT 117.425 164.805 117.715 164.850 ;
        RECT 125.755 164.990 126.045 165.035 ;
        RECT 128.875 164.990 129.165 165.035 ;
        RECT 130.765 164.990 131.055 165.035 ;
        RECT 125.755 164.850 131.055 164.990 ;
        RECT 125.755 164.805 126.045 164.850 ;
        RECT 128.875 164.805 129.165 164.850 ;
        RECT 130.765 164.805 131.055 164.850 ;
        RECT 132.540 164.790 132.860 165.050 ;
        RECT 135.415 164.990 135.705 165.035 ;
        RECT 138.535 164.990 138.825 165.035 ;
        RECT 140.425 164.990 140.715 165.035 ;
        RECT 135.415 164.850 140.715 164.990 ;
        RECT 135.415 164.805 135.705 164.850 ;
        RECT 138.535 164.805 138.825 164.850 ;
        RECT 140.425 164.805 140.715 164.850 ;
        RECT 102.195 164.650 102.485 164.695 ;
        RECT 90.695 164.510 95.970 164.650 ;
        RECT 97.210 164.510 102.485 164.650 ;
        RECT 90.695 164.465 90.985 164.510 ;
        RECT 89.315 164.125 89.605 164.355 ;
        RECT 90.220 164.110 90.540 164.370 ;
        RECT 91.600 164.110 91.920 164.370 ;
        RECT 92.610 164.355 92.750 164.510 ;
        RECT 92.535 164.125 92.825 164.355 ;
        RECT 93.455 164.310 93.745 164.355 ;
        RECT 95.280 164.310 95.600 164.370 ;
        RECT 93.455 164.170 95.600 164.310 ;
        RECT 93.455 164.125 93.745 164.170 ;
        RECT 54.355 163.970 54.645 164.015 ;
        RECT 51.215 163.830 54.645 163.970 ;
        RECT 54.355 163.785 54.645 163.830 ;
        RECT 56.635 163.970 57.285 164.015 ;
        RECT 59.935 163.970 60.525 164.015 ;
        RECT 67.680 163.970 68.000 164.030 ;
        RECT 78.260 163.970 78.580 164.030 ;
        RECT 56.635 163.830 60.525 163.970 ;
        RECT 56.635 163.785 57.285 163.830 ;
        RECT 60.235 163.785 60.525 163.830 ;
        RECT 62.020 163.830 64.230 163.970 ;
        RECT 56.640 163.770 56.960 163.785 ;
        RECT 37.780 163.490 42.610 163.630 ;
        RECT 37.780 163.430 38.100 163.490 ;
        RECT 43.760 163.430 44.080 163.690 ;
        RECT 45.155 163.630 45.445 163.675 ;
        RECT 45.600 163.630 45.920 163.690 ;
        RECT 45.155 163.490 45.920 163.630 ;
        RECT 45.155 163.445 45.445 163.490 ;
        RECT 45.600 163.430 45.920 163.490 ;
        RECT 47.440 163.630 47.760 163.690 ;
        RECT 48.835 163.630 49.125 163.675 ;
        RECT 47.440 163.490 49.125 163.630 ;
        RECT 47.440 163.430 47.760 163.490 ;
        RECT 48.835 163.445 49.125 163.490 ;
        RECT 51.135 163.630 51.425 163.675 ;
        RECT 54.800 163.630 55.120 163.690 ;
        RECT 51.135 163.490 55.120 163.630 ;
        RECT 51.135 163.445 51.425 163.490 ;
        RECT 54.800 163.430 55.120 163.490 ;
        RECT 58.940 163.630 59.260 163.690 ;
        RECT 62.020 163.630 62.160 163.830 ;
        RECT 64.090 163.675 64.230 163.830 ;
        RECT 67.680 163.830 78.580 163.970 ;
        RECT 67.680 163.770 68.000 163.830 ;
        RECT 78.260 163.770 78.580 163.830 ;
        RECT 78.720 163.970 79.040 164.030 ;
        RECT 83.335 163.970 83.625 164.015 ;
        RECT 78.720 163.830 83.625 163.970 ;
        RECT 90.310 163.970 90.450 164.110 ;
        RECT 93.530 163.970 93.670 164.125 ;
        RECT 95.280 164.110 95.600 164.170 ;
        RECT 90.310 163.830 93.670 163.970 ;
        RECT 78.720 163.770 79.040 163.830 ;
        RECT 83.335 163.785 83.625 163.830 ;
        RECT 58.940 163.490 62.160 163.630 ;
        RECT 58.940 163.430 59.260 163.490 ;
        RECT 64.015 163.445 64.305 163.675 ;
        RECT 74.580 163.630 74.900 163.690 ;
        RECT 80.115 163.630 80.405 163.675 ;
        RECT 81.940 163.630 82.260 163.690 ;
        RECT 74.580 163.490 82.260 163.630 ;
        RECT 74.580 163.430 74.900 163.490 ;
        RECT 80.115 163.445 80.405 163.490 ;
        RECT 81.940 163.430 82.260 163.490 ;
        RECT 82.860 163.630 83.180 163.690 ;
        RECT 83.795 163.630 84.085 163.675 ;
        RECT 82.860 163.490 84.085 163.630 ;
        RECT 82.860 163.430 83.180 163.490 ;
        RECT 83.795 163.445 84.085 163.490 ;
        RECT 86.540 163.630 86.860 163.690 ;
        RECT 94.820 163.630 95.140 163.690 ;
        RECT 86.540 163.490 95.140 163.630 ;
        RECT 95.830 163.630 95.970 164.510 ;
        RECT 102.195 164.465 102.485 164.510 ;
        RECT 103.575 164.650 103.865 164.695 ;
        RECT 115.060 164.650 115.380 164.710 ;
        RECT 116.900 164.650 117.220 164.710 ;
        RECT 118.295 164.650 118.585 164.695 ;
        RECT 131.635 164.650 131.925 164.695 ;
        RECT 133.920 164.650 134.240 164.710 ;
        RECT 103.575 164.510 141.510 164.650 ;
        RECT 103.575 164.465 103.865 164.510 ;
        RECT 115.060 164.450 115.380 164.510 ;
        RECT 116.900 164.450 117.220 164.510 ;
        RECT 118.295 164.465 118.585 164.510 ;
        RECT 131.635 164.465 131.925 164.510 ;
        RECT 133.920 164.450 134.240 164.510 ;
        RECT 96.615 164.015 96.905 164.330 ;
        RECT 97.695 164.310 97.985 164.355 ;
        RECT 101.275 164.310 101.565 164.355 ;
        RECT 103.110 164.310 103.400 164.355 ;
        RECT 97.695 164.170 103.400 164.310 ;
        RECT 97.695 164.125 97.985 164.170 ;
        RECT 101.275 164.125 101.565 164.170 ;
        RECT 103.110 164.125 103.400 164.170 ;
        RECT 107.715 164.125 108.005 164.355 ;
        RECT 96.315 163.970 96.905 164.015 ;
        RECT 99.555 163.970 100.205 164.015 ;
        RECT 100.800 163.970 101.120 164.030 ;
        RECT 96.315 163.830 103.330 163.970 ;
        RECT 96.315 163.785 96.605 163.830 ;
        RECT 99.555 163.785 100.205 163.830 ;
        RECT 100.800 163.770 101.120 163.830 ;
        RECT 103.190 163.690 103.330 163.830 ;
        RECT 97.580 163.630 97.900 163.690 ;
        RECT 95.830 163.490 97.900 163.630 ;
        RECT 86.540 163.430 86.860 163.490 ;
        RECT 94.820 163.430 95.140 163.490 ;
        RECT 97.580 163.430 97.900 163.490 ;
        RECT 103.100 163.430 103.420 163.690 ;
        RECT 104.480 163.430 104.800 163.690 ;
        RECT 107.790 163.630 107.930 164.125 ;
        RECT 108.160 164.110 108.480 164.370 ;
        RECT 141.370 164.355 141.510 164.510 ;
        RECT 111.335 164.015 111.625 164.330 ;
        RECT 112.415 164.310 112.705 164.355 ;
        RECT 115.995 164.310 116.285 164.355 ;
        RECT 117.830 164.310 118.120 164.355 ;
        RECT 112.415 164.170 118.120 164.310 ;
        RECT 112.415 164.125 112.705 164.170 ;
        RECT 115.995 164.125 116.285 164.170 ;
        RECT 117.830 164.125 118.120 164.170 ;
        RECT 114.600 164.015 114.920 164.030 ;
        RECT 111.035 163.970 111.625 164.015 ;
        RECT 114.275 163.970 114.925 164.015 ;
        RECT 111.035 163.830 114.925 163.970 ;
        RECT 111.035 163.785 111.325 163.830 ;
        RECT 114.275 163.785 114.925 163.830 ;
        RECT 116.915 163.785 117.205 164.015 ;
        RECT 117.360 163.970 117.680 164.030 ;
        RECT 124.675 164.015 124.965 164.330 ;
        RECT 125.755 164.310 126.045 164.355 ;
        RECT 129.335 164.310 129.625 164.355 ;
        RECT 131.170 164.310 131.460 164.355 ;
        RECT 125.755 164.170 131.460 164.310 ;
        RECT 125.755 164.125 126.045 164.170 ;
        RECT 129.335 164.125 129.625 164.170 ;
        RECT 131.170 164.125 131.460 164.170 ;
        RECT 119.675 163.970 119.965 164.015 ;
        RECT 124.375 163.970 124.965 164.015 ;
        RECT 127.615 163.970 128.265 164.015 ;
        RECT 128.860 163.970 129.180 164.030 ;
        RECT 117.360 163.830 119.965 163.970 ;
        RECT 114.600 163.770 114.920 163.785 ;
        RECT 115.520 163.630 115.840 163.690 ;
        RECT 107.790 163.490 115.840 163.630 ;
        RECT 116.990 163.630 117.130 163.785 ;
        RECT 117.360 163.770 117.680 163.830 ;
        RECT 119.675 163.785 119.965 163.830 ;
        RECT 122.510 163.830 124.030 163.970 ;
        RECT 122.510 163.630 122.650 163.830 ;
        RECT 116.990 163.490 122.650 163.630 ;
        RECT 123.890 163.630 124.030 163.830 ;
        RECT 124.375 163.830 129.180 163.970 ;
        RECT 124.375 163.785 124.665 163.830 ;
        RECT 127.615 163.785 128.265 163.830 ;
        RECT 128.860 163.770 129.180 163.830 ;
        RECT 130.240 163.770 130.560 164.030 ;
        RECT 134.335 164.015 134.625 164.330 ;
        RECT 135.415 164.310 135.705 164.355 ;
        RECT 138.995 164.310 139.285 164.355 ;
        RECT 140.830 164.310 141.120 164.355 ;
        RECT 135.415 164.170 141.120 164.310 ;
        RECT 135.415 164.125 135.705 164.170 ;
        RECT 138.995 164.125 139.285 164.170 ;
        RECT 140.830 164.125 141.120 164.170 ;
        RECT 141.295 164.310 141.585 164.355 ;
        RECT 144.040 164.310 144.360 164.370 ;
        RECT 141.295 164.170 144.360 164.310 ;
        RECT 141.295 164.125 141.585 164.170 ;
        RECT 144.040 164.110 144.360 164.170 ;
        RECT 145.420 164.310 145.740 164.370 ;
        RECT 146.815 164.310 147.105 164.355 ;
        RECT 145.420 164.170 147.105 164.310 ;
        RECT 145.420 164.110 145.740 164.170 ;
        RECT 146.815 164.125 147.105 164.170 ;
        RECT 149.115 164.310 149.405 164.355 ;
        RECT 150.940 164.310 151.260 164.370 ;
        RECT 149.115 164.170 151.260 164.310 ;
        RECT 149.115 164.125 149.405 164.170 ;
        RECT 137.600 164.015 137.920 164.030 ;
        RECT 134.035 163.970 134.625 164.015 ;
        RECT 137.275 163.970 137.925 164.015 ;
        RECT 138.520 163.970 138.840 164.030 ;
        RECT 139.915 163.970 140.205 164.015 ;
        RECT 134.035 163.830 138.290 163.970 ;
        RECT 134.035 163.785 134.325 163.830 ;
        RECT 137.275 163.785 137.925 163.830 ;
        RECT 137.600 163.770 137.920 163.785 ;
        RECT 128.400 163.630 128.720 163.690 ;
        RECT 123.890 163.490 128.720 163.630 ;
        RECT 138.150 163.630 138.290 163.830 ;
        RECT 138.520 163.830 140.205 163.970 ;
        RECT 138.520 163.770 138.840 163.830 ;
        RECT 139.915 163.785 140.205 163.830 ;
        RECT 144.960 163.770 145.280 164.030 ;
        RECT 145.050 163.630 145.190 163.770 ;
        RECT 138.150 163.490 145.190 163.630 ;
        RECT 146.890 163.630 147.030 164.125 ;
        RECT 150.940 164.110 151.260 164.170 ;
        RECT 148.195 163.630 148.485 163.675 ;
        RECT 146.890 163.490 148.485 163.630 ;
        RECT 115.520 163.430 115.840 163.490 ;
        RECT 128.400 163.430 128.720 163.490 ;
        RECT 148.195 163.445 148.485 163.490 ;
        RECT 2.750 162.810 159.030 163.290 ;
        RECT 5.135 162.610 5.425 162.655 ;
        RECT 2.450 162.470 5.425 162.610 ;
        RECT 5.135 162.425 5.425 162.470 ;
        RECT 6.515 162.425 6.805 162.655 ;
        RECT 8.815 162.610 9.105 162.655 ;
        RECT 12.940 162.610 13.260 162.670 ;
        RECT 13.860 162.610 14.180 162.670 ;
        RECT 8.815 162.470 13.260 162.610 ;
        RECT 8.815 162.425 9.105 162.470 ;
        RECT 6.055 161.930 6.345 161.975 ;
        RECT 6.590 161.930 6.730 162.425 ;
        RECT 12.940 162.410 13.260 162.470 ;
        RECT 13.720 162.410 14.180 162.610 ;
        RECT 18.460 162.610 18.780 162.670 ;
        RECT 19.855 162.610 20.145 162.655 ;
        RECT 18.460 162.470 20.145 162.610 ;
        RECT 18.460 162.410 18.780 162.470 ;
        RECT 19.855 162.425 20.145 162.470 ;
        RECT 24.900 162.410 25.220 162.670 ;
        RECT 26.280 162.410 26.600 162.670 ;
        RECT 35.020 162.610 35.340 162.670 ;
        RECT 37.780 162.610 38.100 162.670 ;
        RECT 35.020 162.470 38.100 162.610 ;
        RECT 35.020 162.410 35.340 162.470 ;
        RECT 37.780 162.410 38.100 162.470 ;
        RECT 41.460 162.410 41.780 162.670 ;
        RECT 45.140 162.610 45.460 162.670 ;
        RECT 45.140 162.470 49.050 162.610 ;
        RECT 45.140 162.410 45.460 162.470 ;
        RECT 11.560 162.270 11.880 162.330 ;
        RECT 9.810 162.130 11.880 162.270 ;
        RECT 6.055 161.790 6.730 161.930 ;
        RECT 6.055 161.745 6.345 161.790 ;
        RECT 8.355 161.745 8.645 161.975 ;
        RECT 8.430 161.250 8.570 161.745 ;
        RECT 9.810 161.635 9.950 162.130 ;
        RECT 11.560 162.070 11.880 162.130 ;
        RECT 12.035 162.270 12.325 162.315 ;
        RECT 13.720 162.270 13.860 162.410 ;
        RECT 12.035 162.130 13.860 162.270 ;
        RECT 14.315 162.270 14.965 162.315 ;
        RECT 17.915 162.270 18.205 162.315 ;
        RECT 24.990 162.270 25.130 162.410 ;
        RECT 14.315 162.130 18.205 162.270 ;
        RECT 12.035 162.085 12.325 162.130 ;
        RECT 14.315 162.085 14.965 162.130 ;
        RECT 17.615 162.085 18.205 162.130 ;
        RECT 23.610 162.130 25.130 162.270 ;
        RECT 10.640 161.730 10.960 161.990 ;
        RECT 11.120 161.930 11.410 161.975 ;
        RECT 12.955 161.930 13.245 161.975 ;
        RECT 16.535 161.930 16.825 161.975 ;
        RECT 11.120 161.790 16.825 161.930 ;
        RECT 11.120 161.745 11.410 161.790 ;
        RECT 12.955 161.745 13.245 161.790 ;
        RECT 16.535 161.745 16.825 161.790 ;
        RECT 17.615 161.770 17.905 162.085 ;
        RECT 23.610 161.975 23.750 162.130 ;
        RECT 41.000 162.070 41.320 162.330 ;
        RECT 48.910 162.315 49.050 162.470 ;
        RECT 51.120 162.410 51.440 162.670 ;
        RECT 52.040 162.610 52.360 162.670 ;
        RECT 54.815 162.610 55.105 162.655 ;
        RECT 52.040 162.470 55.105 162.610 ;
        RECT 52.040 162.410 52.360 162.470 ;
        RECT 54.815 162.425 55.105 162.470 ;
        RECT 58.035 162.610 58.325 162.655 ;
        RECT 58.940 162.610 59.260 162.670 ;
        RECT 58.035 162.470 59.260 162.610 ;
        RECT 58.035 162.425 58.325 162.470 ;
        RECT 58.940 162.410 59.260 162.470 ;
        RECT 59.400 162.610 59.720 162.670 ;
        RECT 72.755 162.610 73.045 162.655 ;
        RECT 73.200 162.610 73.520 162.670 ;
        RECT 59.400 162.470 65.610 162.610 ;
        RECT 59.400 162.410 59.720 162.470 ;
        RECT 42.955 162.270 43.245 162.315 ;
        RECT 46.195 162.270 46.845 162.315 ;
        RECT 42.955 162.130 46.845 162.270 ;
        RECT 42.955 162.085 43.545 162.130 ;
        RECT 46.195 162.085 46.845 162.130 ;
        RECT 48.835 162.085 49.125 162.315 ;
        RECT 52.500 162.270 52.820 162.330 ;
        RECT 60.795 162.270 61.085 162.315 ;
        RECT 63.080 162.270 63.400 162.330 ;
        RECT 65.470 162.315 65.610 162.470 ;
        RECT 72.755 162.470 73.520 162.610 ;
        RECT 72.755 162.425 73.045 162.470 ;
        RECT 73.200 162.410 73.520 162.470 ;
        RECT 74.120 162.610 74.440 162.670 ;
        RECT 74.595 162.610 74.885 162.655 ;
        RECT 74.120 162.470 74.885 162.610 ;
        RECT 74.120 162.410 74.440 162.470 ;
        RECT 74.595 162.425 74.885 162.470 ;
        RECT 75.055 162.610 75.345 162.655 ;
        RECT 75.960 162.610 76.280 162.670 ;
        RECT 75.055 162.470 76.280 162.610 ;
        RECT 75.055 162.425 75.345 162.470 ;
        RECT 75.960 162.410 76.280 162.470 ;
        RECT 76.895 162.610 77.185 162.655 ;
        RECT 76.895 162.470 84.010 162.610 ;
        RECT 76.895 162.425 77.185 162.470 ;
        RECT 52.500 162.130 59.170 162.270 ;
        RECT 43.255 161.990 43.545 162.085 ;
        RECT 52.500 162.070 52.820 162.130 ;
        RECT 9.735 161.405 10.025 161.635 ;
        RECT 13.860 161.590 14.180 161.650 ;
        RECT 17.080 161.590 17.400 161.650 ;
        RECT 11.190 161.450 17.400 161.590 ;
        RECT 11.190 161.250 11.330 161.450 ;
        RECT 13.860 161.390 14.180 161.450 ;
        RECT 17.080 161.390 17.400 161.450 ;
        RECT 8.430 161.110 11.330 161.250 ;
        RECT 11.525 161.250 11.815 161.295 ;
        RECT 13.415 161.250 13.705 161.295 ;
        RECT 16.535 161.250 16.825 161.295 ;
        RECT 11.525 161.110 16.825 161.250 ;
        RECT 11.525 161.065 11.815 161.110 ;
        RECT 13.415 161.065 13.705 161.110 ;
        RECT 16.535 161.065 16.825 161.110 ;
        RECT 17.630 160.970 17.770 161.770 ;
        RECT 23.535 161.745 23.825 161.975 ;
        RECT 24.440 161.730 24.760 161.990 ;
        RECT 24.915 161.745 25.205 161.975 ;
        RECT 25.375 161.930 25.665 161.975 ;
        RECT 26.740 161.930 27.060 161.990 ;
        RECT 25.375 161.790 27.060 161.930 ;
        RECT 25.375 161.745 25.665 161.790 ;
        RECT 19.395 161.590 19.685 161.635 ;
        RECT 22.615 161.590 22.905 161.635 ;
        RECT 24.990 161.590 25.130 161.745 ;
        RECT 26.740 161.730 27.060 161.790 ;
        RECT 30.895 161.930 31.185 161.975 ;
        RECT 35.020 161.930 35.340 161.990 ;
        RECT 30.895 161.790 38.010 161.930 ;
        RECT 30.895 161.745 31.185 161.790 ;
        RECT 35.020 161.730 35.340 161.790 ;
        RECT 19.395 161.450 25.130 161.590 ;
        RECT 31.815 161.590 32.105 161.635 ;
        RECT 37.320 161.590 37.640 161.650 ;
        RECT 31.815 161.450 37.640 161.590 ;
        RECT 37.870 161.590 38.010 161.790 ;
        RECT 43.255 161.770 43.620 161.990 ;
        RECT 43.300 161.730 43.620 161.770 ;
        RECT 44.335 161.930 44.625 161.975 ;
        RECT 47.915 161.930 48.205 161.975 ;
        RECT 49.750 161.930 50.040 161.975 ;
        RECT 44.335 161.790 50.040 161.930 ;
        RECT 44.335 161.745 44.625 161.790 ;
        RECT 47.915 161.745 48.205 161.790 ;
        RECT 49.750 161.745 50.040 161.790 ;
        RECT 50.215 161.930 50.505 161.975 ;
        RECT 50.660 161.930 50.980 161.990 ;
        RECT 50.215 161.790 50.980 161.930 ;
        RECT 50.215 161.745 50.505 161.790 ;
        RECT 50.660 161.730 50.980 161.790 ;
        RECT 52.055 161.930 52.345 161.975 ;
        RECT 55.260 161.930 55.580 161.990 ;
        RECT 56.180 161.930 56.500 161.990 ;
        RECT 52.055 161.790 55.030 161.930 ;
        RECT 52.055 161.745 52.345 161.790 ;
        RECT 39.620 161.590 39.940 161.650 ;
        RECT 43.760 161.590 44.080 161.650 ;
        RECT 37.870 161.450 44.080 161.590 ;
        RECT 19.395 161.405 19.685 161.450 ;
        RECT 22.615 161.405 22.905 161.450 ;
        RECT 31.815 161.405 32.105 161.450 ;
        RECT 37.320 161.390 37.640 161.450 ;
        RECT 39.620 161.390 39.940 161.450 ;
        RECT 43.760 161.390 44.080 161.450 ;
        RECT 52.515 161.405 52.805 161.635 ;
        RECT 52.975 161.405 53.265 161.635 ;
        RECT 53.435 161.590 53.725 161.635 ;
        RECT 54.340 161.590 54.660 161.650 ;
        RECT 53.435 161.450 54.660 161.590 ;
        RECT 54.890 161.590 55.030 161.790 ;
        RECT 55.260 161.790 56.500 161.930 ;
        RECT 55.260 161.730 55.580 161.790 ;
        RECT 56.180 161.730 56.500 161.790 ;
        RECT 57.100 161.730 57.420 161.990 ;
        RECT 57.560 161.730 57.880 161.990 ;
        RECT 59.030 161.975 59.170 162.130 ;
        RECT 60.795 162.130 63.400 162.270 ;
        RECT 60.795 162.085 61.085 162.130 ;
        RECT 63.080 162.070 63.400 162.130 ;
        RECT 65.395 162.085 65.685 162.315 ;
        RECT 67.675 162.270 68.325 162.315 ;
        RECT 69.060 162.270 69.380 162.330 ;
        RECT 71.275 162.270 71.565 162.315 ;
        RECT 67.675 162.130 71.565 162.270 ;
        RECT 67.675 162.085 68.325 162.130 ;
        RECT 69.060 162.070 69.380 162.130 ;
        RECT 70.975 162.085 71.565 162.130 ;
        RECT 77.355 162.270 77.645 162.315 ;
        RECT 78.720 162.270 79.040 162.330 ;
        RECT 77.355 162.130 79.040 162.270 ;
        RECT 77.355 162.085 77.645 162.130 ;
        RECT 58.955 161.745 59.245 161.975 ;
        RECT 60.335 161.930 60.625 161.975 ;
        RECT 61.700 161.930 62.020 161.990 ;
        RECT 60.335 161.790 62.020 161.930 ;
        RECT 60.335 161.745 60.625 161.790 ;
        RECT 61.700 161.730 62.020 161.790 ;
        RECT 64.480 161.930 64.770 161.975 ;
        RECT 66.315 161.930 66.605 161.975 ;
        RECT 69.895 161.930 70.185 161.975 ;
        RECT 64.480 161.790 70.185 161.930 ;
        RECT 64.480 161.745 64.770 161.790 ;
        RECT 66.315 161.745 66.605 161.790 ;
        RECT 69.895 161.745 70.185 161.790 ;
        RECT 70.440 161.930 70.760 161.990 ;
        RECT 70.975 161.930 71.265 162.085 ;
        RECT 77.430 161.930 77.570 162.085 ;
        RECT 78.720 162.070 79.040 162.130 ;
        RECT 79.195 162.270 79.485 162.315 ;
        RECT 81.480 162.270 81.800 162.330 ;
        RECT 79.195 162.130 81.800 162.270 ;
        RECT 79.195 162.085 79.485 162.130 ;
        RECT 81.480 162.070 81.800 162.130 ;
        RECT 81.940 162.270 82.260 162.330 ;
        RECT 83.870 162.270 84.010 162.470 ;
        RECT 84.240 162.410 84.560 162.670 ;
        RECT 86.555 162.610 86.845 162.655 ;
        RECT 89.300 162.610 89.620 162.670 ;
        RECT 86.555 162.470 89.620 162.610 ;
        RECT 86.555 162.425 86.845 162.470 ;
        RECT 89.300 162.410 89.620 162.470 ;
        RECT 92.060 162.410 92.380 162.670 ;
        RECT 92.520 162.410 92.840 162.670 ;
        RECT 92.980 162.610 93.300 162.670 ;
        RECT 94.375 162.610 94.665 162.655 ;
        RECT 95.740 162.610 96.060 162.670 ;
        RECT 92.980 162.470 96.060 162.610 ;
        RECT 92.980 162.410 93.300 162.470 ;
        RECT 94.375 162.425 94.665 162.470 ;
        RECT 95.740 162.410 96.060 162.470 ;
        RECT 97.120 162.610 97.440 162.670 ;
        RECT 98.500 162.610 98.820 162.670 ;
        RECT 108.160 162.610 108.480 162.670 ;
        RECT 113.220 162.610 113.540 162.670 ;
        RECT 121.055 162.610 121.345 162.655 ;
        RECT 97.120 162.470 98.820 162.610 ;
        RECT 97.120 162.410 97.440 162.470 ;
        RECT 98.500 162.410 98.820 162.470 ;
        RECT 99.510 162.470 106.550 162.610 ;
        RECT 92.150 162.270 92.290 162.410 ;
        RECT 81.940 162.130 82.630 162.270 ;
        RECT 83.870 162.130 92.290 162.270 ;
        RECT 92.610 162.270 92.750 162.410 ;
        RECT 99.510 162.315 99.650 162.470 ;
        RECT 95.295 162.270 95.585 162.315 ;
        RECT 92.610 162.130 95.585 162.270 ;
        RECT 81.940 162.070 82.260 162.130 ;
        RECT 70.440 161.790 77.570 161.930 ;
        RECT 77.800 161.930 78.120 161.990 ;
        RECT 82.490 161.975 82.630 162.130 ;
        RECT 95.295 162.085 95.585 162.130 ;
        RECT 99.435 162.085 99.725 162.315 ;
        RECT 102.640 162.270 102.960 162.330 ;
        RECT 104.940 162.270 105.260 162.330 ;
        RECT 106.410 162.315 106.550 162.470 ;
        RECT 108.160 162.470 113.540 162.610 ;
        RECT 108.160 162.410 108.480 162.470 ;
        RECT 113.220 162.410 113.540 162.470 ;
        RECT 118.370 162.470 121.345 162.610 ;
        RECT 102.640 162.130 105.260 162.270 ;
        RECT 77.800 161.790 81.710 161.930 ;
        RECT 70.440 161.730 70.760 161.790 ;
        RECT 70.975 161.770 71.265 161.790 ;
        RECT 77.800 161.730 78.120 161.790 ;
        RECT 55.720 161.590 56.040 161.650 ;
        RECT 54.890 161.450 56.040 161.590 ;
        RECT 53.435 161.405 53.725 161.450 ;
        RECT 24.440 161.250 24.760 161.310 ;
        RECT 29.975 161.250 30.265 161.295 ;
        RECT 24.440 161.110 30.265 161.250 ;
        RECT 24.440 161.050 24.760 161.110 ;
        RECT 29.975 161.065 30.265 161.110 ;
        RECT 44.335 161.250 44.625 161.295 ;
        RECT 47.455 161.250 47.745 161.295 ;
        RECT 49.345 161.250 49.635 161.295 ;
        RECT 44.335 161.110 49.635 161.250 ;
        RECT 44.335 161.065 44.625 161.110 ;
        RECT 47.455 161.065 47.745 161.110 ;
        RECT 49.345 161.065 49.635 161.110 ;
        RECT 8.800 160.910 9.120 160.970 ;
        RECT 17.540 160.910 17.860 160.970 ;
        RECT 8.800 160.770 17.860 160.910 ;
        RECT 8.800 160.710 9.120 160.770 ;
        RECT 17.540 160.710 17.860 160.770 ;
        RECT 34.560 160.710 34.880 160.970 ;
        RECT 36.860 160.910 37.180 160.970 ;
        RECT 49.740 160.910 50.060 160.970 ;
        RECT 36.860 160.770 50.060 160.910 ;
        RECT 52.590 160.910 52.730 161.405 ;
        RECT 53.050 161.250 53.190 161.405 ;
        RECT 54.340 161.390 54.660 161.450 ;
        RECT 55.720 161.390 56.040 161.450 ;
        RECT 56.655 161.405 56.945 161.635 ;
        RECT 56.730 161.250 56.870 161.405 ;
        RECT 57.650 161.250 57.790 161.730 ;
        RECT 58.020 161.590 58.340 161.650 ;
        RECT 60.795 161.590 61.085 161.635 ;
        RECT 58.020 161.450 61.085 161.590 ;
        RECT 58.020 161.390 58.340 161.450 ;
        RECT 60.795 161.405 61.085 161.450 ;
        RECT 62.620 161.590 62.940 161.650 ;
        RECT 64.015 161.590 64.305 161.635 ;
        RECT 68.600 161.590 68.920 161.650 ;
        RECT 62.620 161.450 68.920 161.590 ;
        RECT 62.620 161.390 62.940 161.450 ;
        RECT 64.015 161.405 64.305 161.450 ;
        RECT 68.600 161.390 68.920 161.450 ;
        RECT 72.280 161.390 72.600 161.650 ;
        RECT 73.660 161.390 73.980 161.650 ;
        RECT 81.035 161.405 81.325 161.635 ;
        RECT 53.050 161.110 57.790 161.250 ;
        RECT 59.400 161.250 59.720 161.310 ;
        RECT 61.700 161.250 62.020 161.310 ;
        RECT 64.885 161.250 65.175 161.295 ;
        RECT 66.775 161.250 67.065 161.295 ;
        RECT 69.895 161.250 70.185 161.295 ;
        RECT 59.400 161.110 62.020 161.250 ;
        RECT 59.400 161.050 59.720 161.110 ;
        RECT 61.700 161.050 62.020 161.110 ;
        RECT 62.710 161.110 64.695 161.250 ;
        RECT 55.260 160.910 55.580 160.970 ;
        RECT 52.590 160.770 55.580 160.910 ;
        RECT 36.860 160.710 37.180 160.770 ;
        RECT 49.740 160.710 50.060 160.770 ;
        RECT 55.260 160.710 55.580 160.770 ;
        RECT 55.720 160.910 56.040 160.970 ;
        RECT 62.710 160.910 62.850 161.110 ;
        RECT 55.720 160.770 62.850 160.910 ;
        RECT 63.095 160.910 63.385 160.955 ;
        RECT 63.540 160.910 63.860 160.970 ;
        RECT 63.095 160.770 63.860 160.910 ;
        RECT 64.555 160.910 64.695 161.110 ;
        RECT 64.885 161.110 70.185 161.250 ;
        RECT 72.370 161.250 72.510 161.390 ;
        RECT 81.110 161.250 81.250 161.405 ;
        RECT 72.370 161.110 81.250 161.250 ;
        RECT 81.570 161.250 81.710 161.790 ;
        RECT 82.415 161.745 82.705 161.975 ;
        RECT 86.080 161.730 86.400 161.990 ;
        RECT 86.540 161.930 86.860 161.990 ;
        RECT 87.015 161.930 87.305 161.975 ;
        RECT 86.540 161.790 87.305 161.930 ;
        RECT 86.540 161.730 86.860 161.790 ;
        RECT 87.015 161.745 87.305 161.790 ;
        RECT 87.475 161.930 87.765 161.975 ;
        RECT 89.775 161.930 90.065 161.975 ;
        RECT 87.475 161.790 90.065 161.930 ;
        RECT 87.475 161.745 87.765 161.790 ;
        RECT 89.775 161.745 90.065 161.790 ;
        RECT 81.940 161.390 82.260 161.650 ;
        RECT 86.170 161.590 86.310 161.730 ;
        RECT 88.855 161.590 89.145 161.635 ;
        RECT 86.170 161.450 89.145 161.590 ;
        RECT 89.850 161.590 89.990 161.745 ;
        RECT 90.220 161.730 90.540 161.990 ;
        RECT 91.140 161.730 91.460 161.990 ;
        RECT 92.075 161.930 92.365 161.975 ;
        RECT 93.455 161.930 93.745 161.975 ;
        RECT 94.360 161.930 94.680 161.990 ;
        RECT 99.510 161.930 99.650 162.085 ;
        RECT 102.640 162.070 102.960 162.130 ;
        RECT 104.940 162.070 105.260 162.130 ;
        RECT 106.335 162.085 106.625 162.315 ;
        RECT 109.195 162.270 109.485 162.315 ;
        RECT 112.435 162.270 113.085 162.315 ;
        RECT 114.600 162.270 114.920 162.330 ;
        RECT 109.195 162.130 114.920 162.270 ;
        RECT 109.195 162.085 109.785 162.130 ;
        RECT 112.435 162.085 113.085 162.130 ;
        RECT 92.075 161.790 94.680 161.930 ;
        RECT 92.075 161.745 92.365 161.790 ;
        RECT 93.455 161.745 93.745 161.790 ;
        RECT 92.150 161.590 92.290 161.745 ;
        RECT 94.360 161.730 94.680 161.790 ;
        RECT 95.830 161.790 99.650 161.930 ;
        RECT 101.275 161.930 101.565 161.975 ;
        RECT 103.575 161.930 103.865 161.975 ;
        RECT 101.275 161.790 103.865 161.930 ;
        RECT 89.850 161.450 92.290 161.590 ;
        RECT 88.855 161.405 89.145 161.450 ;
        RECT 85.635 161.250 85.925 161.295 ;
        RECT 81.570 161.110 85.925 161.250 ;
        RECT 64.885 161.065 65.175 161.110 ;
        RECT 66.775 161.065 67.065 161.110 ;
        RECT 69.895 161.065 70.185 161.110 ;
        RECT 77.800 160.910 78.120 160.970 ;
        RECT 64.555 160.770 78.120 160.910 ;
        RECT 81.110 160.910 81.250 161.110 ;
        RECT 85.635 161.065 85.925 161.110 ;
        RECT 88.380 161.050 88.700 161.310 ;
        RECT 95.830 161.250 95.970 161.790 ;
        RECT 101.275 161.745 101.565 161.790 ;
        RECT 103.575 161.745 103.865 161.790 ;
        RECT 109.495 161.770 109.785 162.085 ;
        RECT 114.600 162.070 114.920 162.130 ;
        RECT 115.075 162.270 115.365 162.315 ;
        RECT 118.370 162.270 118.510 162.470 ;
        RECT 121.055 162.425 121.345 162.470 ;
        RECT 122.880 162.610 123.200 162.670 ;
        RECT 126.115 162.610 126.405 162.655 ;
        RECT 122.880 162.470 126.405 162.610 ;
        RECT 122.880 162.410 123.200 162.470 ;
        RECT 126.115 162.425 126.405 162.470 ;
        RECT 127.955 162.425 128.245 162.655 ;
        RECT 128.030 162.270 128.170 162.425 ;
        RECT 128.400 162.410 128.720 162.670 ;
        RECT 130.240 162.610 130.560 162.670 ;
        RECT 130.715 162.610 131.005 162.655 ;
        RECT 130.240 162.470 131.005 162.610 ;
        RECT 130.240 162.410 130.560 162.470 ;
        RECT 130.715 162.425 131.005 162.470 ;
        RECT 132.540 162.610 132.860 162.670 ;
        RECT 133.935 162.610 134.225 162.655 ;
        RECT 132.540 162.470 134.225 162.610 ;
        RECT 132.540 162.410 132.860 162.470 ;
        RECT 133.935 162.425 134.225 162.470 ;
        RECT 135.775 162.425 136.065 162.655 ;
        RECT 137.155 162.610 137.445 162.655 ;
        RECT 138.520 162.610 138.840 162.670 ;
        RECT 144.960 162.610 145.280 162.670 ;
        RECT 137.155 162.470 138.840 162.610 ;
        RECT 137.155 162.425 137.445 162.470 ;
        RECT 115.075 162.130 118.510 162.270 ;
        RECT 119.290 162.130 124.950 162.270 ;
        RECT 128.030 162.130 130.010 162.270 ;
        RECT 115.075 162.085 115.365 162.130 ;
        RECT 119.290 161.990 119.430 162.130 ;
        RECT 110.575 161.930 110.865 161.975 ;
        RECT 114.155 161.930 114.445 161.975 ;
        RECT 115.990 161.930 116.280 161.975 ;
        RECT 110.575 161.790 116.280 161.930 ;
        RECT 110.575 161.745 110.865 161.790 ;
        RECT 114.155 161.745 114.445 161.790 ;
        RECT 115.990 161.745 116.280 161.790 ;
        RECT 116.455 161.930 116.745 161.975 ;
        RECT 116.900 161.930 117.220 161.990 ;
        RECT 118.755 161.930 119.045 161.975 ;
        RECT 116.455 161.790 117.220 161.930 ;
        RECT 116.455 161.745 116.745 161.790 ;
        RECT 96.660 161.590 96.980 161.650 ;
        RECT 98.055 161.590 98.345 161.635 ;
        RECT 96.660 161.450 98.345 161.590 ;
        RECT 96.660 161.390 96.980 161.450 ;
        RECT 98.055 161.405 98.345 161.450 ;
        RECT 90.310 161.110 95.970 161.250 ;
        RECT 90.310 160.910 90.450 161.110 ;
        RECT 81.110 160.770 90.450 160.910 ;
        RECT 90.680 160.910 91.000 160.970 ;
        RECT 91.615 160.910 91.905 160.955 ;
        RECT 90.680 160.770 91.905 160.910 ;
        RECT 55.720 160.710 56.040 160.770 ;
        RECT 63.095 160.725 63.385 160.770 ;
        RECT 63.540 160.710 63.860 160.770 ;
        RECT 77.800 160.710 78.120 160.770 ;
        RECT 90.680 160.710 91.000 160.770 ;
        RECT 91.615 160.725 91.905 160.770 ;
        RECT 94.820 160.910 95.140 160.970 ;
        RECT 96.200 160.910 96.520 160.970 ;
        RECT 101.350 160.910 101.490 161.745 ;
        RECT 116.900 161.730 117.220 161.790 ;
        RECT 117.450 161.790 119.045 161.930 ;
        RECT 102.640 161.390 102.960 161.650 ;
        RECT 103.115 161.590 103.405 161.635 ;
        RECT 108.160 161.590 108.480 161.650 ;
        RECT 112.300 161.590 112.620 161.650 ;
        RECT 103.115 161.450 112.620 161.590 ;
        RECT 103.115 161.405 103.405 161.450 ;
        RECT 108.160 161.390 108.480 161.450 ;
        RECT 112.300 161.390 112.620 161.450 ;
        RECT 113.220 161.590 113.540 161.650 ;
        RECT 117.450 161.590 117.590 161.790 ;
        RECT 118.755 161.745 119.045 161.790 ;
        RECT 113.220 161.450 117.590 161.590 ;
        RECT 113.220 161.390 113.540 161.450 ;
        RECT 117.835 161.405 118.125 161.635 ;
        RECT 110.575 161.250 110.865 161.295 ;
        RECT 113.695 161.250 113.985 161.295 ;
        RECT 115.585 161.250 115.875 161.295 ;
        RECT 110.575 161.110 115.875 161.250 ;
        RECT 110.575 161.065 110.865 161.110 ;
        RECT 113.695 161.065 113.985 161.110 ;
        RECT 115.585 161.065 115.875 161.110 ;
        RECT 116.440 161.250 116.760 161.310 ;
        RECT 117.910 161.250 118.050 161.405 ;
        RECT 118.280 161.390 118.600 161.650 ;
        RECT 118.830 161.590 118.970 161.745 ;
        RECT 119.200 161.730 119.520 161.990 ;
        RECT 119.660 161.930 119.980 161.990 ;
        RECT 121.975 161.930 122.265 161.975 ;
        RECT 119.660 161.790 122.265 161.930 ;
        RECT 119.660 161.730 119.980 161.790 ;
        RECT 121.975 161.745 122.265 161.790 ;
        RECT 122.435 161.745 122.725 161.975 ;
        RECT 122.510 161.590 122.650 161.745 ;
        RECT 122.880 161.730 123.200 161.990 ;
        RECT 123.355 161.930 123.645 161.975 ;
        RECT 123.800 161.930 124.120 161.990 ;
        RECT 123.355 161.790 124.120 161.930 ;
        RECT 123.355 161.745 123.645 161.790 ;
        RECT 123.800 161.730 124.120 161.790 ;
        RECT 124.810 161.650 124.950 162.130 ;
        RECT 127.020 161.930 127.340 161.990 ;
        RECT 129.870 161.975 130.010 162.130 ;
        RECT 129.335 161.930 129.625 161.975 ;
        RECT 127.020 161.790 129.625 161.930 ;
        RECT 127.020 161.730 127.340 161.790 ;
        RECT 129.335 161.745 129.625 161.790 ;
        RECT 129.795 161.745 130.085 161.975 ;
        RECT 135.850 161.930 135.990 162.425 ;
        RECT 138.520 162.410 138.840 162.470 ;
        RECT 143.670 162.470 145.280 162.610 ;
        RECT 139.555 162.270 139.845 162.315 ;
        RECT 142.795 162.270 143.445 162.315 ;
        RECT 143.670 162.270 143.810 162.470 ;
        RECT 144.960 162.410 145.280 162.470 ;
        RECT 139.555 162.130 143.810 162.270 ;
        RECT 144.040 162.270 144.360 162.330 ;
        RECT 144.040 162.130 147.030 162.270 ;
        RECT 139.555 162.085 140.145 162.130 ;
        RECT 142.795 162.085 143.445 162.130 ;
        RECT 136.235 161.930 136.525 161.975 ;
        RECT 135.850 161.790 136.525 161.930 ;
        RECT 136.235 161.745 136.525 161.790 ;
        RECT 139.855 161.770 140.145 162.085 ;
        RECT 144.040 162.070 144.360 162.130 ;
        RECT 146.890 161.975 147.030 162.130 ;
        RECT 147.720 162.070 148.040 162.330 ;
        RECT 140.935 161.930 141.225 161.975 ;
        RECT 144.515 161.930 144.805 161.975 ;
        RECT 146.350 161.930 146.640 161.975 ;
        RECT 140.935 161.790 146.640 161.930 ;
        RECT 140.935 161.745 141.225 161.790 ;
        RECT 144.515 161.745 144.805 161.790 ;
        RECT 146.350 161.745 146.640 161.790 ;
        RECT 146.815 161.745 147.105 161.975 ;
        RECT 118.830 161.450 122.650 161.590 ;
        RECT 124.720 161.390 125.040 161.650 ;
        RECT 125.655 161.590 125.945 161.635 ;
        RECT 126.100 161.590 126.420 161.650 ;
        RECT 125.655 161.450 126.420 161.590 ;
        RECT 125.655 161.405 125.945 161.450 ;
        RECT 126.100 161.390 126.420 161.450 ;
        RECT 130.240 161.590 130.560 161.650 ;
        RECT 132.555 161.590 132.845 161.635 ;
        RECT 133.000 161.590 133.320 161.650 ;
        RECT 130.240 161.450 133.320 161.590 ;
        RECT 130.240 161.390 130.560 161.450 ;
        RECT 132.555 161.405 132.845 161.450 ;
        RECT 133.000 161.390 133.320 161.450 ;
        RECT 133.460 161.390 133.780 161.650 ;
        RECT 138.060 161.390 138.380 161.650 ;
        RECT 145.435 161.590 145.725 161.635 ;
        RECT 147.810 161.590 147.950 162.070 ;
        RECT 145.435 161.450 147.950 161.590 ;
        RECT 145.435 161.405 145.725 161.450 ;
        RECT 118.740 161.250 119.060 161.310 ;
        RECT 116.440 161.110 119.060 161.250 ;
        RECT 116.440 161.050 116.760 161.110 ;
        RECT 118.740 161.050 119.060 161.110 ;
        RECT 120.595 161.250 120.885 161.295 ;
        RECT 127.020 161.250 127.340 161.310 ;
        RECT 120.595 161.110 127.340 161.250 ;
        RECT 120.595 161.065 120.885 161.110 ;
        RECT 127.020 161.050 127.340 161.110 ;
        RECT 140.935 161.250 141.225 161.295 ;
        RECT 144.055 161.250 144.345 161.295 ;
        RECT 145.945 161.250 146.235 161.295 ;
        RECT 140.935 161.110 146.235 161.250 ;
        RECT 140.935 161.065 141.225 161.110 ;
        RECT 144.055 161.065 144.345 161.110 ;
        RECT 145.945 161.065 146.235 161.110 ;
        RECT 94.820 160.770 101.490 160.910 ;
        RECT 105.415 160.910 105.705 160.955 ;
        RECT 119.660 160.910 119.980 160.970 ;
        RECT 105.415 160.770 119.980 160.910 ;
        RECT 94.820 160.710 95.140 160.770 ;
        RECT 96.200 160.710 96.520 160.770 ;
        RECT 105.415 160.725 105.705 160.770 ;
        RECT 119.660 160.710 119.980 160.770 ;
        RECT 124.720 160.910 125.040 160.970 ;
        RECT 129.320 160.910 129.640 160.970 ;
        RECT 124.720 160.770 129.640 160.910 ;
        RECT 124.720 160.710 125.040 160.770 ;
        RECT 129.320 160.710 129.640 160.770 ;
        RECT 2.750 160.090 158.230 160.570 ;
        RECT 19.380 159.890 19.700 159.950 ;
        RECT 31.340 159.890 31.660 159.950 ;
        RECT 19.380 159.750 31.660 159.890 ;
        RECT 19.380 159.690 19.700 159.750 ;
        RECT 31.340 159.690 31.660 159.750 ;
        RECT 35.020 159.690 35.340 159.950 ;
        RECT 40.080 159.890 40.400 159.950 ;
        RECT 44.680 159.890 45.000 159.950 ;
        RECT 57.560 159.890 57.880 159.950 ;
        RECT 40.080 159.750 45.000 159.890 ;
        RECT 40.080 159.690 40.400 159.750 ;
        RECT 44.680 159.690 45.000 159.750 ;
        RECT 54.890 159.750 57.880 159.890 ;
        RECT 5.085 159.550 5.375 159.595 ;
        RECT 6.975 159.550 7.265 159.595 ;
        RECT 10.095 159.550 10.385 159.595 ;
        RECT 5.085 159.410 10.385 159.550 ;
        RECT 5.085 159.365 5.375 159.410 ;
        RECT 6.975 159.365 7.265 159.410 ;
        RECT 10.095 159.365 10.385 159.410 ;
        RECT 12.480 159.550 12.800 159.610 ;
        RECT 12.480 159.410 18.690 159.550 ;
        RECT 12.480 159.350 12.800 159.410 ;
        RECT 18.550 159.255 18.690 159.410 ;
        RECT 19.470 159.255 19.610 159.690 ;
        RECT 24.900 159.550 25.220 159.610 ;
        RECT 32.260 159.550 32.580 159.610 ;
        RECT 22.230 159.410 25.220 159.550 ;
        RECT 4.215 159.210 4.505 159.255 ;
        RECT 12.955 159.210 13.245 159.255 ;
        RECT 4.215 159.070 10.870 159.210 ;
        RECT 4.215 159.025 4.505 159.070 ;
        RECT 10.730 158.930 10.870 159.070 ;
        RECT 12.955 159.070 18.230 159.210 ;
        RECT 12.955 159.025 13.245 159.070 ;
        RECT 4.680 158.870 4.970 158.915 ;
        RECT 6.515 158.870 6.805 158.915 ;
        RECT 10.095 158.870 10.385 158.915 ;
        RECT 4.680 158.730 10.385 158.870 ;
        RECT 4.680 158.685 4.970 158.730 ;
        RECT 6.515 158.685 6.805 158.730 ;
        RECT 10.095 158.685 10.385 158.730 ;
        RECT 10.640 158.670 10.960 158.930 ;
        RECT 18.090 158.915 18.230 159.070 ;
        RECT 18.475 159.025 18.765 159.255 ;
        RECT 19.395 159.025 19.685 159.255 ;
        RECT 5.595 158.345 5.885 158.575 ;
        RECT 7.875 158.530 8.525 158.575 ;
        RECT 8.800 158.530 9.120 158.590 ;
        RECT 11.175 158.575 11.465 158.890 ;
        RECT 14.335 158.870 14.625 158.915 ;
        RECT 18.015 158.870 18.305 158.915 ;
        RECT 22.230 158.870 22.370 159.410 ;
        RECT 24.900 159.350 25.220 159.410 ;
        RECT 30.050 159.410 32.580 159.550 ;
        RECT 24.990 159.210 25.130 159.350 ;
        RECT 30.050 159.255 30.190 159.410 ;
        RECT 32.260 159.350 32.580 159.410 ;
        RECT 32.720 159.350 33.040 159.610 ;
        RECT 24.990 159.070 26.510 159.210 ;
        RECT 14.335 158.730 16.390 158.870 ;
        RECT 14.335 158.685 14.625 158.730 ;
        RECT 11.175 158.530 11.765 158.575 ;
        RECT 7.875 158.390 11.765 158.530 ;
        RECT 7.875 158.345 8.525 158.390 ;
        RECT 5.670 158.190 5.810 158.345 ;
        RECT 8.800 158.330 9.120 158.390 ;
        RECT 11.475 158.345 11.765 158.390 ;
        RECT 16.250 158.235 16.390 158.730 ;
        RECT 18.015 158.730 22.370 158.870 ;
        RECT 18.015 158.685 18.305 158.730 ;
        RECT 22.600 158.670 22.920 158.930 ;
        RECT 23.520 158.915 23.840 158.930 ;
        RECT 23.355 158.685 23.840 158.915 ;
        RECT 24.455 158.685 24.745 158.915 ;
        RECT 25.145 158.870 25.435 158.915 ;
        RECT 25.820 158.870 26.140 158.930 ;
        RECT 25.145 158.730 26.140 158.870 ;
        RECT 26.370 158.870 26.510 159.070 ;
        RECT 29.975 159.025 30.265 159.255 ;
        RECT 35.110 159.210 35.250 159.690 ;
        RECT 37.780 159.350 38.100 159.610 ;
        RECT 41.935 159.550 42.225 159.595 ;
        RECT 44.220 159.550 44.540 159.610 ;
        RECT 41.935 159.410 44.540 159.550 ;
        RECT 41.935 159.365 42.225 159.410 ;
        RECT 44.220 159.350 44.540 159.410 ;
        RECT 52.515 159.550 52.805 159.595 ;
        RECT 54.890 159.550 55.030 159.750 ;
        RECT 57.560 159.690 57.880 159.750 ;
        RECT 58.020 159.890 58.340 159.950 ;
        RECT 58.940 159.890 59.260 159.950 ;
        RECT 58.020 159.750 59.260 159.890 ;
        RECT 58.020 159.690 58.340 159.750 ;
        RECT 58.940 159.690 59.260 159.750 ;
        RECT 59.860 159.890 60.180 159.950 ;
        RECT 63.540 159.890 63.860 159.950 ;
        RECT 68.140 159.890 68.460 159.950 ;
        RECT 59.860 159.750 63.310 159.890 ;
        RECT 59.860 159.690 60.180 159.750 ;
        RECT 52.515 159.410 55.030 159.550 ;
        RECT 55.375 159.550 55.665 159.595 ;
        RECT 58.495 159.550 58.785 159.595 ;
        RECT 60.385 159.550 60.675 159.595 ;
        RECT 62.620 159.550 62.940 159.610 ;
        RECT 55.375 159.410 60.675 159.550 ;
        RECT 52.515 159.365 52.805 159.410 ;
        RECT 55.375 159.365 55.665 159.410 ;
        RECT 58.495 159.365 58.785 159.410 ;
        RECT 60.385 159.365 60.675 159.410 ;
        RECT 61.330 159.410 62.940 159.550 ;
        RECT 37.870 159.210 38.010 159.350 ;
        RECT 39.620 159.210 39.940 159.270 ;
        RECT 45.140 159.210 45.460 159.270 ;
        RECT 48.820 159.210 49.140 159.270 ;
        RECT 35.110 159.070 35.710 159.210 ;
        RECT 37.870 159.070 38.475 159.210 ;
        RECT 30.435 158.870 30.725 158.915 ;
        RECT 26.370 158.730 30.725 158.870 ;
        RECT 25.145 158.685 25.435 158.730 ;
        RECT 23.520 158.670 23.840 158.685 ;
        RECT 20.760 158.530 21.080 158.590 ;
        RECT 23.995 158.530 24.285 158.575 ;
        RECT 20.760 158.390 24.285 158.530 ;
        RECT 24.530 158.530 24.670 158.685 ;
        RECT 25.820 158.670 26.140 158.730 ;
        RECT 30.435 158.685 30.725 158.730 ;
        RECT 32.260 158.870 32.580 158.930 ;
        RECT 35.020 158.915 35.340 158.930 ;
        RECT 35.570 158.915 35.710 159.070 ;
        RECT 34.115 158.870 34.405 158.915 ;
        RECT 32.260 158.730 34.405 158.870 ;
        RECT 32.260 158.670 32.580 158.730 ;
        RECT 34.115 158.685 34.405 158.730 ;
        RECT 34.855 158.685 35.340 158.915 ;
        RECT 35.495 158.685 35.785 158.915 ;
        RECT 35.020 158.670 35.340 158.685 ;
        RECT 35.940 158.670 36.260 158.930 ;
        RECT 36.860 158.915 37.180 158.930 ;
        RECT 38.335 158.915 38.475 159.070 ;
        RECT 39.620 159.070 40.770 159.210 ;
        RECT 39.620 159.010 39.940 159.070 ;
        RECT 36.645 158.685 37.180 158.915 ;
        RECT 37.795 158.685 38.085 158.915 ;
        RECT 38.260 158.685 38.550 158.915 ;
        RECT 38.790 158.730 39.850 158.870 ;
        RECT 36.860 158.670 37.180 158.685 ;
        RECT 27.200 158.530 27.520 158.590 ;
        RECT 30.895 158.530 31.185 158.575 ;
        RECT 37.870 158.530 38.010 158.685 ;
        RECT 24.530 158.390 31.185 158.530 ;
        RECT 20.760 158.330 21.080 158.390 ;
        RECT 23.610 158.250 23.750 158.390 ;
        RECT 23.995 158.345 24.285 158.390 ;
        RECT 27.200 158.330 27.520 158.390 ;
        RECT 30.895 158.345 31.185 158.390 ;
        RECT 37.410 158.390 38.010 158.530 ;
        RECT 13.415 158.190 13.705 158.235 ;
        RECT 5.670 158.050 13.705 158.190 ;
        RECT 13.415 158.005 13.705 158.050 ;
        RECT 16.175 158.005 16.465 158.235 ;
        RECT 23.520 157.990 23.840 158.250 ;
        RECT 25.835 158.190 26.125 158.235 ;
        RECT 26.280 158.190 26.600 158.250 ;
        RECT 37.410 158.235 37.550 158.390 ;
        RECT 25.835 158.050 26.600 158.190 ;
        RECT 25.835 158.005 26.125 158.050 ;
        RECT 26.280 157.990 26.600 158.050 ;
        RECT 37.335 158.005 37.625 158.235 ;
        RECT 37.780 158.190 38.100 158.250 ;
        RECT 38.790 158.190 38.930 158.730 ;
        RECT 39.710 158.575 39.850 158.730 ;
        RECT 40.120 158.685 40.410 158.915 ;
        RECT 40.630 158.870 40.770 159.070 ;
        RECT 45.140 159.070 49.140 159.210 ;
        RECT 45.140 159.010 45.460 159.070 ;
        RECT 48.820 159.010 49.140 159.070 ;
        RECT 41.460 158.870 41.780 158.930 ;
        RECT 43.775 158.870 44.065 158.915 ;
        RECT 40.630 158.730 44.065 158.870 ;
        RECT 39.175 158.345 39.465 158.575 ;
        RECT 39.635 158.345 39.925 158.575 ;
        RECT 40.195 158.530 40.335 158.685 ;
        RECT 41.460 158.670 41.780 158.730 ;
        RECT 43.775 158.685 44.065 158.730 ;
        RECT 46.075 158.870 46.365 158.915 ;
        RECT 50.200 158.870 50.520 158.930 ;
        RECT 52.590 158.870 52.730 159.365 ;
        RECT 58.020 159.210 58.340 159.270 ;
        RECT 61.330 159.255 61.470 159.410 ;
        RECT 62.620 159.350 62.940 159.410 ;
        RECT 59.875 159.210 60.165 159.255 ;
        RECT 58.020 159.070 60.165 159.210 ;
        RECT 58.020 159.010 58.340 159.070 ;
        RECT 59.875 159.025 60.165 159.070 ;
        RECT 61.255 159.025 61.545 159.255 ;
        RECT 63.170 159.210 63.310 159.750 ;
        RECT 63.540 159.750 68.460 159.890 ;
        RECT 63.540 159.690 63.860 159.750 ;
        RECT 68.140 159.690 68.460 159.750 ;
        RECT 68.600 159.690 68.920 159.950 ;
        RECT 86.555 159.890 86.845 159.935 ;
        RECT 87.000 159.890 87.320 159.950 ;
        RECT 86.555 159.750 87.320 159.890 ;
        RECT 86.555 159.705 86.845 159.750 ;
        RECT 87.000 159.690 87.320 159.750 ;
        RECT 88.380 159.890 88.700 159.950 ;
        RECT 91.140 159.890 91.460 159.950 ;
        RECT 105.860 159.890 106.180 159.950 ;
        RECT 106.795 159.890 107.085 159.935 ;
        RECT 88.380 159.750 95.510 159.890 ;
        RECT 88.380 159.690 88.700 159.750 ;
        RECT 91.140 159.690 91.460 159.750 ;
        RECT 65.380 159.550 65.700 159.610 ;
        RECT 68.690 159.550 68.830 159.690 ;
        RECT 65.380 159.410 68.830 159.550 ;
        RECT 65.380 159.350 65.700 159.410 ;
        RECT 64.460 159.210 64.780 159.270 ;
        RECT 65.855 159.210 66.145 159.255 ;
        RECT 63.170 159.070 66.145 159.210 ;
        RECT 64.460 159.010 64.780 159.070 ;
        RECT 65.855 159.025 66.145 159.070 ;
        RECT 68.155 159.210 68.445 159.255 ;
        RECT 68.690 159.210 68.830 159.410 ;
        RECT 69.025 159.550 69.315 159.595 ;
        RECT 70.915 159.550 71.205 159.595 ;
        RECT 74.035 159.550 74.325 159.595 ;
        RECT 69.025 159.410 74.325 159.550 ;
        RECT 69.025 159.365 69.315 159.410 ;
        RECT 70.915 159.365 71.205 159.410 ;
        RECT 74.035 159.365 74.325 159.410 ;
        RECT 77.800 159.350 78.120 159.610 ;
        RECT 81.940 159.550 82.260 159.610 ;
        RECT 78.810 159.410 82.260 159.550 ;
        RECT 68.155 159.070 68.830 159.210 ;
        RECT 69.980 159.210 70.300 159.270 ;
        RECT 76.880 159.210 77.200 159.270 ;
        RECT 78.810 159.210 78.950 159.410 ;
        RECT 81.940 159.350 82.260 159.410 ;
        RECT 83.335 159.365 83.625 159.595 ;
        RECT 69.980 159.070 75.270 159.210 ;
        RECT 68.155 159.025 68.445 159.070 ;
        RECT 46.075 158.730 49.970 158.870 ;
        RECT 46.075 158.685 46.365 158.730 ;
        RECT 40.195 158.390 43.990 158.530 ;
        RECT 37.780 158.050 38.930 158.190 ;
        RECT 39.250 158.190 39.390 158.345 ;
        RECT 40.080 158.190 40.400 158.250 ;
        RECT 39.250 158.050 40.400 158.190 ;
        RECT 37.780 157.990 38.100 158.050 ;
        RECT 40.080 157.990 40.400 158.050 ;
        RECT 41.015 158.190 41.305 158.235 ;
        RECT 43.300 158.190 43.620 158.250 ;
        RECT 41.015 158.050 43.620 158.190 ;
        RECT 43.850 158.190 43.990 158.390 ;
        RECT 44.220 158.330 44.540 158.590 ;
        RECT 46.980 158.330 47.300 158.590 ;
        RECT 47.915 158.530 48.205 158.575 ;
        RECT 49.280 158.530 49.600 158.590 ;
        RECT 47.915 158.390 49.600 158.530 ;
        RECT 49.830 158.530 49.970 158.730 ;
        RECT 50.200 158.730 52.730 158.870 ;
        RECT 50.200 158.670 50.520 158.730 ;
        RECT 54.295 158.575 54.585 158.890 ;
        RECT 55.375 158.870 55.665 158.915 ;
        RECT 58.955 158.870 59.245 158.915 ;
        RECT 60.790 158.870 61.080 158.915 ;
        RECT 55.375 158.730 61.080 158.870 ;
        RECT 55.375 158.685 55.665 158.730 ;
        RECT 58.955 158.685 59.245 158.730 ;
        RECT 60.790 158.685 61.080 158.730 ;
        RECT 61.700 158.670 62.020 158.930 ;
        RECT 62.620 158.870 62.940 158.930 ;
        RECT 62.620 158.730 66.530 158.870 ;
        RECT 62.620 158.670 62.940 158.730 ;
        RECT 57.560 158.575 57.880 158.590 ;
        RECT 53.995 158.530 54.585 158.575 ;
        RECT 57.235 158.530 57.885 158.575 ;
        RECT 49.830 158.390 53.650 158.530 ;
        RECT 47.915 158.345 48.205 158.390 ;
        RECT 49.280 158.330 49.600 158.390 ;
        RECT 44.680 158.190 45.000 158.250 ;
        RECT 43.850 158.050 45.000 158.190 ;
        RECT 41.015 158.005 41.305 158.050 ;
        RECT 43.300 157.990 43.620 158.050 ;
        RECT 44.680 157.990 45.000 158.050 ;
        RECT 49.755 158.190 50.045 158.235 ;
        RECT 50.660 158.190 50.980 158.250 ;
        RECT 49.755 158.050 50.980 158.190 ;
        RECT 49.755 158.005 50.045 158.050 ;
        RECT 50.660 157.990 50.980 158.050 ;
        RECT 52.055 158.190 52.345 158.235 ;
        RECT 52.500 158.190 52.820 158.250 ;
        RECT 52.055 158.050 52.820 158.190 ;
        RECT 53.510 158.190 53.650 158.390 ;
        RECT 53.995 158.390 57.885 158.530 ;
        RECT 53.995 158.345 54.285 158.390 ;
        RECT 57.235 158.345 57.885 158.390 ;
        RECT 58.480 158.530 58.800 158.590 ;
        RECT 65.840 158.530 66.160 158.590 ;
        RECT 58.480 158.390 63.310 158.530 ;
        RECT 57.560 158.330 57.880 158.345 ;
        RECT 58.480 158.330 58.800 158.390 ;
        RECT 59.860 158.190 60.180 158.250 ;
        RECT 53.510 158.050 60.180 158.190 ;
        RECT 52.055 158.005 52.345 158.050 ;
        RECT 52.500 157.990 52.820 158.050 ;
        RECT 59.860 157.990 60.180 158.050 ;
        RECT 62.620 157.990 62.940 158.250 ;
        RECT 63.170 158.235 63.310 158.390 ;
        RECT 64.090 158.390 66.160 158.530 ;
        RECT 64.090 158.250 64.230 158.390 ;
        RECT 63.095 158.005 63.385 158.235 ;
        RECT 64.000 157.990 64.320 158.250 ;
        RECT 64.920 157.990 65.240 158.250 ;
        RECT 65.470 158.235 65.610 158.390 ;
        RECT 65.840 158.330 66.160 158.390 ;
        RECT 65.395 158.005 65.685 158.235 ;
        RECT 66.390 158.190 66.530 158.730 ;
        RECT 68.230 158.530 68.370 159.025 ;
        RECT 69.980 159.010 70.300 159.070 ;
        RECT 68.620 158.870 68.910 158.915 ;
        RECT 70.455 158.870 70.745 158.915 ;
        RECT 74.035 158.870 74.325 158.915 ;
        RECT 75.130 158.890 75.270 159.070 ;
        RECT 76.880 159.070 78.950 159.210 ;
        RECT 79.180 159.210 79.500 159.270 ;
        RECT 79.655 159.210 79.945 159.255 ;
        RECT 79.180 159.070 79.945 159.210 ;
        RECT 83.410 159.210 83.550 159.365 ;
        RECT 83.780 159.350 84.100 159.610 ;
        RECT 86.095 159.550 86.385 159.595 ;
        RECT 86.095 159.410 90.450 159.550 ;
        RECT 86.095 159.365 86.385 159.410 ;
        RECT 84.255 159.210 84.545 159.255 ;
        RECT 87.920 159.210 88.240 159.270 ;
        RECT 83.410 159.070 88.240 159.210 ;
        RECT 76.880 159.010 77.200 159.070 ;
        RECT 79.180 159.010 79.500 159.070 ;
        RECT 79.655 159.025 79.945 159.070 ;
        RECT 84.255 159.025 84.545 159.070 ;
        RECT 87.920 159.010 88.240 159.070 ;
        RECT 68.620 158.730 74.325 158.870 ;
        RECT 68.620 158.685 68.910 158.730 ;
        RECT 70.455 158.685 70.745 158.730 ;
        RECT 74.035 158.685 74.325 158.730 ;
        RECT 75.115 158.870 75.405 158.890 ;
        RECT 77.340 158.870 77.660 158.930 ;
        RECT 82.860 158.870 83.180 158.930 ;
        RECT 75.115 158.730 83.180 158.870 ;
        RECT 69.060 158.530 69.380 158.590 ;
        RECT 75.115 158.575 75.405 158.730 ;
        RECT 77.340 158.670 77.660 158.730 ;
        RECT 82.860 158.670 83.180 158.730 ;
        RECT 87.000 158.670 87.320 158.930 ;
        RECT 88.380 158.670 88.700 158.930 ;
        RECT 90.310 158.915 90.450 159.410 ;
        RECT 95.370 159.210 95.510 159.750 ;
        RECT 105.860 159.750 107.085 159.890 ;
        RECT 105.860 159.690 106.180 159.750 ;
        RECT 106.795 159.705 107.085 159.750 ;
        RECT 108.620 159.690 108.940 159.950 ;
        RECT 116.900 159.890 117.220 159.950 ;
        RECT 150.940 159.890 151.260 159.950 ;
        RECT 116.900 159.750 151.260 159.890 ;
        RECT 116.900 159.690 117.220 159.750 ;
        RECT 150.940 159.690 151.260 159.750 ;
        RECT 98.005 159.550 98.295 159.595 ;
        RECT 99.895 159.550 100.185 159.595 ;
        RECT 103.015 159.550 103.305 159.595 ;
        RECT 98.005 159.410 103.305 159.550 ;
        RECT 98.005 159.365 98.295 159.410 ;
        RECT 99.895 159.365 100.185 159.410 ;
        RECT 103.015 159.365 103.305 159.410 ;
        RECT 104.940 159.550 105.260 159.610 ;
        RECT 109.080 159.550 109.400 159.610 ;
        RECT 117.360 159.550 117.680 159.610 ;
        RECT 104.940 159.410 117.680 159.550 ;
        RECT 104.940 159.350 105.260 159.410 ;
        RECT 109.080 159.350 109.400 159.410 ;
        RECT 117.360 159.350 117.680 159.410 ;
        RECT 117.820 159.550 118.140 159.610 ;
        RECT 124.720 159.550 125.040 159.610 ;
        RECT 129.795 159.550 130.085 159.595 ;
        RECT 117.820 159.410 122.650 159.550 ;
        RECT 117.820 159.350 118.140 159.410 ;
        RECT 95.370 159.070 121.270 159.210 ;
        RECT 90.235 158.870 90.525 158.915 ;
        RECT 92.980 158.870 93.300 158.930 ;
        RECT 95.370 158.915 95.510 159.070 ;
        RECT 90.235 158.730 93.300 158.870 ;
        RECT 90.235 158.685 90.525 158.730 ;
        RECT 92.980 158.670 93.300 158.730 ;
        RECT 94.375 158.685 94.665 158.915 ;
        RECT 95.295 158.685 95.585 158.915 ;
        RECT 68.230 158.390 69.380 158.530 ;
        RECT 69.060 158.330 69.380 158.390 ;
        RECT 69.535 158.345 69.825 158.575 ;
        RECT 71.815 158.530 72.465 158.575 ;
        RECT 75.115 158.530 75.705 158.575 ;
        RECT 71.815 158.390 75.705 158.530 ;
        RECT 71.815 158.345 72.465 158.390 ;
        RECT 75.415 158.345 75.705 158.390 ;
        RECT 80.575 158.530 80.865 158.575 ;
        RECT 81.480 158.530 81.800 158.590 ;
        RECT 80.575 158.390 81.800 158.530 ;
        RECT 80.575 158.345 80.865 158.390 ;
        RECT 69.610 158.190 69.750 158.345 ;
        RECT 81.480 158.330 81.800 158.390 ;
        RECT 81.940 158.530 82.260 158.590 ;
        RECT 94.450 158.530 94.590 158.685 ;
        RECT 95.740 158.670 96.060 158.930 ;
        RECT 96.200 158.870 96.520 158.930 ;
        RECT 106.410 158.915 106.550 159.070 ;
        RECT 97.135 158.870 97.425 158.915 ;
        RECT 96.200 158.730 97.425 158.870 ;
        RECT 96.200 158.670 96.520 158.730 ;
        RECT 97.135 158.685 97.425 158.730 ;
        RECT 97.600 158.870 97.890 158.915 ;
        RECT 99.435 158.870 99.725 158.915 ;
        RECT 103.015 158.870 103.305 158.915 ;
        RECT 97.600 158.730 103.305 158.870 ;
        RECT 97.600 158.685 97.890 158.730 ;
        RECT 99.435 158.685 99.725 158.730 ;
        RECT 103.015 158.685 103.305 158.730 ;
        RECT 98.040 158.530 98.360 158.590 ;
        RECT 81.940 158.390 94.130 158.530 ;
        RECT 94.450 158.390 98.360 158.530 ;
        RECT 81.940 158.330 82.260 158.390 ;
        RECT 66.390 158.050 69.750 158.190 ;
        RECT 76.880 157.990 77.200 158.250 ;
        RECT 80.115 158.190 80.405 158.235 ;
        RECT 82.860 158.190 83.180 158.250 ;
        RECT 86.540 158.190 86.860 158.250 ;
        RECT 80.115 158.050 86.860 158.190 ;
        RECT 80.115 158.005 80.405 158.050 ;
        RECT 82.860 157.990 83.180 158.050 ;
        RECT 86.540 157.990 86.860 158.050 ;
        RECT 87.935 158.190 88.225 158.235 ;
        RECT 88.840 158.190 89.160 158.250 ;
        RECT 87.935 158.050 89.160 158.190 ;
        RECT 87.935 158.005 88.225 158.050 ;
        RECT 88.840 157.990 89.160 158.050 ;
        RECT 89.300 157.990 89.620 158.250 ;
        RECT 92.520 158.190 92.840 158.250 ;
        RECT 93.455 158.190 93.745 158.235 ;
        RECT 92.520 158.050 93.745 158.190 ;
        RECT 93.990 158.190 94.130 158.390 ;
        RECT 98.040 158.330 98.360 158.390 ;
        RECT 98.515 158.530 98.805 158.575 ;
        RECT 99.880 158.530 100.200 158.590 ;
        RECT 104.095 158.575 104.385 158.890 ;
        RECT 106.335 158.685 106.625 158.915 ;
        RECT 109.540 158.670 109.860 158.930 ;
        RECT 116.900 158.870 117.220 158.930 ;
        RECT 110.090 158.730 117.220 158.870 ;
        RECT 110.090 158.590 110.230 158.730 ;
        RECT 116.900 158.670 117.220 158.730 ;
        RECT 120.580 158.870 120.900 158.930 ;
        RECT 121.130 158.915 121.270 159.070 ;
        RECT 121.960 159.010 122.280 159.270 ;
        RECT 122.510 159.210 122.650 159.410 ;
        RECT 124.720 159.410 130.085 159.550 ;
        RECT 124.720 159.350 125.040 159.410 ;
        RECT 129.795 159.365 130.085 159.410 ;
        RECT 135.315 159.210 135.605 159.255 ;
        RECT 140.375 159.210 140.665 159.255 ;
        RECT 140.820 159.210 141.140 159.270 ;
        RECT 122.510 159.070 130.930 159.210 ;
        RECT 121.055 158.870 121.345 158.915 ;
        RECT 120.580 158.730 121.345 158.870 ;
        RECT 120.580 158.670 120.900 158.730 ;
        RECT 121.055 158.685 121.345 158.730 ;
        RECT 121.500 158.870 121.820 158.930 ;
        RECT 123.355 158.870 123.645 158.915 ;
        RECT 121.500 158.730 123.645 158.870 ;
        RECT 121.500 158.670 121.820 158.730 ;
        RECT 123.355 158.685 123.645 158.730 ;
        RECT 128.400 158.670 128.720 158.930 ;
        RECT 130.790 158.915 130.930 159.070 ;
        RECT 131.250 159.070 141.140 159.210 ;
        RECT 130.715 158.685 131.005 158.915 ;
        RECT 98.515 158.390 100.200 158.530 ;
        RECT 98.515 158.345 98.805 158.390 ;
        RECT 99.880 158.330 100.200 158.390 ;
        RECT 100.795 158.530 101.445 158.575 ;
        RECT 104.095 158.530 104.685 158.575 ;
        RECT 104.940 158.530 105.260 158.590 ;
        RECT 110.000 158.530 110.320 158.590 ;
        RECT 124.735 158.530 125.025 158.575 ;
        RECT 125.640 158.530 125.960 158.590 ;
        RECT 100.795 158.390 110.320 158.530 ;
        RECT 100.795 158.345 101.445 158.390 ;
        RECT 104.395 158.345 104.685 158.390 ;
        RECT 104.940 158.330 105.260 158.390 ;
        RECT 110.000 158.330 110.320 158.390 ;
        RECT 112.390 158.390 121.730 158.530 ;
        RECT 96.660 158.190 96.980 158.250 ;
        RECT 102.640 158.190 102.960 158.250 ;
        RECT 93.990 158.050 102.960 158.190 ;
        RECT 92.520 157.990 92.840 158.050 ;
        RECT 93.455 158.005 93.745 158.050 ;
        RECT 96.660 157.990 96.980 158.050 ;
        RECT 102.640 157.990 102.960 158.050 ;
        RECT 103.100 158.190 103.420 158.250 ;
        RECT 108.620 158.190 108.940 158.250 ;
        RECT 112.390 158.190 112.530 158.390 ;
        RECT 103.100 158.050 112.530 158.190 ;
        RECT 112.760 158.190 113.080 158.250 ;
        RECT 115.995 158.190 116.285 158.235 ;
        RECT 112.760 158.050 116.285 158.190 ;
        RECT 103.100 157.990 103.420 158.050 ;
        RECT 108.620 157.990 108.940 158.050 ;
        RECT 112.760 157.990 113.080 158.050 ;
        RECT 115.995 158.005 116.285 158.050 ;
        RECT 116.440 158.190 116.760 158.250 ;
        RECT 121.590 158.235 121.730 158.390 ;
        RECT 124.735 158.390 125.960 158.530 ;
        RECT 124.735 158.345 125.025 158.390 ;
        RECT 125.640 158.330 125.960 158.390 ;
        RECT 126.115 158.530 126.405 158.575 ;
        RECT 126.560 158.530 126.880 158.590 ;
        RECT 126.115 158.390 126.880 158.530 ;
        RECT 126.115 158.345 126.405 158.390 ;
        RECT 126.560 158.330 126.880 158.390 ;
        RECT 127.020 158.330 127.340 158.590 ;
        RECT 128.875 158.530 129.165 158.575 ;
        RECT 127.570 158.390 129.165 158.530 ;
        RECT 119.215 158.190 119.505 158.235 ;
        RECT 116.440 158.050 119.505 158.190 ;
        RECT 116.440 157.990 116.760 158.050 ;
        RECT 119.215 158.005 119.505 158.050 ;
        RECT 121.515 158.005 121.805 158.235 ;
        RECT 121.960 158.190 122.280 158.250 ;
        RECT 127.570 158.190 127.710 158.390 ;
        RECT 128.875 158.345 129.165 158.390 ;
        RECT 129.320 158.530 129.640 158.590 ;
        RECT 131.250 158.530 131.390 159.070 ;
        RECT 135.315 159.025 135.605 159.070 ;
        RECT 140.375 159.025 140.665 159.070 ;
        RECT 140.820 159.010 141.140 159.070 ;
        RECT 144.500 159.010 144.820 159.270 ;
        RECT 133.460 158.870 133.780 158.930 ;
        RECT 139.455 158.870 139.745 158.915 ;
        RECT 144.590 158.870 144.730 159.010 ;
        RECT 133.460 158.730 144.730 158.870 ;
        RECT 133.460 158.670 133.780 158.730 ;
        RECT 139.455 158.685 139.745 158.730 ;
        RECT 135.760 158.530 136.080 158.590 ;
        RECT 129.320 158.390 131.390 158.530 ;
        RECT 131.710 158.390 136.080 158.530 ;
        RECT 129.320 158.330 129.640 158.390 ;
        RECT 131.710 158.250 131.850 158.390 ;
        RECT 121.960 158.050 127.710 158.190 ;
        RECT 127.955 158.190 128.245 158.235 ;
        RECT 130.240 158.190 130.560 158.250 ;
        RECT 127.955 158.050 130.560 158.190 ;
        RECT 121.960 157.990 122.280 158.050 ;
        RECT 127.955 158.005 128.245 158.050 ;
        RECT 130.240 157.990 130.560 158.050 ;
        RECT 131.620 157.990 131.940 158.250 ;
        RECT 132.080 157.990 132.400 158.250 ;
        RECT 133.920 157.990 134.240 158.250 ;
        RECT 134.470 158.235 134.610 158.390 ;
        RECT 135.760 158.330 136.080 158.390 ;
        RECT 134.395 158.005 134.685 158.235 ;
        RECT 137.155 158.190 137.445 158.235 ;
        RECT 137.600 158.190 137.920 158.250 ;
        RECT 137.155 158.050 137.920 158.190 ;
        RECT 137.155 158.005 137.445 158.050 ;
        RECT 137.600 157.990 137.920 158.050 ;
        RECT 138.980 158.190 139.300 158.250 ;
        RECT 141.740 158.190 142.060 158.250 ;
        RECT 138.980 158.050 142.060 158.190 ;
        RECT 138.980 157.990 139.300 158.050 ;
        RECT 141.740 157.990 142.060 158.050 ;
        RECT 2.750 157.370 159.030 157.850 ;
        RECT 7.895 157.170 8.185 157.215 ;
        RECT 10.180 157.170 10.500 157.230 ;
        RECT 12.940 157.170 13.260 157.230 ;
        RECT 22.600 157.170 22.920 157.230 ;
        RECT 23.535 157.170 23.825 157.215 ;
        RECT 27.660 157.170 27.980 157.230 ;
        RECT 7.895 157.030 13.260 157.170 ;
        RECT 7.895 156.985 8.185 157.030 ;
        RECT 10.180 156.970 10.500 157.030 ;
        RECT 12.940 156.970 13.260 157.030 ;
        RECT 13.720 157.030 19.610 157.170 ;
        RECT 13.720 156.830 13.860 157.030 ;
        RECT 19.470 156.890 19.610 157.030 ;
        RECT 22.600 157.030 23.825 157.170 ;
        RECT 22.600 156.970 22.920 157.030 ;
        RECT 23.535 156.985 23.825 157.030 ;
        RECT 24.070 157.030 27.980 157.170 ;
        RECT 7.510 156.690 13.860 156.830 ;
        RECT 14.315 156.830 14.965 156.875 ;
        RECT 17.915 156.830 18.205 156.875 ;
        RECT 14.315 156.690 18.205 156.830 ;
        RECT 7.510 156.195 7.650 156.690 ;
        RECT 14.315 156.645 14.965 156.690 ;
        RECT 17.615 156.645 18.205 156.690 ;
        RECT 17.615 156.550 17.905 156.645 ;
        RECT 19.380 156.630 19.700 156.890 ;
        RECT 8.355 156.305 8.645 156.535 ;
        RECT 7.435 155.965 7.725 156.195 ;
        RECT 8.430 156.150 8.570 156.305 ;
        RECT 10.640 156.290 10.960 156.550 ;
        RECT 11.120 156.490 11.410 156.535 ;
        RECT 12.955 156.490 13.245 156.535 ;
        RECT 16.535 156.490 16.825 156.535 ;
        RECT 11.120 156.350 16.825 156.490 ;
        RECT 11.120 156.305 11.410 156.350 ;
        RECT 12.955 156.305 13.245 156.350 ;
        RECT 16.535 156.305 16.825 156.350 ;
        RECT 17.540 156.490 17.905 156.550 ;
        RECT 24.070 156.490 24.210 157.030 ;
        RECT 27.660 156.970 27.980 157.030 ;
        RECT 29.055 156.985 29.345 157.215 ;
        RECT 24.530 156.690 26.970 156.830 ;
        RECT 24.530 156.535 24.670 156.690 ;
        RECT 17.540 156.350 24.210 156.490 ;
        RECT 17.540 156.330 17.905 156.350 ;
        RECT 17.540 156.290 17.860 156.330 ;
        RECT 24.455 156.305 24.745 156.535 ;
        RECT 8.430 156.010 10.870 156.150 ;
        RECT 10.180 155.270 10.500 155.530 ;
        RECT 10.730 155.470 10.870 156.010 ;
        RECT 12.020 155.950 12.340 156.210 ;
        RECT 19.395 156.150 19.685 156.195 ;
        RECT 20.760 156.150 21.080 156.210 ;
        RECT 22.615 156.150 22.905 156.195 ;
        RECT 19.395 156.010 22.905 156.150 ;
        RECT 19.395 155.965 19.685 156.010 ;
        RECT 20.760 155.950 21.080 156.010 ;
        RECT 22.615 155.965 22.905 156.010 ;
        RECT 23.980 156.150 24.300 156.210 ;
        RECT 24.530 156.150 24.670 156.305 ;
        RECT 24.900 156.290 25.220 156.550 ;
        RECT 25.375 156.305 25.665 156.535 ;
        RECT 25.820 156.490 26.140 156.550 ;
        RECT 26.295 156.490 26.585 156.535 ;
        RECT 25.820 156.350 26.585 156.490 ;
        RECT 25.450 156.150 25.590 156.305 ;
        RECT 25.820 156.290 26.140 156.350 ;
        RECT 26.295 156.305 26.585 156.350 ;
        RECT 23.980 156.010 24.670 156.150 ;
        RECT 24.990 156.010 25.590 156.150 ;
        RECT 26.830 156.150 26.970 156.690 ;
        RECT 27.675 156.490 27.965 156.535 ;
        RECT 29.130 156.490 29.270 156.985 ;
        RECT 38.240 156.970 38.560 157.230 ;
        RECT 42.380 157.170 42.700 157.230 ;
        RECT 46.120 157.170 46.410 157.215 ;
        RECT 42.380 157.030 46.410 157.170 ;
        RECT 42.380 156.970 42.700 157.030 ;
        RECT 46.120 156.985 46.410 157.030 ;
        RECT 30.895 156.830 31.185 156.875 ;
        RECT 31.800 156.830 32.120 156.890 ;
        RECT 38.330 156.830 38.470 156.970 ;
        RECT 38.715 156.830 39.005 156.875 ;
        RECT 30.895 156.690 32.120 156.830 ;
        RECT 30.895 156.645 31.185 156.690 ;
        RECT 27.675 156.350 29.270 156.490 ;
        RECT 27.675 156.305 27.965 156.350 ;
        RECT 28.120 156.150 28.440 156.210 ;
        RECT 26.830 156.010 28.440 156.150 ;
        RECT 23.980 155.950 24.300 156.010 ;
        RECT 11.525 155.810 11.815 155.855 ;
        RECT 13.415 155.810 13.705 155.855 ;
        RECT 16.535 155.810 16.825 155.855 ;
        RECT 11.525 155.670 16.825 155.810 ;
        RECT 11.525 155.625 11.815 155.670 ;
        RECT 13.415 155.625 13.705 155.670 ;
        RECT 16.535 155.625 16.825 155.670 ;
        RECT 18.000 155.810 18.320 155.870 ;
        RECT 24.070 155.810 24.210 155.950 ;
        RECT 18.000 155.670 24.210 155.810 ;
        RECT 24.990 155.810 25.130 156.010 ;
        RECT 28.120 155.950 28.440 156.010 ;
        RECT 30.970 155.810 31.110 156.645 ;
        RECT 31.800 156.630 32.120 156.690 ;
        RECT 34.190 156.690 39.005 156.830 ;
        RECT 32.260 156.490 32.580 156.550 ;
        RECT 34.190 156.535 34.330 156.690 ;
        RECT 38.715 156.645 39.005 156.690 ;
        RECT 41.935 156.830 42.225 156.875 ;
        RECT 42.840 156.830 43.160 156.890 ;
        RECT 41.935 156.690 43.160 156.830 ;
        RECT 41.935 156.645 42.225 156.690 ;
        RECT 42.840 156.630 43.160 156.690 ;
        RECT 43.775 156.830 44.065 156.875 ;
        RECT 45.140 156.830 45.460 156.890 ;
        RECT 43.775 156.690 45.460 156.830 ;
        RECT 46.195 156.830 46.335 156.985 ;
        RECT 47.900 156.970 48.220 157.230 ;
        RECT 52.500 157.170 52.820 157.230 ;
        RECT 48.450 157.030 52.820 157.170 ;
        RECT 48.450 156.830 48.590 157.030 ;
        RECT 52.500 156.970 52.820 157.030 ;
        RECT 53.880 157.170 54.200 157.230 ;
        RECT 55.275 157.170 55.565 157.215 ;
        RECT 53.880 157.030 55.565 157.170 ;
        RECT 53.880 156.970 54.200 157.030 ;
        RECT 55.275 156.985 55.565 157.030 ;
        RECT 56.180 156.970 56.500 157.230 ;
        RECT 61.700 156.970 62.020 157.230 ;
        RECT 63.540 156.970 63.860 157.230 ;
        RECT 81.940 157.170 82.260 157.230 ;
        RECT 64.090 157.030 78.030 157.170 ;
        RECT 51.120 156.830 51.440 156.890 ;
        RECT 53.435 156.830 53.725 156.875 ;
        RECT 57.115 156.830 57.405 156.875 ;
        RECT 64.090 156.830 64.230 157.030 ;
        RECT 77.890 156.890 78.030 157.030 ;
        RECT 78.350 157.030 82.260 157.170 ;
        RECT 46.195 156.690 48.590 156.830 ;
        RECT 49.375 156.690 64.230 156.830 ;
        RECT 69.515 156.830 70.165 156.875 ;
        RECT 70.440 156.830 70.760 156.890 ;
        RECT 73.115 156.830 73.405 156.875 ;
        RECT 69.515 156.690 73.405 156.830 ;
        RECT 43.775 156.645 44.065 156.690 ;
        RECT 45.140 156.630 45.460 156.690 ;
        RECT 35.020 156.535 35.340 156.550 ;
        RECT 36.400 156.535 36.720 156.550 ;
        RECT 34.115 156.490 34.405 156.535 ;
        RECT 32.260 156.350 34.405 156.490 ;
        RECT 32.260 156.290 32.580 156.350 ;
        RECT 34.115 156.305 34.405 156.350 ;
        RECT 34.855 156.305 35.340 156.535 ;
        RECT 35.495 156.305 35.785 156.535 ;
        RECT 35.955 156.305 36.245 156.535 ;
        RECT 36.400 156.490 36.730 156.535 ;
        RECT 37.320 156.490 37.640 156.550 ;
        RECT 38.240 156.490 38.560 156.550 ;
        RECT 44.235 156.490 44.525 156.535 ;
        RECT 49.375 156.490 49.515 156.690 ;
        RECT 51.120 156.630 51.440 156.690 ;
        RECT 53.435 156.645 53.725 156.690 ;
        RECT 57.115 156.645 57.405 156.690 ;
        RECT 69.515 156.645 70.165 156.690 ;
        RECT 70.440 156.630 70.760 156.690 ;
        RECT 72.815 156.645 73.405 156.690 ;
        RECT 36.400 156.350 36.915 156.490 ;
        RECT 37.320 156.480 47.210 156.490 ;
        RECT 47.530 156.480 49.515 156.490 ;
        RECT 37.320 156.350 49.515 156.480 ;
        RECT 50.675 156.490 50.965 156.535 ;
        RECT 51.580 156.490 51.900 156.550 ;
        RECT 55.720 156.490 56.040 156.550 ;
        RECT 50.675 156.350 56.040 156.490 ;
        RECT 36.400 156.305 36.730 156.350 ;
        RECT 35.020 156.290 35.340 156.305 ;
        RECT 31.340 155.950 31.660 156.210 ;
        RECT 31.800 155.950 32.120 156.210 ;
        RECT 35.570 155.870 35.710 156.305 ;
        RECT 36.030 156.150 36.170 156.305 ;
        RECT 36.400 156.290 36.720 156.305 ;
        RECT 37.320 156.290 37.640 156.350 ;
        RECT 38.240 156.290 38.560 156.350 ;
        RECT 44.235 156.305 44.525 156.350 ;
        RECT 47.070 156.340 47.670 156.350 ;
        RECT 50.675 156.305 50.965 156.350 ;
        RECT 51.580 156.290 51.900 156.350 ;
        RECT 55.720 156.290 56.040 156.350 ;
        RECT 58.495 156.490 58.785 156.535 ;
        RECT 59.860 156.490 60.180 156.550 ;
        RECT 58.495 156.350 60.180 156.490 ;
        RECT 58.495 156.305 58.785 156.350 ;
        RECT 59.860 156.290 60.180 156.350 ;
        RECT 60.320 156.290 60.640 156.550 ;
        RECT 61.240 156.490 61.560 156.550 ;
        RECT 64.015 156.490 64.305 156.535 ;
        RECT 64.920 156.490 65.240 156.550 ;
        RECT 61.240 156.350 65.240 156.490 ;
        RECT 61.240 156.290 61.560 156.350 ;
        RECT 64.015 156.305 64.305 156.350 ;
        RECT 64.920 156.290 65.240 156.350 ;
        RECT 65.380 156.490 65.700 156.550 ;
        RECT 65.855 156.490 66.145 156.535 ;
        RECT 65.380 156.350 66.145 156.490 ;
        RECT 65.380 156.290 65.700 156.350 ;
        RECT 65.855 156.305 66.145 156.350 ;
        RECT 66.320 156.490 66.610 156.535 ;
        RECT 68.155 156.490 68.445 156.535 ;
        RECT 71.735 156.490 72.025 156.535 ;
        RECT 66.320 156.350 72.025 156.490 ;
        RECT 66.320 156.305 66.610 156.350 ;
        RECT 68.155 156.305 68.445 156.350 ;
        RECT 71.735 156.305 72.025 156.350 ;
        RECT 72.815 156.330 73.105 156.645 ;
        RECT 77.800 156.630 78.120 156.890 ;
        RECT 49.280 156.150 49.600 156.210 ;
        RECT 55.260 156.150 55.580 156.210 ;
        RECT 36.030 156.010 49.120 156.150 ;
        RECT 34.100 155.810 34.420 155.870 ;
        RECT 24.990 155.670 30.650 155.810 ;
        RECT 30.970 155.670 34.420 155.810 ;
        RECT 18.000 155.610 18.320 155.670 ;
        RECT 24.990 155.530 25.130 155.670 ;
        RECT 15.700 155.470 16.020 155.530 ;
        RECT 10.730 155.330 16.020 155.470 ;
        RECT 15.700 155.270 16.020 155.330 ;
        RECT 19.840 155.270 20.160 155.530 ;
        RECT 23.060 155.470 23.380 155.530 ;
        RECT 23.980 155.470 24.300 155.530 ;
        RECT 23.060 155.330 24.300 155.470 ;
        RECT 23.060 155.270 23.380 155.330 ;
        RECT 23.980 155.270 24.300 155.330 ;
        RECT 24.900 155.270 25.220 155.530 ;
        RECT 25.820 155.470 26.140 155.530 ;
        RECT 26.755 155.470 27.045 155.515 ;
        RECT 25.820 155.330 27.045 155.470 ;
        RECT 30.510 155.470 30.650 155.670 ;
        RECT 34.100 155.610 34.420 155.670 ;
        RECT 35.480 155.610 35.800 155.870 ;
        RECT 40.080 155.810 40.400 155.870 ;
        RECT 36.950 155.670 40.400 155.810 ;
        RECT 36.950 155.470 37.090 155.670 ;
        RECT 40.080 155.610 40.400 155.670 ;
        RECT 40.540 155.810 40.860 155.870 ;
        RECT 42.840 155.810 43.160 155.870 ;
        RECT 43.760 155.810 44.080 155.870 ;
        RECT 40.540 155.670 44.080 155.810 ;
        RECT 40.540 155.610 40.860 155.670 ;
        RECT 42.840 155.610 43.160 155.670 ;
        RECT 43.760 155.610 44.080 155.670 ;
        RECT 44.680 155.810 45.000 155.870 ;
        RECT 46.995 155.810 47.285 155.855 ;
        RECT 44.680 155.670 47.285 155.810 ;
        RECT 48.980 155.810 49.120 156.010 ;
        RECT 49.280 156.010 55.580 156.150 ;
        RECT 49.280 155.950 49.600 156.010 ;
        RECT 55.260 155.950 55.580 156.010 ;
        RECT 64.460 155.950 64.780 156.210 ;
        RECT 67.220 155.950 67.540 156.210 ;
        RECT 67.680 156.150 68.000 156.210 ;
        RECT 69.520 156.150 69.840 156.210 ;
        RECT 74.595 156.150 74.885 156.195 ;
        RECT 67.680 156.010 74.885 156.150 ;
        RECT 67.680 155.950 68.000 156.010 ;
        RECT 69.520 155.950 69.840 156.010 ;
        RECT 74.595 155.965 74.885 156.010 ;
        RECT 76.880 156.150 77.200 156.210 ;
        RECT 78.350 156.195 78.490 157.030 ;
        RECT 81.940 156.970 82.260 157.030 ;
        RECT 88.840 157.170 89.160 157.230 ;
        RECT 88.840 157.030 90.450 157.170 ;
        RECT 88.840 156.970 89.160 157.030 ;
        RECT 78.735 156.830 79.025 156.875 ;
        RECT 84.355 156.830 84.645 156.875 ;
        RECT 85.160 156.830 85.480 156.890 ;
        RECT 90.310 156.875 90.450 157.030 ;
        RECT 92.610 157.030 96.660 157.170 ;
        RECT 87.595 156.830 88.245 156.875 ;
        RECT 78.735 156.690 81.250 156.830 ;
        RECT 78.735 156.645 79.025 156.690 ;
        RECT 81.110 156.535 81.250 156.690 ;
        RECT 84.355 156.690 88.245 156.830 ;
        RECT 84.355 156.645 84.945 156.690 ;
        RECT 81.035 156.305 81.325 156.535 ;
        RECT 81.480 156.490 81.800 156.550 ;
        RECT 81.480 156.350 83.550 156.490 ;
        RECT 78.275 156.150 78.565 156.195 ;
        RECT 76.880 156.010 78.565 156.150 ;
        RECT 76.880 155.950 77.200 156.010 ;
        RECT 78.275 155.965 78.565 156.010 ;
        RECT 79.195 155.965 79.485 156.195 ;
        RECT 81.110 156.150 81.250 156.305 ;
        RECT 81.480 156.290 81.800 156.350 ;
        RECT 82.875 156.150 83.165 156.195 ;
        RECT 81.110 156.010 83.165 156.150 ;
        RECT 82.875 155.965 83.165 156.010 ;
        RECT 83.410 156.150 83.550 156.350 ;
        RECT 84.655 156.330 84.945 156.645 ;
        RECT 85.160 156.630 85.480 156.690 ;
        RECT 87.595 156.645 88.245 156.690 ;
        RECT 90.235 156.645 90.525 156.875 ;
        RECT 85.735 156.490 86.025 156.535 ;
        RECT 89.315 156.490 89.605 156.535 ;
        RECT 91.150 156.490 91.440 156.535 ;
        RECT 85.735 156.350 91.440 156.490 ;
        RECT 85.735 156.305 86.025 156.350 ;
        RECT 89.315 156.305 89.605 156.350 ;
        RECT 91.150 156.305 91.440 156.350 ;
        RECT 91.615 156.490 91.905 156.535 ;
        RECT 92.060 156.490 92.380 156.550 ;
        RECT 92.610 156.535 92.750 157.030 ;
        RECT 96.520 156.830 96.660 157.030 ;
        RECT 99.435 156.985 99.725 157.215 ;
        RECT 96.520 156.690 99.190 156.830 ;
        RECT 91.615 156.350 92.380 156.490 ;
        RECT 91.615 156.305 91.905 156.350 ;
        RECT 92.060 156.290 92.380 156.350 ;
        RECT 92.535 156.305 92.825 156.535 ;
        RECT 97.595 156.490 97.885 156.535 ;
        RECT 93.990 156.350 97.885 156.490 ;
        RECT 92.610 156.150 92.750 156.305 ;
        RECT 83.410 156.010 92.750 156.150 ;
        RECT 92.980 156.150 93.300 156.210 ;
        RECT 93.990 156.195 94.130 156.350 ;
        RECT 97.595 156.305 97.885 156.350 ;
        RECT 93.915 156.150 94.205 156.195 ;
        RECT 92.980 156.010 94.205 156.150 ;
        RECT 63.540 155.810 63.860 155.870 ;
        RECT 48.980 155.670 63.860 155.810 ;
        RECT 64.550 155.810 64.690 155.950 ;
        RECT 65.380 155.810 65.700 155.870 ;
        RECT 64.550 155.670 65.700 155.810 ;
        RECT 44.680 155.610 45.000 155.670 ;
        RECT 46.995 155.625 47.285 155.670 ;
        RECT 63.540 155.610 63.860 155.670 ;
        RECT 65.380 155.610 65.700 155.670 ;
        RECT 66.725 155.810 67.015 155.855 ;
        RECT 68.615 155.810 68.905 155.855 ;
        RECT 71.735 155.810 72.025 155.855 ;
        RECT 66.725 155.670 72.025 155.810 ;
        RECT 79.270 155.810 79.410 155.965 ;
        RECT 83.410 155.810 83.550 156.010 ;
        RECT 92.980 155.950 93.300 156.010 ;
        RECT 93.915 155.965 94.205 156.010 ;
        RECT 96.200 155.950 96.520 156.210 ;
        RECT 96.675 155.965 96.965 156.195 ;
        RECT 97.135 156.150 97.425 156.195 ;
        RECT 98.500 156.150 98.820 156.210 ;
        RECT 97.135 156.010 98.820 156.150 ;
        RECT 99.050 156.150 99.190 156.690 ;
        RECT 99.510 156.490 99.650 156.985 ;
        RECT 99.880 156.970 100.200 157.230 ;
        RECT 101.260 157.170 101.580 157.230 ;
        RECT 102.655 157.170 102.945 157.215 ;
        RECT 106.335 157.170 106.625 157.215 ;
        RECT 101.260 157.030 102.945 157.170 ;
        RECT 101.260 156.970 101.580 157.030 ;
        RECT 102.655 156.985 102.945 157.030 ;
        RECT 103.650 157.030 106.625 157.170 ;
        RECT 100.815 156.490 101.105 156.535 ;
        RECT 99.510 156.350 101.105 156.490 ;
        RECT 100.815 156.305 101.105 156.350 ;
        RECT 101.735 156.490 102.025 156.535 ;
        RECT 103.650 156.490 103.790 157.030 ;
        RECT 106.335 156.985 106.625 157.030 ;
        RECT 106.780 157.170 107.100 157.230 ;
        RECT 108.175 157.170 108.465 157.215 ;
        RECT 106.780 157.030 108.465 157.170 ;
        RECT 106.780 156.970 107.100 157.030 ;
        RECT 108.175 156.985 108.465 157.030 ;
        RECT 108.620 156.970 108.940 157.230 ;
        RECT 120.580 157.170 120.900 157.230 ;
        RECT 122.895 157.170 123.185 157.215 ;
        RECT 120.580 157.030 123.185 157.170 ;
        RECT 120.580 156.970 120.900 157.030 ;
        RECT 122.895 156.985 123.185 157.030 ;
        RECT 127.955 157.170 128.245 157.215 ;
        RECT 129.780 157.170 130.100 157.230 ;
        RECT 127.955 157.030 130.100 157.170 ;
        RECT 127.955 156.985 128.245 157.030 ;
        RECT 129.780 156.970 130.100 157.030 ;
        RECT 132.080 156.970 132.400 157.230 ;
        RECT 141.740 157.170 142.060 157.230 ;
        RECT 150.495 157.170 150.785 157.215 ;
        RECT 141.740 157.030 150.785 157.170 ;
        RECT 141.740 156.970 142.060 157.030 ;
        RECT 150.495 156.985 150.785 157.030 ;
        RECT 104.955 156.830 105.245 156.875 ;
        RECT 105.860 156.830 106.180 156.890 ;
        RECT 104.955 156.690 106.180 156.830 ;
        RECT 104.955 156.645 105.245 156.690 ;
        RECT 105.860 156.630 106.180 156.690 ;
        RECT 112.760 156.830 113.080 156.890 ;
        RECT 112.760 156.690 114.370 156.830 ;
        RECT 112.760 156.630 113.080 156.690 ;
        RECT 111.395 156.490 111.685 156.535 ;
        RECT 111.840 156.490 112.160 156.550 ;
        RECT 101.735 156.350 103.790 156.490 ;
        RECT 104.110 156.350 112.160 156.490 ;
        RECT 101.735 156.305 102.025 156.350 ;
        RECT 103.575 156.150 103.865 156.195 ;
        RECT 104.110 156.150 104.250 156.350 ;
        RECT 111.395 156.305 111.685 156.350 ;
        RECT 111.840 156.290 112.160 156.350 ;
        RECT 112.315 156.490 112.605 156.535 ;
        RECT 113.680 156.490 114.000 156.550 ;
        RECT 114.230 156.535 114.370 156.690 ;
        RECT 115.520 156.630 115.840 156.890 ;
        RECT 117.815 156.830 118.465 156.875 ;
        RECT 121.415 156.830 121.705 156.875 ;
        RECT 122.420 156.830 122.740 156.890 ;
        RECT 117.815 156.690 122.740 156.830 ;
        RECT 117.815 156.645 118.465 156.690 ;
        RECT 121.115 156.645 121.705 156.690 ;
        RECT 112.315 156.350 114.000 156.490 ;
        RECT 112.315 156.305 112.605 156.350 ;
        RECT 113.680 156.290 114.000 156.350 ;
        RECT 114.155 156.305 114.445 156.535 ;
        RECT 114.620 156.490 114.910 156.535 ;
        RECT 116.455 156.490 116.745 156.535 ;
        RECT 120.035 156.490 120.325 156.535 ;
        RECT 114.620 156.350 120.325 156.490 ;
        RECT 114.620 156.305 114.910 156.350 ;
        RECT 116.455 156.305 116.745 156.350 ;
        RECT 120.035 156.305 120.325 156.350 ;
        RECT 121.115 156.330 121.405 156.645 ;
        RECT 122.420 156.630 122.740 156.690 ;
        RECT 124.260 156.830 124.580 156.890 ;
        RECT 127.495 156.830 127.785 156.875 ;
        RECT 124.260 156.690 130.010 156.830 ;
        RECT 124.260 156.630 124.580 156.690 ;
        RECT 127.495 156.645 127.785 156.690 ;
        RECT 125.195 156.490 125.485 156.535 ;
        RECT 125.195 156.350 125.870 156.490 ;
        RECT 125.195 156.305 125.485 156.350 ;
        RECT 99.050 156.010 104.250 156.150 ;
        RECT 97.135 155.965 97.425 156.010 ;
        RECT 79.270 155.670 83.550 155.810 ;
        RECT 85.735 155.810 86.025 155.855 ;
        RECT 88.855 155.810 89.145 155.855 ;
        RECT 90.745 155.810 91.035 155.855 ;
        RECT 85.735 155.670 91.035 155.810 ;
        RECT 66.725 155.625 67.015 155.670 ;
        RECT 68.615 155.625 68.905 155.670 ;
        RECT 71.735 155.625 72.025 155.670 ;
        RECT 85.735 155.625 86.025 155.670 ;
        RECT 88.855 155.625 89.145 155.670 ;
        RECT 90.745 155.625 91.035 155.670 ;
        RECT 92.060 155.810 92.380 155.870 ;
        RECT 93.440 155.810 93.760 155.870 ;
        RECT 96.290 155.810 96.430 155.950 ;
        RECT 92.060 155.670 96.430 155.810 ;
        RECT 96.750 155.810 96.890 155.965 ;
        RECT 98.500 155.950 98.820 156.010 ;
        RECT 103.575 155.965 103.865 156.010 ;
        RECT 109.080 155.950 109.400 156.210 ;
        RECT 110.920 156.150 111.240 156.210 ;
        RECT 118.740 156.150 119.060 156.210 ;
        RECT 110.920 156.010 119.060 156.150 ;
        RECT 110.920 155.950 111.240 156.010 ;
        RECT 113.770 155.855 113.910 156.010 ;
        RECT 118.740 155.950 119.060 156.010 ;
        RECT 125.730 155.855 125.870 156.350 ;
        RECT 129.320 156.290 129.640 156.550 ;
        RECT 128.875 156.150 129.165 156.195 ;
        RECT 129.410 156.150 129.550 156.290 ;
        RECT 128.875 156.010 129.550 156.150 ;
        RECT 129.870 156.150 130.010 156.690 ;
        RECT 130.255 156.490 130.545 156.535 ;
        RECT 132.170 156.490 132.310 156.970 ;
        RECT 137.140 156.875 137.460 156.890 ;
        RECT 145.420 156.875 145.740 156.890 ;
        RECT 134.035 156.830 134.325 156.875 ;
        RECT 137.140 156.830 137.925 156.875 ;
        RECT 134.035 156.690 137.925 156.830 ;
        RECT 134.035 156.645 134.625 156.690 ;
        RECT 130.255 156.350 132.310 156.490 ;
        RECT 130.255 156.305 130.545 156.350 ;
        RECT 134.335 156.330 134.625 156.645 ;
        RECT 137.140 156.645 137.925 156.690 ;
        RECT 145.415 156.830 146.065 156.875 ;
        RECT 149.015 156.830 149.305 156.875 ;
        RECT 145.415 156.690 149.305 156.830 ;
        RECT 145.415 156.645 146.065 156.690 ;
        RECT 148.715 156.645 149.305 156.690 ;
        RECT 137.140 156.630 137.460 156.645 ;
        RECT 145.420 156.630 145.740 156.645 ;
        RECT 135.415 156.490 135.705 156.535 ;
        RECT 138.995 156.490 139.285 156.535 ;
        RECT 140.830 156.490 141.120 156.535 ;
        RECT 135.415 156.350 141.120 156.490 ;
        RECT 135.415 156.305 135.705 156.350 ;
        RECT 138.995 156.305 139.285 156.350 ;
        RECT 140.830 156.305 141.120 156.350 ;
        RECT 142.220 156.490 142.510 156.535 ;
        RECT 144.055 156.490 144.345 156.535 ;
        RECT 147.635 156.490 147.925 156.535 ;
        RECT 142.220 156.350 147.925 156.490 ;
        RECT 142.220 156.305 142.510 156.350 ;
        RECT 144.055 156.305 144.345 156.350 ;
        RECT 147.635 156.305 147.925 156.350 ;
        RECT 148.715 156.330 149.005 156.645 ;
        RECT 130.700 156.150 131.020 156.210 ;
        RECT 139.915 156.150 140.205 156.195 ;
        RECT 141.295 156.150 141.585 156.195 ;
        RECT 141.755 156.150 142.045 156.195 ;
        RECT 129.870 156.010 131.020 156.150 ;
        RECT 128.875 155.965 129.165 156.010 ;
        RECT 130.700 155.950 131.020 156.010 ;
        RECT 131.250 156.010 140.205 156.150 ;
        RECT 131.250 155.855 131.390 156.010 ;
        RECT 139.915 155.965 140.205 156.010 ;
        RECT 140.910 156.010 142.045 156.150 ;
        RECT 96.750 155.670 97.350 155.810 ;
        RECT 92.060 155.610 92.380 155.670 ;
        RECT 93.440 155.610 93.760 155.670 ;
        RECT 30.510 155.330 37.090 155.470 ;
        RECT 25.820 155.270 26.140 155.330 ;
        RECT 26.755 155.285 27.045 155.330 ;
        RECT 37.320 155.270 37.640 155.530 ;
        RECT 41.920 155.470 42.240 155.530 ;
        RECT 46.075 155.470 46.365 155.515 ;
        RECT 47.440 155.470 47.760 155.530 ;
        RECT 41.920 155.330 47.760 155.470 ;
        RECT 41.920 155.270 42.240 155.330 ;
        RECT 46.075 155.285 46.365 155.330 ;
        RECT 47.440 155.270 47.760 155.330 ;
        RECT 48.360 155.470 48.680 155.530 ;
        RECT 48.835 155.470 49.125 155.515 ;
        RECT 48.360 155.330 49.125 155.470 ;
        RECT 48.360 155.270 48.680 155.330 ;
        RECT 48.835 155.285 49.125 155.330 ;
        RECT 49.740 155.470 50.060 155.530 ;
        RECT 51.595 155.470 51.885 155.515 ;
        RECT 49.740 155.330 51.885 155.470 ;
        RECT 49.740 155.270 50.060 155.330 ;
        RECT 51.595 155.285 51.885 155.330 ;
        RECT 52.515 155.470 52.805 155.515 ;
        RECT 53.420 155.470 53.740 155.530 ;
        RECT 56.195 155.470 56.485 155.515 ;
        RECT 56.640 155.470 56.960 155.530 ;
        RECT 76.435 155.470 76.725 155.515 ;
        RECT 52.515 155.330 76.725 155.470 ;
        RECT 52.515 155.285 52.805 155.330 ;
        RECT 53.420 155.270 53.740 155.330 ;
        RECT 56.195 155.285 56.485 155.330 ;
        RECT 56.640 155.270 56.960 155.330 ;
        RECT 76.435 155.285 76.725 155.330 ;
        RECT 81.940 155.470 82.260 155.530 ;
        RECT 83.780 155.470 84.100 155.530 ;
        RECT 81.940 155.330 84.100 155.470 ;
        RECT 81.940 155.270 82.260 155.330 ;
        RECT 83.780 155.270 84.100 155.330 ;
        RECT 84.240 155.470 84.560 155.530 ;
        RECT 97.210 155.470 97.350 155.670 ;
        RECT 113.695 155.625 113.985 155.855 ;
        RECT 115.025 155.810 115.315 155.855 ;
        RECT 116.915 155.810 117.205 155.855 ;
        RECT 120.035 155.810 120.325 155.855 ;
        RECT 115.025 155.670 120.325 155.810 ;
        RECT 115.025 155.625 115.315 155.670 ;
        RECT 116.915 155.625 117.205 155.670 ;
        RECT 120.035 155.625 120.325 155.670 ;
        RECT 123.890 155.670 124.950 155.810 ;
        RECT 123.890 155.530 124.030 155.670 ;
        RECT 103.560 155.470 103.880 155.530 ;
        RECT 84.240 155.330 103.880 155.470 ;
        RECT 84.240 155.270 84.560 155.330 ;
        RECT 103.560 155.270 103.880 155.330 ;
        RECT 123.800 155.270 124.120 155.530 ;
        RECT 124.260 155.270 124.580 155.530 ;
        RECT 124.810 155.470 124.950 155.670 ;
        RECT 125.655 155.625 125.945 155.855 ;
        RECT 131.175 155.625 131.465 155.855 ;
        RECT 133.000 155.810 133.320 155.870 ;
        RECT 135.415 155.810 135.705 155.855 ;
        RECT 138.535 155.810 138.825 155.855 ;
        RECT 140.425 155.810 140.715 155.855 ;
        RECT 133.000 155.670 135.070 155.810 ;
        RECT 133.000 155.610 133.320 155.670 ;
        RECT 132.555 155.470 132.845 155.515 ;
        RECT 133.920 155.470 134.240 155.530 ;
        RECT 124.810 155.330 134.240 155.470 ;
        RECT 134.930 155.470 135.070 155.670 ;
        RECT 135.415 155.670 140.715 155.810 ;
        RECT 135.415 155.625 135.705 155.670 ;
        RECT 138.535 155.625 138.825 155.670 ;
        RECT 140.425 155.625 140.715 155.670 ;
        RECT 140.910 155.470 141.050 156.010 ;
        RECT 141.295 155.965 141.585 156.010 ;
        RECT 141.755 155.965 142.045 156.010 ;
        RECT 143.120 155.950 143.440 156.210 ;
        RECT 142.625 155.810 142.915 155.855 ;
        RECT 144.515 155.810 144.805 155.855 ;
        RECT 147.635 155.810 147.925 155.855 ;
        RECT 142.625 155.670 147.925 155.810 ;
        RECT 142.625 155.625 142.915 155.670 ;
        RECT 144.515 155.625 144.805 155.670 ;
        RECT 147.635 155.625 147.925 155.670 ;
        RECT 134.930 155.330 141.050 155.470 ;
        RECT 132.555 155.285 132.845 155.330 ;
        RECT 133.920 155.270 134.240 155.330 ;
        RECT 2.750 154.650 158.230 155.130 ;
        RECT 12.020 154.450 12.340 154.510 ;
        RECT 13.415 154.450 13.705 154.495 ;
        RECT 12.020 154.310 13.705 154.450 ;
        RECT 12.020 154.250 12.340 154.310 ;
        RECT 13.415 154.265 13.705 154.310 ;
        RECT 15.790 154.310 18.230 154.450 ;
        RECT 5.085 154.110 5.375 154.155 ;
        RECT 6.975 154.110 7.265 154.155 ;
        RECT 10.095 154.110 10.385 154.155 ;
        RECT 5.085 153.970 10.385 154.110 ;
        RECT 5.085 153.925 5.375 153.970 ;
        RECT 6.975 153.925 7.265 153.970 ;
        RECT 10.095 153.925 10.385 153.970 ;
        RECT 12.480 154.110 12.800 154.170 ;
        RECT 15.790 154.110 15.930 154.310 ;
        RECT 12.480 153.970 15.930 154.110 ;
        RECT 12.480 153.910 12.800 153.970 ;
        RECT 16.175 153.925 16.465 154.155 ;
        RECT 4.200 153.230 4.520 153.490 ;
        RECT 4.680 153.430 4.970 153.475 ;
        RECT 6.515 153.430 6.805 153.475 ;
        RECT 10.095 153.430 10.385 153.475 ;
        RECT 4.680 153.290 10.385 153.430 ;
        RECT 4.680 153.245 4.970 153.290 ;
        RECT 6.515 153.245 6.805 153.290 ;
        RECT 10.095 153.245 10.385 153.290 ;
        RECT 5.595 153.090 5.885 153.135 ;
        RECT 6.040 153.090 6.360 153.150 ;
        RECT 11.175 153.135 11.465 153.450 ;
        RECT 14.335 153.430 14.625 153.475 ;
        RECT 16.250 153.430 16.390 153.925 ;
        RECT 18.090 153.475 18.230 154.310 ;
        RECT 19.840 154.250 20.160 154.510 ;
        RECT 20.760 154.250 21.080 154.510 ;
        RECT 21.220 154.450 21.540 154.510 ;
        RECT 24.440 154.450 24.760 154.510 ;
        RECT 21.220 154.310 24.760 154.450 ;
        RECT 21.220 154.250 21.540 154.310 ;
        RECT 24.440 154.250 24.760 154.310 ;
        RECT 25.310 154.450 25.600 154.495 ;
        RECT 25.820 154.450 26.140 154.510 ;
        RECT 25.310 154.310 26.140 154.450 ;
        RECT 25.310 154.265 25.600 154.310 ;
        RECT 25.820 154.250 26.140 154.310 ;
        RECT 31.340 154.450 31.660 154.510 ;
        RECT 33.195 154.450 33.485 154.495 ;
        RECT 31.340 154.310 33.485 154.450 ;
        RECT 31.340 154.250 31.660 154.310 ;
        RECT 33.195 154.265 33.485 154.310 ;
        RECT 34.100 154.450 34.420 154.510 ;
        RECT 35.480 154.450 35.800 154.510 ;
        RECT 34.100 154.310 35.800 154.450 ;
        RECT 34.100 154.250 34.420 154.310 ;
        RECT 35.480 154.250 35.800 154.310 ;
        RECT 37.780 154.250 38.100 154.510 ;
        RECT 38.715 154.265 39.005 154.495 ;
        RECT 39.635 154.450 39.925 154.495 ;
        RECT 40.080 154.450 40.400 154.510 ;
        RECT 39.635 154.310 40.400 154.450 ;
        RECT 39.635 154.265 39.925 154.310 ;
        RECT 19.930 154.110 20.070 154.250 ;
        RECT 18.550 153.970 20.070 154.110 ;
        RECT 18.550 153.815 18.690 153.970 ;
        RECT 18.475 153.585 18.765 153.815 ;
        RECT 19.380 153.570 19.700 153.830 ;
        RECT 14.335 153.290 16.390 153.430 ;
        RECT 14.335 153.245 14.625 153.290 ;
        RECT 18.015 153.245 18.305 153.475 ;
        RECT 20.315 153.245 20.605 153.475 ;
        RECT 20.850 153.430 20.990 154.250 ;
        RECT 24.865 154.110 25.155 154.155 ;
        RECT 26.755 154.110 27.045 154.155 ;
        RECT 29.875 154.110 30.165 154.155 ;
        RECT 24.865 153.970 30.165 154.110 ;
        RECT 24.865 153.925 25.155 153.970 ;
        RECT 26.755 153.925 27.045 153.970 ;
        RECT 29.875 153.925 30.165 153.970 ;
        RECT 32.735 154.110 33.025 154.155 ;
        RECT 32.735 153.970 36.630 154.110 ;
        RECT 32.735 153.925 33.025 153.970 ;
        RECT 36.490 153.815 36.630 153.970 ;
        RECT 23.995 153.770 24.285 153.815 ;
        RECT 36.415 153.770 36.705 153.815 ;
        RECT 37.870 153.770 38.010 154.250 ;
        RECT 38.790 154.110 38.930 154.265 ;
        RECT 40.080 154.250 40.400 154.310 ;
        RECT 41.920 154.250 42.240 154.510 ;
        RECT 43.315 154.450 43.605 154.495 ;
        RECT 45.140 154.450 45.460 154.510 ;
        RECT 43.315 154.310 45.460 154.450 ;
        RECT 43.315 154.265 43.605 154.310 ;
        RECT 45.140 154.250 45.460 154.310 ;
        RECT 46.520 154.250 46.840 154.510 ;
        RECT 49.280 154.250 49.600 154.510 ;
        RECT 51.120 154.450 51.440 154.510 ;
        RECT 49.830 154.310 51.440 154.450 ;
        RECT 42.010 154.110 42.150 154.250 ;
        RECT 38.790 153.970 42.150 154.110 ;
        RECT 42.395 153.925 42.685 154.155 ;
        RECT 49.830 154.110 49.970 154.310 ;
        RECT 51.120 154.250 51.440 154.310 ;
        RECT 51.580 154.250 51.900 154.510 ;
        RECT 56.640 154.450 56.960 154.510 ;
        RECT 55.810 154.310 56.960 154.450 ;
        RECT 51.670 154.110 51.810 154.250 ;
        RECT 53.420 154.110 53.740 154.170 ;
        RECT 45.230 153.970 49.970 154.110 ;
        RECT 50.290 153.970 51.810 154.110 ;
        RECT 52.130 153.970 53.740 154.110 ;
        RECT 23.995 153.630 34.790 153.770 ;
        RECT 23.995 153.585 24.285 153.630 ;
        RECT 34.650 153.490 34.790 153.630 ;
        RECT 36.415 153.630 38.010 153.770 ;
        RECT 41.920 153.770 42.240 153.830 ;
        RECT 42.470 153.770 42.610 153.925 ;
        RECT 41.920 153.630 42.610 153.770 ;
        RECT 43.300 153.770 43.620 153.830 ;
        RECT 43.300 153.630 43.990 153.770 ;
        RECT 36.415 153.585 36.705 153.630 ;
        RECT 41.920 153.570 42.240 153.630 ;
        RECT 43.300 153.570 43.620 153.630 ;
        RECT 21.695 153.430 21.985 153.475 ;
        RECT 20.850 153.290 21.985 153.430 ;
        RECT 21.695 153.245 21.985 153.290 ;
        RECT 22.155 153.245 22.445 153.475 ;
        RECT 24.460 153.430 24.750 153.475 ;
        RECT 26.295 153.430 26.585 153.475 ;
        RECT 29.875 153.430 30.165 153.475 ;
        RECT 24.460 153.290 30.165 153.430 ;
        RECT 24.460 153.245 24.750 153.290 ;
        RECT 26.295 153.245 26.585 153.290 ;
        RECT 29.875 153.245 30.165 153.290 ;
        RECT 5.595 152.950 6.360 153.090 ;
        RECT 5.595 152.905 5.885 152.950 ;
        RECT 6.040 152.890 6.360 152.950 ;
        RECT 7.875 153.090 8.525 153.135 ;
        RECT 11.175 153.090 11.765 153.135 ;
        RECT 14.780 153.090 15.100 153.150 ;
        RECT 7.875 152.950 15.100 153.090 ;
        RECT 7.875 152.905 8.525 152.950 ;
        RECT 11.475 152.905 11.765 152.950 ;
        RECT 14.780 152.890 15.100 152.950 ;
        RECT 15.240 153.090 15.560 153.150 ;
        RECT 20.390 153.090 20.530 153.245 ;
        RECT 15.240 152.950 20.530 153.090 ;
        RECT 15.240 152.890 15.560 152.950 ;
        RECT 21.220 152.890 21.540 153.150 ;
        RECT 22.230 153.090 22.370 153.245 ;
        RECT 23.520 153.090 23.840 153.150 ;
        RECT 27.660 153.135 27.980 153.150 ;
        RECT 30.955 153.135 31.245 153.450 ;
        RECT 34.560 153.230 34.880 153.490 ;
        RECT 36.875 153.430 37.165 153.475 ;
        RECT 38.240 153.430 38.560 153.490 ;
        RECT 36.875 153.290 38.560 153.430 ;
        RECT 36.875 153.245 37.165 153.290 ;
        RECT 38.240 153.230 38.560 153.290 ;
        RECT 22.230 152.950 23.840 153.090 ;
        RECT 12.955 152.750 13.245 152.795 ;
        RECT 15.700 152.750 16.020 152.810 ;
        RECT 12.955 152.610 16.020 152.750 ;
        RECT 12.955 152.565 13.245 152.610 ;
        RECT 15.700 152.550 16.020 152.610 ;
        RECT 17.080 152.750 17.400 152.810 ;
        RECT 22.230 152.750 22.370 152.950 ;
        RECT 23.520 152.890 23.840 152.950 ;
        RECT 27.655 153.090 28.305 153.135 ;
        RECT 30.955 153.090 31.545 153.135 ;
        RECT 27.655 152.950 31.545 153.090 ;
        RECT 27.655 152.905 28.305 152.950 ;
        RECT 31.255 152.905 31.545 152.950 ;
        RECT 35.020 153.090 35.340 153.150 ;
        RECT 38.945 153.090 39.235 153.135 ;
        RECT 41.920 153.090 42.240 153.150 ;
        RECT 35.020 152.950 42.240 153.090 ;
        RECT 27.660 152.890 27.980 152.905 ;
        RECT 35.020 152.890 35.340 152.950 ;
        RECT 38.945 152.905 39.235 152.950 ;
        RECT 41.920 152.890 42.240 152.950 ;
        RECT 17.080 152.610 22.370 152.750 ;
        RECT 17.080 152.550 17.400 152.610 ;
        RECT 23.060 152.550 23.380 152.810 ;
        RECT 25.820 152.750 26.140 152.810 ;
        RECT 26.740 152.750 27.060 152.810 ;
        RECT 33.640 152.750 33.960 152.810 ;
        RECT 25.820 152.610 33.960 152.750 ;
        RECT 25.820 152.550 26.140 152.610 ;
        RECT 26.740 152.550 27.060 152.610 ;
        RECT 33.640 152.550 33.960 152.610 ;
        RECT 38.240 152.750 38.560 152.810 ;
        RECT 42.380 152.750 42.700 152.810 ;
        RECT 43.270 152.750 43.560 152.795 ;
        RECT 38.240 152.610 43.560 152.750 ;
        RECT 43.850 152.750 43.990 153.630 ;
        RECT 45.230 153.475 45.370 153.970 ;
        RECT 48.375 153.770 48.665 153.815 ;
        RECT 50.290 153.770 50.430 153.970 ;
        RECT 52.130 153.770 52.270 153.970 ;
        RECT 53.420 153.910 53.740 153.970 ;
        RECT 54.355 154.110 54.645 154.155 ;
        RECT 55.810 154.110 55.950 154.310 ;
        RECT 56.640 154.250 56.960 154.310 ;
        RECT 57.560 154.450 57.880 154.510 ;
        RECT 61.700 154.450 62.020 154.510 ;
        RECT 57.560 154.310 62.020 154.450 ;
        RECT 57.560 154.250 57.880 154.310 ;
        RECT 61.700 154.250 62.020 154.310 ;
        RECT 65.855 154.450 66.145 154.495 ;
        RECT 66.300 154.450 66.620 154.510 ;
        RECT 65.855 154.310 66.620 154.450 ;
        RECT 65.855 154.265 66.145 154.310 ;
        RECT 66.300 154.250 66.620 154.310 ;
        RECT 66.775 154.450 67.065 154.495 ;
        RECT 75.500 154.450 75.820 154.510 ;
        RECT 78.275 154.450 78.565 154.495 ;
        RECT 66.775 154.310 75.270 154.450 ;
        RECT 66.775 154.265 67.065 154.310 ;
        RECT 54.355 153.970 55.950 154.110 ;
        RECT 56.145 154.110 56.435 154.155 ;
        RECT 58.035 154.110 58.325 154.155 ;
        RECT 61.155 154.110 61.445 154.155 ;
        RECT 67.220 154.110 67.540 154.170 ;
        RECT 56.145 153.970 61.445 154.110 ;
        RECT 54.355 153.925 54.645 153.970 ;
        RECT 56.145 153.925 56.435 153.970 ;
        RECT 58.035 153.925 58.325 153.970 ;
        RECT 61.155 153.925 61.445 153.970 ;
        RECT 61.790 153.970 67.540 154.110 ;
        RECT 48.375 153.630 50.430 153.770 ;
        RECT 50.750 153.630 52.270 153.770 ;
        RECT 52.500 153.770 52.820 153.830 ;
        RECT 55.275 153.770 55.565 153.815 ;
        RECT 59.860 153.770 60.180 153.830 ;
        RECT 52.500 153.630 55.030 153.770 ;
        RECT 48.375 153.585 48.665 153.630 ;
        RECT 45.155 153.245 45.445 153.475 ;
        RECT 45.615 153.430 45.905 153.475 ;
        RECT 47.900 153.430 48.220 153.490 ;
        RECT 45.615 153.290 48.220 153.430 ;
        RECT 45.615 153.245 45.905 153.290 ;
        RECT 47.900 153.230 48.220 153.290 ;
        RECT 48.820 153.430 49.140 153.490 ;
        RECT 49.740 153.430 50.060 153.490 ;
        RECT 50.750 153.430 50.890 153.630 ;
        RECT 52.500 153.570 52.820 153.630 ;
        RECT 54.890 153.475 55.030 153.630 ;
        RECT 55.275 153.630 60.180 153.770 ;
        RECT 55.275 153.585 55.565 153.630 ;
        RECT 59.860 153.570 60.180 153.630 ;
        RECT 60.320 153.770 60.640 153.830 ;
        RECT 61.790 153.770 61.930 153.970 ;
        RECT 67.220 153.910 67.540 153.970 ;
        RECT 60.320 153.630 61.930 153.770 ;
        RECT 60.320 153.570 60.640 153.630 ;
        RECT 64.920 153.570 65.240 153.830 ;
        RECT 65.380 153.770 65.700 153.830 ;
        RECT 70.455 153.770 70.745 153.815 ;
        RECT 65.380 153.630 70.745 153.770 ;
        RECT 65.380 153.570 65.700 153.630 ;
        RECT 70.455 153.585 70.745 153.630 ;
        RECT 53.435 153.430 53.725 153.475 ;
        RECT 48.820 153.290 50.890 153.430 ;
        RECT 51.670 153.290 53.725 153.430 ;
        RECT 48.820 153.230 49.140 153.290 ;
        RECT 49.740 153.230 50.060 153.290 ;
        RECT 51.670 153.150 51.810 153.290 ;
        RECT 53.435 153.245 53.725 153.290 ;
        RECT 54.815 153.245 55.105 153.475 ;
        RECT 55.740 153.430 56.030 153.475 ;
        RECT 57.575 153.430 57.865 153.475 ;
        RECT 61.155 153.430 61.445 153.475 ;
        RECT 55.740 153.290 61.445 153.430 ;
        RECT 55.740 153.245 56.030 153.290 ;
        RECT 57.575 153.245 57.865 153.290 ;
        RECT 61.155 153.245 61.445 153.290 ;
        RECT 51.135 152.905 51.425 153.135 ;
        RECT 51.580 153.090 51.900 153.150 ;
        RECT 52.500 153.090 52.820 153.150 ;
        RECT 51.580 152.950 52.820 153.090 ;
        RECT 46.520 152.750 46.840 152.810 ;
        RECT 43.850 152.610 46.840 152.750 ;
        RECT 38.240 152.550 38.560 152.610 ;
        RECT 42.380 152.550 42.700 152.610 ;
        RECT 43.270 152.565 43.560 152.610 ;
        RECT 46.520 152.550 46.840 152.610 ;
        RECT 46.980 152.550 47.300 152.810 ;
        RECT 50.660 152.750 50.980 152.810 ;
        RECT 51.210 152.750 51.350 152.905 ;
        RECT 51.580 152.890 51.900 152.950 ;
        RECT 52.500 152.890 52.820 152.950 ;
        RECT 56.640 152.890 56.960 153.150 ;
        RECT 62.235 153.135 62.525 153.450 ;
        RECT 65.855 153.430 66.145 153.475 ;
        RECT 66.760 153.430 67.080 153.490 ;
        RECT 65.855 153.290 67.080 153.430 ;
        RECT 65.855 153.245 66.145 153.290 ;
        RECT 66.760 153.230 67.080 153.290 ;
        RECT 71.820 153.230 72.140 153.490 ;
        RECT 74.120 153.230 74.440 153.490 ;
        RECT 74.595 153.245 74.885 153.475 ;
        RECT 75.130 153.430 75.270 154.310 ;
        RECT 75.500 154.310 78.565 154.450 ;
        RECT 75.500 154.250 75.820 154.310 ;
        RECT 78.275 154.265 78.565 154.310 ;
        RECT 78.720 154.450 79.040 154.510 ;
        RECT 80.115 154.450 80.405 154.495 ;
        RECT 78.720 154.310 80.405 154.450 ;
        RECT 78.720 154.250 79.040 154.310 ;
        RECT 80.115 154.265 80.405 154.310 ;
        RECT 82.400 154.250 82.720 154.510 ;
        RECT 82.860 154.250 83.180 154.510 ;
        RECT 87.000 154.250 87.320 154.510 ;
        RECT 88.380 154.450 88.700 154.510 ;
        RECT 88.855 154.450 89.145 154.495 ;
        RECT 88.380 154.310 89.145 154.450 ;
        RECT 88.380 154.250 88.700 154.310 ;
        RECT 88.855 154.265 89.145 154.310 ;
        RECT 95.740 154.250 96.060 154.510 ;
        RECT 101.275 154.450 101.565 154.495 ;
        RECT 101.720 154.450 102.040 154.510 ;
        RECT 101.275 154.310 102.040 154.450 ;
        RECT 101.275 154.265 101.565 154.310 ;
        RECT 101.720 154.250 102.040 154.310 ;
        RECT 106.780 154.450 107.100 154.510 ;
        RECT 112.315 154.450 112.605 154.495 ;
        RECT 106.780 154.310 112.605 154.450 ;
        RECT 106.780 154.250 107.100 154.310 ;
        RECT 112.315 154.265 112.605 154.310 ;
        RECT 114.155 154.450 114.445 154.495 ;
        RECT 115.520 154.450 115.840 154.510 ;
        RECT 114.155 154.310 115.840 154.450 ;
        RECT 114.155 154.265 114.445 154.310 ;
        RECT 115.520 154.250 115.840 154.310 ;
        RECT 117.820 154.450 118.140 154.510 ;
        RECT 118.295 154.450 118.585 154.495 ;
        RECT 117.820 154.310 118.585 154.450 ;
        RECT 117.820 154.250 118.140 154.310 ;
        RECT 118.295 154.265 118.585 154.310 ;
        RECT 119.660 154.250 119.980 154.510 ;
        RECT 121.500 154.250 121.820 154.510 ;
        RECT 123.290 154.450 123.580 154.495 ;
        RECT 124.260 154.450 124.580 154.510 ;
        RECT 123.290 154.310 124.580 154.450 ;
        RECT 123.290 154.265 123.580 154.310 ;
        RECT 124.260 154.250 124.580 154.310 ;
        RECT 130.700 154.250 131.020 154.510 ;
        RECT 131.160 154.450 131.480 154.510 ;
        RECT 132.095 154.450 132.385 154.495 ;
        RECT 131.160 154.310 132.385 154.450 ;
        RECT 131.160 154.250 131.480 154.310 ;
        RECT 132.095 154.265 132.385 154.310 ;
        RECT 75.960 154.110 76.280 154.170 ;
        RECT 80.575 154.110 80.865 154.155 ;
        RECT 82.950 154.110 83.090 154.250 ;
        RECT 75.960 153.970 80.865 154.110 ;
        RECT 75.960 153.910 76.280 153.970 ;
        RECT 80.575 153.925 80.865 153.970 ;
        RECT 82.030 153.970 83.090 154.110 ;
        RECT 83.320 154.110 83.640 154.170 ;
        RECT 93.455 154.110 93.745 154.155 ;
        RECT 83.320 153.970 93.745 154.110 ;
        RECT 76.420 153.770 76.740 153.830 ;
        RECT 82.030 153.815 82.170 153.970 ;
        RECT 83.320 153.910 83.640 153.970 ;
        RECT 93.455 153.925 93.745 153.970 ;
        RECT 76.420 153.630 79.410 153.770 ;
        RECT 76.420 153.570 76.740 153.630 ;
        RECT 78.275 153.430 78.565 153.475 ;
        RECT 75.130 153.290 78.565 153.430 ;
        RECT 78.275 153.245 78.565 153.290 ;
        RECT 78.735 153.245 79.025 153.475 ;
        RECT 79.270 153.430 79.410 153.630 ;
        RECT 81.955 153.585 82.245 153.815 ;
        RECT 84.240 153.570 84.560 153.830 ;
        RECT 84.700 153.570 85.020 153.830 ;
        RECT 91.615 153.770 91.905 153.815 ;
        RECT 85.710 153.630 91.905 153.770 ;
        RECT 82.415 153.430 82.705 153.475 ;
        RECT 79.270 153.290 82.705 153.430 ;
        RECT 82.415 153.245 82.705 153.290 ;
        RECT 83.780 153.430 84.100 153.490 ;
        RECT 85.175 153.430 85.465 153.475 ;
        RECT 83.780 153.290 85.465 153.430 ;
        RECT 58.935 153.090 59.585 153.135 ;
        RECT 62.235 153.090 62.825 153.135 ;
        RECT 63.540 153.090 63.860 153.150 ;
        RECT 58.935 152.950 63.860 153.090 ;
        RECT 58.935 152.905 59.585 152.950 ;
        RECT 62.535 152.905 62.825 152.950 ;
        RECT 63.540 152.890 63.860 152.950 ;
        RECT 64.460 152.890 64.780 153.150 ;
        RECT 70.900 153.090 71.220 153.150 ;
        RECT 74.210 153.090 74.350 153.230 ;
        RECT 67.770 152.950 71.220 153.090 ;
        RECT 50.660 152.610 51.350 152.750 ;
        RECT 53.880 152.750 54.200 152.810 ;
        RECT 64.000 152.750 64.320 152.810 ;
        RECT 67.770 152.795 67.910 152.950 ;
        RECT 70.900 152.890 71.220 152.950 ;
        RECT 72.370 152.950 74.350 153.090 ;
        RECT 74.670 153.090 74.810 153.245 ;
        RECT 74.670 152.950 76.650 153.090 ;
        RECT 53.880 152.610 64.320 152.750 ;
        RECT 50.660 152.550 50.980 152.610 ;
        RECT 53.880 152.550 54.200 152.610 ;
        RECT 64.000 152.550 64.320 152.610 ;
        RECT 67.695 152.565 67.985 152.795 ;
        RECT 68.140 152.750 68.460 152.810 ;
        RECT 69.520 152.750 69.840 152.810 ;
        RECT 68.140 152.610 69.840 152.750 ;
        RECT 68.140 152.550 68.460 152.610 ;
        RECT 69.520 152.550 69.840 152.610 ;
        RECT 69.980 152.750 70.300 152.810 ;
        RECT 72.370 152.750 72.510 152.950 ;
        RECT 69.980 152.610 72.510 152.750 ;
        RECT 69.980 152.550 70.300 152.610 ;
        RECT 75.960 152.550 76.280 152.810 ;
        RECT 76.510 152.750 76.650 152.950 ;
        RECT 77.340 152.890 77.660 153.150 ;
        RECT 78.810 153.090 78.950 153.245 ;
        RECT 78.810 152.950 82.170 153.090 ;
        RECT 82.030 152.810 82.170 152.950 ;
        RECT 77.800 152.750 78.120 152.810 ;
        RECT 76.510 152.610 78.120 152.750 ;
        RECT 77.800 152.550 78.120 152.610 ;
        RECT 81.940 152.550 82.260 152.810 ;
        RECT 82.490 152.750 82.630 153.245 ;
        RECT 83.780 153.230 84.100 153.290 ;
        RECT 85.175 153.245 85.465 153.290 ;
        RECT 82.860 153.090 83.180 153.150 ;
        RECT 85.710 153.090 85.850 153.630 ;
        RECT 91.615 153.585 91.905 153.630 ;
        RECT 89.760 153.230 90.080 153.490 ;
        RECT 90.220 153.430 90.540 153.490 ;
        RECT 94.375 153.430 94.665 153.475 ;
        RECT 90.220 153.290 94.665 153.430 ;
        RECT 90.220 153.230 90.540 153.290 ;
        RECT 94.375 153.245 94.665 153.290 ;
        RECT 89.850 153.090 89.990 153.230 ;
        RECT 90.695 153.090 90.985 153.135 ;
        RECT 82.860 152.950 85.850 153.090 ;
        RECT 86.170 152.950 89.990 153.090 ;
        RECT 90.310 152.950 90.985 153.090 ;
        RECT 82.860 152.890 83.180 152.950 ;
        RECT 86.170 152.750 86.310 152.950 ;
        RECT 82.490 152.610 86.310 152.750 ;
        RECT 89.760 152.750 90.080 152.810 ;
        RECT 90.310 152.750 90.450 152.950 ;
        RECT 90.695 152.905 90.985 152.950 ;
        RECT 91.155 153.090 91.445 153.135 ;
        RECT 92.060 153.090 92.380 153.150 ;
        RECT 91.155 152.950 92.380 153.090 ;
        RECT 95.830 153.090 95.970 154.250 ;
        RECT 96.200 154.110 96.520 154.170 ;
        RECT 104.445 154.110 104.735 154.155 ;
        RECT 106.335 154.110 106.625 154.155 ;
        RECT 109.455 154.110 109.745 154.155 ;
        RECT 122.845 154.110 123.135 154.155 ;
        RECT 124.735 154.110 125.025 154.155 ;
        RECT 127.855 154.110 128.145 154.155 ;
        RECT 96.200 153.970 103.790 154.110 ;
        RECT 96.200 153.910 96.520 153.970 ;
        RECT 98.515 153.585 98.805 153.815 ;
        RECT 98.590 153.430 98.730 153.585 ;
        RECT 98.960 153.570 99.280 153.830 ;
        RECT 102.180 153.570 102.500 153.830 ;
        RECT 103.650 153.815 103.790 153.970 ;
        RECT 104.445 153.970 109.745 154.110 ;
        RECT 104.445 153.925 104.735 153.970 ;
        RECT 106.335 153.925 106.625 153.970 ;
        RECT 109.455 153.925 109.745 153.970 ;
        RECT 112.850 153.970 122.190 154.110 ;
        RECT 112.850 153.830 112.990 153.970 ;
        RECT 103.575 153.770 103.865 153.815 ;
        RECT 112.760 153.770 113.080 153.830 ;
        RECT 103.575 153.630 113.080 153.770 ;
        RECT 103.575 153.585 103.865 153.630 ;
        RECT 112.760 153.570 113.080 153.630 ;
        RECT 115.520 153.570 115.840 153.830 ;
        RECT 115.980 153.570 116.300 153.830 ;
        RECT 116.440 153.570 116.760 153.830 ;
        RECT 118.740 153.570 119.060 153.830 ;
        RECT 122.050 153.815 122.190 153.970 ;
        RECT 122.845 153.970 128.145 154.110 ;
        RECT 122.845 153.925 123.135 153.970 ;
        RECT 124.735 153.925 125.025 153.970 ;
        RECT 127.855 153.925 128.145 153.970 ;
        RECT 121.975 153.770 122.265 153.815 ;
        RECT 123.340 153.770 123.660 153.830 ;
        RECT 121.975 153.630 123.660 153.770 ;
        RECT 132.170 153.770 132.310 154.265 ;
        RECT 137.600 154.250 137.920 154.510 ;
        RECT 138.995 154.450 139.285 154.495 ;
        RECT 143.120 154.450 143.440 154.510 ;
        RECT 138.995 154.310 143.440 154.450 ;
        RECT 138.995 154.265 139.285 154.310 ;
        RECT 143.120 154.250 143.440 154.310 ;
        RECT 137.140 153.910 137.460 154.170 ;
        RECT 134.855 153.770 135.145 153.815 ;
        RECT 132.170 153.630 135.145 153.770 ;
        RECT 121.975 153.585 122.265 153.630 ;
        RECT 123.340 153.570 123.660 153.630 ;
        RECT 134.855 153.585 135.145 153.630 ;
        RECT 102.270 153.430 102.410 153.570 ;
        RECT 98.590 153.290 102.410 153.430 ;
        RECT 104.040 153.430 104.330 153.475 ;
        RECT 105.875 153.430 106.165 153.475 ;
        RECT 109.455 153.430 109.745 153.475 ;
        RECT 104.040 153.290 109.745 153.430 ;
        RECT 104.040 153.245 104.330 153.290 ;
        RECT 105.875 153.245 106.165 153.290 ;
        RECT 109.455 153.245 109.745 153.290 ;
        RECT 110.000 153.430 110.320 153.490 ;
        RECT 110.535 153.430 110.825 153.450 ;
        RECT 110.000 153.290 110.825 153.430 ;
        RECT 110.000 153.230 110.320 153.290 ;
        RECT 99.435 153.090 99.725 153.135 ;
        RECT 95.830 152.950 99.725 153.090 ;
        RECT 91.155 152.905 91.445 152.950 ;
        RECT 92.060 152.890 92.380 152.950 ;
        RECT 99.435 152.905 99.725 152.950 ;
        RECT 101.260 153.090 101.580 153.150 ;
        RECT 110.535 153.135 110.825 153.290 ;
        RECT 112.300 153.230 112.620 153.490 ;
        RECT 113.235 153.430 113.525 153.475 ;
        RECT 116.530 153.430 116.670 153.570 ;
        RECT 113.235 153.290 116.670 153.430 ;
        RECT 118.830 153.430 118.970 153.570 ;
        RECT 119.240 153.430 119.530 153.475 ;
        RECT 122.440 153.430 122.730 153.475 ;
        RECT 124.275 153.430 124.565 153.475 ;
        RECT 127.855 153.430 128.145 153.475 ;
        RECT 118.830 153.290 122.190 153.430 ;
        RECT 113.235 153.245 113.525 153.290 ;
        RECT 119.240 153.245 119.530 153.290 ;
        RECT 104.955 153.090 105.245 153.135 ;
        RECT 101.260 152.950 105.245 153.090 ;
        RECT 101.260 152.890 101.580 152.950 ;
        RECT 104.955 152.905 105.245 152.950 ;
        RECT 107.235 153.090 107.885 153.135 ;
        RECT 110.535 153.090 111.125 153.135 ;
        RECT 107.235 152.950 111.125 153.090 ;
        RECT 112.390 153.090 112.530 153.230 ;
        RECT 119.660 153.090 119.980 153.150 ;
        RECT 112.390 152.950 119.980 153.090 ;
        RECT 122.050 153.090 122.190 153.290 ;
        RECT 122.440 153.290 128.145 153.430 ;
        RECT 122.440 153.245 122.730 153.290 ;
        RECT 124.275 153.245 124.565 153.290 ;
        RECT 127.855 153.245 128.145 153.290 ;
        RECT 128.860 153.450 129.180 153.490 ;
        RECT 128.860 153.230 129.225 153.450 ;
        RECT 137.690 153.430 137.830 154.250 ;
        RECT 138.075 153.430 138.365 153.475 ;
        RECT 123.800 153.090 124.120 153.150 ;
        RECT 128.935 153.135 129.225 153.230 ;
        RECT 133.550 153.290 135.070 153.430 ;
        RECT 137.690 153.290 138.365 153.430 ;
        RECT 133.550 153.150 133.690 153.290 ;
        RECT 122.050 152.950 124.120 153.090 ;
        RECT 107.235 152.905 107.885 152.950 ;
        RECT 110.835 152.905 111.125 152.950 ;
        RECT 119.660 152.890 119.980 152.950 ;
        RECT 123.800 152.890 124.120 152.950 ;
        RECT 125.635 153.090 126.285 153.135 ;
        RECT 128.935 153.090 129.525 153.135 ;
        RECT 125.635 152.950 129.525 153.090 ;
        RECT 125.635 152.905 126.285 152.950 ;
        RECT 129.235 152.905 129.525 152.950 ;
        RECT 133.460 152.890 133.780 153.150 ;
        RECT 134.930 153.135 135.070 153.290 ;
        RECT 138.075 153.245 138.365 153.290 ;
        RECT 140.375 153.430 140.665 153.475 ;
        RECT 140.820 153.430 141.140 153.490 ;
        RECT 140.375 153.290 141.140 153.430 ;
        RECT 140.375 153.245 140.665 153.290 ;
        RECT 140.820 153.230 141.140 153.290 ;
        RECT 134.395 152.905 134.685 153.135 ;
        RECT 134.855 152.905 135.145 153.135 ;
        RECT 89.760 152.610 90.450 152.750 ;
        RECT 97.580 152.750 97.900 152.810 ;
        RECT 108.620 152.750 108.940 152.810 ;
        RECT 97.580 152.610 108.940 152.750 ;
        RECT 89.760 152.550 90.080 152.610 ;
        RECT 97.580 152.550 97.900 152.610 ;
        RECT 108.620 152.550 108.940 152.610 ;
        RECT 116.455 152.750 116.745 152.795 ;
        RECT 116.900 152.750 117.220 152.810 ;
        RECT 116.455 152.610 117.220 152.750 ;
        RECT 116.455 152.565 116.745 152.610 ;
        RECT 116.900 152.550 117.220 152.610 ;
        RECT 117.820 152.750 118.140 152.810 ;
        RECT 126.560 152.750 126.880 152.810 ;
        RECT 134.470 152.750 134.610 152.905 ;
        RECT 117.820 152.610 134.610 152.750 ;
        RECT 139.455 152.750 139.745 152.795 ;
        RECT 139.900 152.750 140.220 152.810 ;
        RECT 139.455 152.610 140.220 152.750 ;
        RECT 117.820 152.550 118.140 152.610 ;
        RECT 126.560 152.550 126.880 152.610 ;
        RECT 139.455 152.565 139.745 152.610 ;
        RECT 139.900 152.550 140.220 152.610 ;
        RECT 2.750 151.930 159.030 152.410 ;
        RECT 7.880 151.730 8.200 151.790 ;
        RECT 18.460 151.730 18.780 151.790 ;
        RECT 7.880 151.590 18.780 151.730 ;
        RECT 7.880 151.530 8.200 151.590 ;
        RECT 18.460 151.530 18.780 151.590 ;
        RECT 23.995 151.730 24.285 151.775 ;
        RECT 35.020 151.730 35.340 151.790 ;
        RECT 23.995 151.590 35.340 151.730 ;
        RECT 23.995 151.545 24.285 151.590 ;
        RECT 35.020 151.530 35.340 151.590 ;
        RECT 37.780 151.730 38.100 151.790 ;
        RECT 44.220 151.730 44.540 151.790 ;
        RECT 50.200 151.730 50.520 151.790 ;
        RECT 37.780 151.590 44.540 151.730 ;
        RECT 37.780 151.530 38.100 151.590 ;
        RECT 44.220 151.530 44.540 151.590 ;
        RECT 45.230 151.590 49.510 151.730 ;
        RECT 8.800 151.390 9.120 151.450 ;
        RECT 11.115 151.390 11.405 151.435 ;
        RECT 8.800 151.250 11.405 151.390 ;
        RECT 8.800 151.190 9.120 151.250 ;
        RECT 11.115 151.205 11.405 151.250 ;
        RECT 13.395 151.390 14.045 151.435 ;
        RECT 16.995 151.390 17.285 151.435 ;
        RECT 38.240 151.390 38.560 151.450 ;
        RECT 13.395 151.250 17.285 151.390 ;
        RECT 13.395 151.205 14.045 151.250 ;
        RECT 16.695 151.205 17.285 151.250 ;
        RECT 24.530 151.250 38.560 151.390 ;
        RECT 5.135 151.050 5.425 151.095 ;
        RECT 3.830 150.910 5.425 151.050 ;
        RECT 3.830 150.030 3.970 150.910 ;
        RECT 5.135 150.865 5.425 150.910 ;
        RECT 5.580 151.050 5.900 151.110 ;
        RECT 6.515 151.050 6.805 151.095 ;
        RECT 5.580 150.910 6.805 151.050 ;
        RECT 5.580 150.850 5.900 150.910 ;
        RECT 6.515 150.865 6.805 150.910 ;
        RECT 6.975 151.050 7.265 151.095 ;
        RECT 7.420 151.050 7.740 151.110 ;
        RECT 6.975 150.910 7.740 151.050 ;
        RECT 6.975 150.865 7.265 150.910 ;
        RECT 7.420 150.850 7.740 150.910 ;
        RECT 7.880 150.850 8.200 151.110 ;
        RECT 8.355 150.865 8.645 151.095 ;
        RECT 10.200 151.050 10.490 151.095 ;
        RECT 12.035 151.050 12.325 151.095 ;
        RECT 15.615 151.050 15.905 151.095 ;
        RECT 10.200 150.910 15.905 151.050 ;
        RECT 10.200 150.865 10.490 150.910 ;
        RECT 12.035 150.865 12.325 150.910 ;
        RECT 15.615 150.865 15.905 150.910 ;
        RECT 16.695 150.890 16.985 151.205 ;
        RECT 24.530 151.095 24.670 151.250 ;
        RECT 38.240 151.190 38.560 151.250 ;
        RECT 41.460 151.390 41.780 151.450 ;
        RECT 42.855 151.390 43.145 151.435 ;
        RECT 41.460 151.250 43.530 151.390 ;
        RECT 41.460 151.190 41.780 151.250 ;
        RECT 42.855 151.205 43.145 151.250 ;
        RECT 43.390 151.110 43.530 151.250 ;
        RECT 8.430 150.430 8.570 150.865 ;
        RECT 9.720 150.510 10.040 150.770 ;
        RECT 11.100 150.710 11.420 150.770 ;
        RECT 16.710 150.710 16.850 150.890 ;
        RECT 24.455 150.865 24.745 151.095 ;
        RECT 26.280 150.850 26.600 151.110 ;
        RECT 26.740 150.850 27.060 151.110 ;
        RECT 27.200 151.050 27.520 151.110 ;
        RECT 27.200 150.910 27.890 151.050 ;
        RECT 27.200 150.850 27.520 150.910 ;
        RECT 11.100 150.570 16.850 150.710 ;
        RECT 17.540 150.710 17.860 150.770 ;
        RECT 18.475 150.710 18.765 150.755 ;
        RECT 21.695 150.710 21.985 150.755 ;
        RECT 17.540 150.570 21.985 150.710 ;
        RECT 27.750 150.710 27.890 150.910 ;
        RECT 28.580 150.850 28.900 151.110 ;
        RECT 29.040 151.050 29.360 151.110 ;
        RECT 30.435 151.050 30.725 151.095 ;
        RECT 29.040 150.910 30.725 151.050 ;
        RECT 29.040 150.850 29.360 150.910 ;
        RECT 30.435 150.865 30.725 150.910 ;
        RECT 30.895 151.050 31.185 151.095 ;
        RECT 30.895 150.910 31.570 151.050 ;
        RECT 30.895 150.865 31.185 150.910 ;
        RECT 28.135 150.710 28.425 150.755 ;
        RECT 27.750 150.570 28.425 150.710 ;
        RECT 28.670 150.710 28.810 150.850 ;
        RECT 29.515 150.710 29.805 150.755 ;
        RECT 28.670 150.570 29.805 150.710 ;
        RECT 11.100 150.510 11.420 150.570 ;
        RECT 17.540 150.510 17.860 150.570 ;
        RECT 18.475 150.525 18.765 150.570 ;
        RECT 21.695 150.525 21.985 150.570 ;
        RECT 28.135 150.525 28.425 150.570 ;
        RECT 29.515 150.525 29.805 150.570 ;
        RECT 6.055 150.185 6.345 150.415 ;
        RECT 2.450 149.890 3.970 150.030 ;
        RECT 6.130 150.030 6.270 150.185 ;
        RECT 8.340 150.170 8.660 150.430 ;
        RECT 10.605 150.370 10.895 150.415 ;
        RECT 12.495 150.370 12.785 150.415 ;
        RECT 15.615 150.370 15.905 150.415 ;
        RECT 19.840 150.370 20.160 150.430 ;
        RECT 10.605 150.230 15.905 150.370 ;
        RECT 10.605 150.185 10.895 150.230 ;
        RECT 12.495 150.185 12.785 150.230 ;
        RECT 15.615 150.185 15.905 150.230 ;
        RECT 18.550 150.230 20.160 150.370 ;
        RECT 8.800 150.030 9.120 150.090 ;
        RECT 6.130 149.890 9.120 150.030 ;
        RECT 2.450 149.010 2.590 149.890 ;
        RECT 8.800 149.830 9.120 149.890 ;
        RECT 9.275 150.030 9.565 150.075 ;
        RECT 18.550 150.030 18.690 150.230 ;
        RECT 19.840 150.170 20.160 150.230 ;
        RECT 26.280 150.370 26.600 150.430 ;
        RECT 31.430 150.370 31.570 150.910 ;
        RECT 32.260 150.850 32.580 151.110 ;
        RECT 33.640 150.850 33.960 151.110 ;
        RECT 34.100 150.850 34.420 151.110 ;
        RECT 35.020 150.850 35.340 151.110 ;
        RECT 35.495 150.865 35.785 151.095 ;
        RECT 39.635 150.865 39.925 151.095 ;
        RECT 40.080 151.050 40.400 151.110 ;
        RECT 41.935 151.050 42.225 151.095 ;
        RECT 40.080 150.910 42.225 151.050 ;
        RECT 31.815 150.710 32.105 150.755 ;
        RECT 35.570 150.710 35.710 150.865 ;
        RECT 36.860 150.710 37.180 150.770 ;
        RECT 31.815 150.570 34.560 150.710 ;
        RECT 35.570 150.570 37.180 150.710 ;
        RECT 31.815 150.525 32.105 150.570 ;
        RECT 26.280 150.230 31.570 150.370 ;
        RECT 26.280 150.170 26.600 150.230 ;
        RECT 9.275 149.890 18.690 150.030 ;
        RECT 9.275 149.845 9.565 149.890 ;
        RECT 18.920 149.830 19.240 150.090 ;
        RECT 23.520 150.030 23.840 150.090 ;
        RECT 24.440 150.030 24.760 150.090 ;
        RECT 23.520 149.890 24.760 150.030 ;
        RECT 23.520 149.830 23.840 149.890 ;
        RECT 24.440 149.830 24.760 149.890 ;
        RECT 25.375 150.030 25.665 150.075 ;
        RECT 27.200 150.030 27.520 150.090 ;
        RECT 25.375 149.890 27.520 150.030 ;
        RECT 25.375 149.845 25.665 149.890 ;
        RECT 27.200 149.830 27.520 149.890 ;
        RECT 27.675 150.030 27.965 150.075 ;
        RECT 28.580 150.030 28.900 150.090 ;
        RECT 31.890 150.030 32.030 150.525 ;
        RECT 34.420 150.370 34.560 150.570 ;
        RECT 36.860 150.510 37.180 150.570 ;
        RECT 37.320 150.710 37.640 150.770 ;
        RECT 39.710 150.710 39.850 150.865 ;
        RECT 40.080 150.850 40.400 150.910 ;
        RECT 41.935 150.865 42.225 150.910 ;
        RECT 37.320 150.570 39.850 150.710 ;
        RECT 42.010 150.710 42.150 150.865 ;
        RECT 42.380 150.850 42.700 151.110 ;
        RECT 43.300 150.850 43.620 151.110 ;
        RECT 43.760 150.850 44.080 151.110 ;
        RECT 44.310 151.050 44.450 151.530 ;
        RECT 44.310 150.910 44.730 151.050 ;
        RECT 42.840 150.710 43.160 150.770 ;
        RECT 42.010 150.570 43.160 150.710 ;
        RECT 44.590 150.710 44.730 150.910 ;
        RECT 45.230 150.710 45.370 151.590 ;
        RECT 49.370 151.435 49.510 151.590 ;
        RECT 49.830 151.590 50.520 151.730 ;
        RECT 49.830 151.435 49.970 151.590 ;
        RECT 50.200 151.530 50.520 151.590 ;
        RECT 53.420 151.530 53.740 151.790 ;
        RECT 55.260 151.530 55.580 151.790 ;
        RECT 55.735 151.730 56.025 151.775 ;
        RECT 60.320 151.730 60.640 151.790 ;
        RECT 55.735 151.590 60.640 151.730 ;
        RECT 55.735 151.545 56.025 151.590 ;
        RECT 60.320 151.530 60.640 151.590 ;
        RECT 62.175 151.730 62.465 151.775 ;
        RECT 64.920 151.730 65.240 151.790 ;
        RECT 65.840 151.730 66.160 151.790 ;
        RECT 62.175 151.590 66.160 151.730 ;
        RECT 62.175 151.545 62.465 151.590 ;
        RECT 64.920 151.530 65.240 151.590 ;
        RECT 65.840 151.530 66.160 151.590 ;
        RECT 71.820 151.530 72.140 151.790 ;
        RECT 77.800 151.730 78.120 151.790 ;
        RECT 82.860 151.730 83.180 151.790 ;
        RECT 77.800 151.590 83.180 151.730 ;
        RECT 77.800 151.530 78.120 151.590 ;
        RECT 82.860 151.530 83.180 151.590 ;
        RECT 83.780 151.730 84.100 151.790 ;
        RECT 120.580 151.730 120.900 151.790 ;
        RECT 83.780 151.590 120.900 151.730 ;
        RECT 83.780 151.530 84.100 151.590 ;
        RECT 120.580 151.530 120.900 151.590 ;
        RECT 122.420 151.530 122.740 151.790 ;
        RECT 123.340 151.730 123.660 151.790 ;
        RECT 127.035 151.730 127.325 151.775 ;
        RECT 128.400 151.730 128.720 151.790 ;
        RECT 123.340 151.590 125.870 151.730 ;
        RECT 123.340 151.530 123.660 151.590 ;
        RECT 49.295 151.205 49.585 151.435 ;
        RECT 49.755 151.205 50.045 151.435 ;
        RECT 55.350 151.390 55.490 151.530 ;
        RECT 62.635 151.390 62.925 151.435 ;
        RECT 55.350 151.250 62.925 151.390 ;
        RECT 62.635 151.205 62.925 151.250 ;
        RECT 64.000 151.390 64.320 151.450 ;
        RECT 64.000 151.250 65.610 151.390 ;
        RECT 45.615 150.865 45.905 151.095 ;
        RECT 46.075 151.050 46.365 151.095 ;
        RECT 46.520 151.050 46.840 151.110 ;
        RECT 46.075 150.910 46.840 151.050 ;
        RECT 46.075 150.865 46.365 150.910 ;
        RECT 44.590 150.570 45.370 150.710 ;
        RECT 37.320 150.510 37.640 150.570 ;
        RECT 42.840 150.510 43.160 150.570 ;
        RECT 35.020 150.370 35.340 150.430 ;
        RECT 39.620 150.370 39.940 150.430 ;
        RECT 34.420 150.230 35.340 150.370 ;
        RECT 35.020 150.170 35.340 150.230 ;
        RECT 35.570 150.230 39.940 150.370 ;
        RECT 35.570 150.090 35.710 150.230 ;
        RECT 39.620 150.170 39.940 150.230 ;
        RECT 43.300 150.370 43.620 150.430 ;
        RECT 45.690 150.370 45.830 150.865 ;
        RECT 46.520 150.850 46.840 150.910 ;
        RECT 48.360 150.850 48.680 151.110 ;
        RECT 50.215 151.050 50.505 151.095 ;
        RECT 52.515 151.050 52.805 151.095 ;
        RECT 49.370 150.910 50.505 151.050 ;
        RECT 49.370 150.770 49.510 150.910 ;
        RECT 50.215 150.865 50.505 150.910 ;
        RECT 51.210 150.910 52.805 151.050 ;
        RECT 47.455 150.525 47.745 150.755 ;
        RECT 43.300 150.230 45.830 150.370 ;
        RECT 47.530 150.370 47.670 150.525 ;
        RECT 49.280 150.510 49.600 150.770 ;
        RECT 49.740 150.510 50.060 150.770 ;
        RECT 49.830 150.370 49.970 150.510 ;
        RECT 51.210 150.415 51.350 150.910 ;
        RECT 52.515 150.865 52.805 150.910 ;
        RECT 53.880 150.850 54.200 151.110 ;
        RECT 54.800 150.850 55.120 151.110 ;
        RECT 58.035 151.050 58.325 151.095 ;
        RECT 62.710 151.050 62.850 151.205 ;
        RECT 64.000 151.190 64.320 151.250 ;
        RECT 64.920 151.050 65.240 151.110 ;
        RECT 55.350 150.910 57.790 151.050 ;
        RECT 51.580 150.710 51.900 150.770 ;
        RECT 53.420 150.710 53.740 150.770 ;
        RECT 55.350 150.710 55.490 150.910 ;
        RECT 51.580 150.570 55.490 150.710 ;
        RECT 57.650 150.710 57.790 150.910 ;
        RECT 58.035 150.910 62.160 151.050 ;
        RECT 62.710 150.910 65.240 151.050 ;
        RECT 58.035 150.865 58.325 150.910 ;
        RECT 58.495 150.710 58.785 150.755 ;
        RECT 58.940 150.710 59.260 150.770 ;
        RECT 57.650 150.570 59.260 150.710 ;
        RECT 51.580 150.510 51.900 150.570 ;
        RECT 53.420 150.510 53.740 150.570 ;
        RECT 58.495 150.525 58.785 150.570 ;
        RECT 58.940 150.510 59.260 150.570 ;
        RECT 59.400 150.510 59.720 150.770 ;
        RECT 47.530 150.230 49.970 150.370 ;
        RECT 43.300 150.170 43.620 150.230 ;
        RECT 51.135 150.185 51.425 150.415 ;
        RECT 55.260 150.370 55.580 150.430 ;
        RECT 60.335 150.370 60.625 150.415 ;
        RECT 55.260 150.230 60.625 150.370 ;
        RECT 62.020 150.370 62.160 150.910 ;
        RECT 64.920 150.850 65.240 150.910 ;
        RECT 63.080 150.510 63.400 150.770 ;
        RECT 65.470 150.710 65.610 151.250 ;
        RECT 66.760 151.050 67.080 151.110 ;
        RECT 68.155 151.050 68.445 151.095 ;
        RECT 66.760 150.910 68.445 151.050 ;
        RECT 66.760 150.850 67.080 150.910 ;
        RECT 68.155 150.865 68.445 150.910 ;
        RECT 69.075 151.050 69.365 151.095 ;
        RECT 71.910 151.050 72.050 151.530 ;
        RECT 78.260 151.190 78.580 151.450 ;
        RECT 81.955 151.390 82.245 151.435 ;
        RECT 83.320 151.390 83.640 151.450 ;
        RECT 81.955 151.250 83.640 151.390 ;
        RECT 81.955 151.205 82.245 151.250 ;
        RECT 83.320 151.190 83.640 151.250 ;
        RECT 84.235 151.390 84.885 151.435 ;
        RECT 85.160 151.390 85.480 151.450 ;
        RECT 87.835 151.390 88.125 151.435 ;
        RECT 94.820 151.390 95.140 151.450 ;
        RECT 98.500 151.435 98.820 151.450 ;
        RECT 84.235 151.250 88.125 151.390 ;
        RECT 84.235 151.205 84.885 151.250 ;
        RECT 85.160 151.190 85.480 151.250 ;
        RECT 87.535 151.205 88.125 151.250 ;
        RECT 91.690 151.250 95.140 151.390 ;
        RECT 69.075 150.910 72.050 151.050 ;
        RECT 81.040 151.050 81.330 151.095 ;
        RECT 82.875 151.050 83.165 151.095 ;
        RECT 86.455 151.050 86.745 151.095 ;
        RECT 81.040 150.910 86.745 151.050 ;
        RECT 69.075 150.865 69.365 150.910 ;
        RECT 81.040 150.865 81.330 150.910 ;
        RECT 82.875 150.865 83.165 150.910 ;
        RECT 86.455 150.865 86.745 150.910 ;
        RECT 87.535 150.890 87.825 151.205 ;
        RECT 88.010 150.910 90.910 151.050 ;
        RECT 67.235 150.710 67.525 150.755 ;
        RECT 65.470 150.570 67.525 150.710 ;
        RECT 68.230 150.710 68.370 150.865 ;
        RECT 88.010 150.770 88.150 150.910 ;
        RECT 76.420 150.710 76.740 150.770 ;
        RECT 68.230 150.570 76.740 150.710 ;
        RECT 67.235 150.525 67.525 150.570 ;
        RECT 76.420 150.510 76.740 150.570 ;
        RECT 80.575 150.525 80.865 150.755 ;
        RECT 85.160 150.710 85.480 150.770 ;
        RECT 85.160 150.570 87.690 150.710 ;
        RECT 64.475 150.370 64.765 150.415 ;
        RECT 71.835 150.370 72.125 150.415 ;
        RECT 80.650 150.370 80.790 150.525 ;
        RECT 85.160 150.510 85.480 150.570 ;
        RECT 62.020 150.230 64.765 150.370 ;
        RECT 55.260 150.170 55.580 150.230 ;
        RECT 60.335 150.185 60.625 150.230 ;
        RECT 64.475 150.185 64.765 150.230 ;
        RECT 67.310 150.230 80.790 150.370 ;
        RECT 81.445 150.370 81.735 150.415 ;
        RECT 83.335 150.370 83.625 150.415 ;
        RECT 86.455 150.370 86.745 150.415 ;
        RECT 81.445 150.230 86.745 150.370 ;
        RECT 87.550 150.370 87.690 150.570 ;
        RECT 87.920 150.510 88.240 150.770 ;
        RECT 88.380 150.710 88.700 150.770 ;
        RECT 89.315 150.710 89.605 150.755 ;
        RECT 88.380 150.570 89.605 150.710 ;
        RECT 90.770 150.710 90.910 150.910 ;
        RECT 91.140 150.850 91.460 151.110 ;
        RECT 91.690 151.095 91.830 151.250 ;
        RECT 94.820 151.190 95.140 151.250 ;
        RECT 98.425 151.205 98.820 151.435 ;
        RECT 100.815 151.205 101.105 151.435 ;
        RECT 101.275 151.390 101.565 151.435 ;
        RECT 102.180 151.390 102.500 151.450 ;
        RECT 101.275 151.250 102.500 151.390 ;
        RECT 101.275 151.205 101.565 151.250 ;
        RECT 98.500 151.190 98.820 151.205 ;
        RECT 91.615 150.865 91.905 151.095 ;
        RECT 92.535 151.050 92.825 151.095 ;
        RECT 92.980 151.050 93.300 151.110 ;
        RECT 92.535 150.910 93.300 151.050 ;
        RECT 92.535 150.865 92.825 150.910 ;
        RECT 92.610 150.710 92.750 150.865 ;
        RECT 92.980 150.850 93.300 150.910 ;
        RECT 96.660 151.050 96.980 151.110 ;
        RECT 99.895 151.050 100.185 151.095 ;
        RECT 96.660 150.910 100.185 151.050 ;
        RECT 100.890 151.050 101.030 151.205 ;
        RECT 102.180 151.190 102.500 151.250 ;
        RECT 102.640 151.390 102.960 151.450 ;
        RECT 103.115 151.390 103.405 151.435 ;
        RECT 107.255 151.390 107.545 151.435 ;
        RECT 102.640 151.250 107.545 151.390 ;
        RECT 102.640 151.190 102.960 151.250 ;
        RECT 103.115 151.205 103.405 151.250 ;
        RECT 107.255 151.205 107.545 151.250 ;
        RECT 113.680 151.390 114.000 151.450 ;
        RECT 114.155 151.390 114.445 151.435 ;
        RECT 117.820 151.390 118.140 151.450 ;
        RECT 113.680 151.250 118.140 151.390 ;
        RECT 113.680 151.190 114.000 151.250 ;
        RECT 114.155 151.205 114.445 151.250 ;
        RECT 117.820 151.190 118.140 151.250 ;
        RECT 118.395 151.390 118.685 151.435 ;
        RECT 121.635 151.390 122.285 151.435 ;
        RECT 122.510 151.390 122.650 151.530 ;
        RECT 118.395 151.250 122.650 151.390 ;
        RECT 124.275 151.390 124.565 151.435 ;
        RECT 124.720 151.390 125.040 151.450 ;
        RECT 124.275 151.250 125.040 151.390 ;
        RECT 118.395 151.205 118.985 151.250 ;
        RECT 121.635 151.205 122.285 151.250 ;
        RECT 124.275 151.205 124.565 151.250 ;
        RECT 105.860 151.050 106.180 151.110 ;
        RECT 109.095 151.050 109.385 151.095 ;
        RECT 100.890 150.910 103.330 151.050 ;
        RECT 96.660 150.850 96.980 150.910 ;
        RECT 99.895 150.865 100.185 150.910 ;
        RECT 103.190 150.770 103.330 150.910 ;
        RECT 105.860 150.910 109.385 151.050 ;
        RECT 105.860 150.850 106.180 150.910 ;
        RECT 109.095 150.865 109.385 150.910 ;
        RECT 111.840 150.850 112.160 151.110 ;
        RECT 115.075 150.865 115.365 151.095 ;
        RECT 118.695 150.890 118.985 151.205 ;
        RECT 124.720 151.190 125.040 151.250 ;
        RECT 125.730 151.390 125.870 151.590 ;
        RECT 127.035 151.590 128.720 151.730 ;
        RECT 127.035 151.545 127.325 151.590 ;
        RECT 128.400 151.530 128.720 151.590 ;
        RECT 128.860 151.730 129.180 151.790 ;
        RECT 141.280 151.730 141.600 151.790 ;
        RECT 145.420 151.730 145.740 151.790 ;
        RECT 128.860 151.590 133.230 151.730 ;
        RECT 128.860 151.530 129.180 151.590 ;
        RECT 133.090 151.390 133.230 151.590 ;
        RECT 135.850 151.590 145.740 151.730 ;
        RECT 135.850 151.390 135.990 151.590 ;
        RECT 141.280 151.530 141.600 151.590 ;
        RECT 145.420 151.530 145.740 151.590 ;
        RECT 136.215 151.390 136.865 151.435 ;
        RECT 139.815 151.390 140.105 151.435 ;
        RECT 125.730 151.250 132.770 151.390 ;
        RECT 133.090 151.250 140.105 151.390 ;
        RECT 125.730 151.095 125.870 151.250 ;
        RECT 132.630 151.110 132.770 151.250 ;
        RECT 136.215 151.205 136.865 151.250 ;
        RECT 139.515 151.205 140.105 151.250 ;
        RECT 119.775 151.050 120.065 151.095 ;
        RECT 123.355 151.050 123.645 151.095 ;
        RECT 125.190 151.050 125.480 151.095 ;
        RECT 119.775 150.910 125.480 151.050 ;
        RECT 119.775 150.865 120.065 150.910 ;
        RECT 123.355 150.865 123.645 150.910 ;
        RECT 125.190 150.865 125.480 150.910 ;
        RECT 125.655 150.865 125.945 151.095 ;
        RECT 126.115 150.865 126.405 151.095 ;
        RECT 90.770 150.570 92.750 150.710 ;
        RECT 94.835 150.710 95.125 150.755 ;
        RECT 95.280 150.710 95.600 150.770 ;
        RECT 94.835 150.570 95.600 150.710 ;
        RECT 88.380 150.510 88.700 150.570 ;
        RECT 89.315 150.525 89.605 150.570 ;
        RECT 94.835 150.525 95.125 150.570 ;
        RECT 95.280 150.510 95.600 150.570 ;
        RECT 95.740 150.710 96.060 150.770 ;
        RECT 95.740 150.570 101.490 150.710 ;
        RECT 95.740 150.510 96.060 150.570 ;
        RECT 100.800 150.370 101.120 150.430 ;
        RECT 87.550 150.230 101.120 150.370 ;
        RECT 101.350 150.370 101.490 150.570 ;
        RECT 103.100 150.510 103.420 150.770 ;
        RECT 104.940 150.710 105.260 150.770 ;
        RECT 108.175 150.710 108.465 150.755 ;
        RECT 104.940 150.570 108.465 150.710 ;
        RECT 104.940 150.510 105.260 150.570 ;
        RECT 108.175 150.525 108.465 150.570 ;
        RECT 109.540 150.710 109.860 150.770 ;
        RECT 112.775 150.710 113.065 150.755 ;
        RECT 114.600 150.710 114.920 150.770 ;
        RECT 109.540 150.570 114.920 150.710 ;
        RECT 109.540 150.510 109.860 150.570 ;
        RECT 112.775 150.525 113.065 150.570 ;
        RECT 114.600 150.510 114.920 150.570 ;
        RECT 101.350 150.230 104.710 150.370 ;
        RECT 67.310 150.090 67.450 150.230 ;
        RECT 71.835 150.185 72.125 150.230 ;
        RECT 81.445 150.185 81.735 150.230 ;
        RECT 83.335 150.185 83.625 150.230 ;
        RECT 86.455 150.185 86.745 150.230 ;
        RECT 100.800 150.170 101.120 150.230 ;
        RECT 27.675 149.890 32.030 150.030 ;
        RECT 32.735 150.030 33.025 150.075 ;
        RECT 33.180 150.030 33.500 150.090 ;
        RECT 32.735 149.890 33.500 150.030 ;
        RECT 27.675 149.845 27.965 149.890 ;
        RECT 28.580 149.830 28.900 149.890 ;
        RECT 32.735 149.845 33.025 149.890 ;
        RECT 33.180 149.830 33.500 149.890 ;
        RECT 35.480 149.830 35.800 150.090 ;
        RECT 36.860 149.830 37.180 150.090 ;
        RECT 40.540 150.030 40.860 150.090 ;
        RECT 41.015 150.030 41.305 150.075 ;
        RECT 40.540 149.890 41.305 150.030 ;
        RECT 40.540 149.830 40.860 149.890 ;
        RECT 41.015 149.845 41.305 149.890 ;
        RECT 44.680 149.830 45.000 150.090 ;
        RECT 46.520 150.030 46.840 150.090 ;
        RECT 46.995 150.030 47.285 150.075 ;
        RECT 46.520 149.890 47.285 150.030 ;
        RECT 46.520 149.830 46.840 149.890 ;
        RECT 46.995 149.845 47.285 149.890 ;
        RECT 49.280 150.030 49.600 150.090 ;
        RECT 51.595 150.030 51.885 150.075 ;
        RECT 49.280 149.890 51.885 150.030 ;
        RECT 49.280 149.830 49.600 149.890 ;
        RECT 51.595 149.845 51.885 149.890 ;
        RECT 56.180 149.830 56.500 150.090 ;
        RECT 59.860 150.030 60.180 150.090 ;
        RECT 67.220 150.030 67.540 150.090 ;
        RECT 59.860 149.890 67.540 150.030 ;
        RECT 59.860 149.830 60.180 149.890 ;
        RECT 67.220 149.830 67.540 149.890 ;
        RECT 68.615 150.030 68.905 150.075 ;
        RECT 69.980 150.030 70.300 150.090 ;
        RECT 68.615 149.890 70.300 150.030 ;
        RECT 68.615 149.845 68.905 149.890 ;
        RECT 69.980 149.830 70.300 149.890 ;
        RECT 82.400 150.030 82.720 150.090 ;
        RECT 103.560 150.030 103.880 150.090 ;
        RECT 82.400 149.890 103.880 150.030 ;
        RECT 82.400 149.830 82.720 149.890 ;
        RECT 103.560 149.830 103.880 149.890 ;
        RECT 104.020 149.830 104.340 150.090 ;
        RECT 104.570 150.030 104.710 150.230 ;
        RECT 115.150 150.030 115.290 150.865 ;
        RECT 116.900 150.510 117.220 150.770 ;
        RECT 119.200 150.710 119.520 150.770 ;
        RECT 121.960 150.710 122.280 150.770 ;
        RECT 126.190 150.710 126.330 150.865 ;
        RECT 127.020 150.850 127.340 151.110 ;
        RECT 129.320 150.850 129.640 151.110 ;
        RECT 132.540 150.850 132.860 151.110 ;
        RECT 133.020 151.050 133.310 151.095 ;
        RECT 134.855 151.050 135.145 151.095 ;
        RECT 138.435 151.050 138.725 151.095 ;
        RECT 133.020 150.910 138.725 151.050 ;
        RECT 133.020 150.865 133.310 150.910 ;
        RECT 134.855 150.865 135.145 150.910 ;
        RECT 138.435 150.865 138.725 150.910 ;
        RECT 139.515 150.890 139.805 151.205 ;
        RECT 143.580 150.850 143.900 151.110 ;
        RECT 119.200 150.570 122.280 150.710 ;
        RECT 119.200 150.510 119.520 150.570 ;
        RECT 121.960 150.510 122.280 150.570 ;
        RECT 125.730 150.570 126.330 150.710 ;
        RECT 127.480 150.710 127.800 150.770 ;
        RECT 127.955 150.710 128.245 150.755 ;
        RECT 128.875 150.710 129.165 150.755 ;
        RECT 127.480 150.570 128.245 150.710 ;
        RECT 125.730 150.430 125.870 150.570 ;
        RECT 127.480 150.510 127.800 150.570 ;
        RECT 127.955 150.525 128.245 150.570 ;
        RECT 128.490 150.570 129.165 150.710 ;
        RECT 119.775 150.370 120.065 150.415 ;
        RECT 122.895 150.370 123.185 150.415 ;
        RECT 124.785 150.370 125.075 150.415 ;
        RECT 115.610 150.230 119.430 150.370 ;
        RECT 115.610 150.090 115.750 150.230 ;
        RECT 104.570 149.890 115.290 150.030 ;
        RECT 115.520 149.830 115.840 150.090 ;
        RECT 115.995 150.030 116.285 150.075 ;
        RECT 117.820 150.030 118.140 150.090 ;
        RECT 115.995 149.890 118.140 150.030 ;
        RECT 119.290 150.030 119.430 150.230 ;
        RECT 119.775 150.230 125.075 150.370 ;
        RECT 119.775 150.185 120.065 150.230 ;
        RECT 122.895 150.185 123.185 150.230 ;
        RECT 124.785 150.185 125.075 150.230 ;
        RECT 125.640 150.170 125.960 150.430 ;
        RECT 126.100 150.030 126.420 150.090 ;
        RECT 128.490 150.030 128.630 150.570 ;
        RECT 128.875 150.525 129.165 150.570 ;
        RECT 133.935 150.710 134.225 150.755 ;
        RECT 140.360 150.710 140.680 150.770 ;
        RECT 133.935 150.570 140.680 150.710 ;
        RECT 133.935 150.525 134.225 150.570 ;
        RECT 140.360 150.510 140.680 150.570 ;
        RECT 141.295 150.710 141.585 150.755 ;
        RECT 143.670 150.710 143.810 150.850 ;
        RECT 141.295 150.570 143.810 150.710 ;
        RECT 141.295 150.525 141.585 150.570 ;
        RECT 133.425 150.370 133.715 150.415 ;
        RECT 135.315 150.370 135.605 150.415 ;
        RECT 138.435 150.370 138.725 150.415 ;
        RECT 133.425 150.230 138.725 150.370 ;
        RECT 133.425 150.185 133.715 150.230 ;
        RECT 135.315 150.185 135.605 150.230 ;
        RECT 138.435 150.185 138.725 150.230 ;
        RECT 141.740 150.370 142.060 150.430 ;
        RECT 142.215 150.370 142.505 150.415 ;
        RECT 141.740 150.230 142.505 150.370 ;
        RECT 141.740 150.170 142.060 150.230 ;
        RECT 142.215 150.185 142.505 150.230 ;
        RECT 119.290 149.890 128.630 150.030 ;
        RECT 131.175 150.030 131.465 150.075 ;
        RECT 142.660 150.030 142.980 150.090 ;
        RECT 131.175 149.890 142.980 150.030 ;
        RECT 115.995 149.845 116.285 149.890 ;
        RECT 117.820 149.830 118.140 149.890 ;
        RECT 126.100 149.830 126.420 149.890 ;
        RECT 131.175 149.845 131.465 149.890 ;
        RECT 142.660 149.830 142.980 149.890 ;
        RECT 2.750 149.210 158.230 149.690 ;
        RECT 16.175 149.010 16.465 149.055 ;
        RECT 2.450 148.870 16.465 149.010 ;
        RECT 16.175 148.825 16.465 148.870 ;
        RECT 18.920 148.810 19.240 149.070 ;
        RECT 24.440 149.010 24.760 149.070 ;
        RECT 24.440 148.870 27.430 149.010 ;
        RECT 24.440 148.810 24.760 148.870 ;
        RECT 5.085 148.670 5.375 148.715 ;
        RECT 6.975 148.670 7.265 148.715 ;
        RECT 10.095 148.670 10.385 148.715 ;
        RECT 13.415 148.670 13.705 148.715 ;
        RECT 5.085 148.530 10.385 148.670 ;
        RECT 5.085 148.485 5.375 148.530 ;
        RECT 6.975 148.485 7.265 148.530 ;
        RECT 10.095 148.485 10.385 148.530 ;
        RECT 10.730 148.530 13.705 148.670 ;
        RECT 6.040 148.330 6.360 148.390 ;
        RECT 10.730 148.330 10.870 148.530 ;
        RECT 13.415 148.485 13.705 148.530 ;
        RECT 13.860 148.670 14.180 148.730 ;
        RECT 14.780 148.670 15.100 148.730 ;
        RECT 19.010 148.670 19.150 148.810 ;
        RECT 13.860 148.530 15.100 148.670 ;
        RECT 13.860 148.470 14.180 148.530 ;
        RECT 14.780 148.470 15.100 148.530 ;
        RECT 18.550 148.530 19.150 148.670 ;
        RECT 23.980 148.670 24.300 148.730 ;
        RECT 27.290 148.670 27.430 148.870 ;
        RECT 28.595 148.825 28.885 149.055 ;
        RECT 29.500 149.010 29.820 149.070 ;
        RECT 31.815 149.010 32.105 149.055 ;
        RECT 29.500 148.870 32.105 149.010 ;
        RECT 28.670 148.670 28.810 148.825 ;
        RECT 29.500 148.810 29.820 148.870 ;
        RECT 31.815 148.825 32.105 148.870 ;
        RECT 32.735 149.010 33.025 149.055 ;
        RECT 33.640 149.010 33.960 149.070 ;
        RECT 32.735 148.870 33.960 149.010 ;
        RECT 32.735 148.825 33.025 148.870 ;
        RECT 33.640 148.810 33.960 148.870 ;
        RECT 35.020 149.010 35.340 149.070 ;
        RECT 46.520 149.010 46.840 149.070 ;
        RECT 48.375 149.010 48.665 149.055 ;
        RECT 51.120 149.010 51.440 149.070 ;
        RECT 35.020 148.870 47.210 149.010 ;
        RECT 35.020 148.810 35.340 148.870 ;
        RECT 46.520 148.810 46.840 148.870 ;
        RECT 33.180 148.670 33.500 148.730 ;
        RECT 39.160 148.670 39.480 148.730 ;
        RECT 41.000 148.670 41.320 148.730 ;
        RECT 42.395 148.670 42.685 148.715 ;
        RECT 23.980 148.530 26.050 148.670 ;
        RECT 27.290 148.530 27.890 148.670 ;
        RECT 28.670 148.530 32.950 148.670 ;
        RECT 18.550 148.375 18.690 148.530 ;
        RECT 23.980 148.470 24.300 148.530 ;
        RECT 6.040 148.190 10.870 148.330 ;
        RECT 12.955 148.330 13.245 148.375 ;
        RECT 12.955 148.190 18.230 148.330 ;
        RECT 6.040 148.130 6.360 148.190 ;
        RECT 12.955 148.145 13.245 148.190 ;
        RECT 4.200 147.790 4.520 148.050 ;
        RECT 4.680 147.990 4.970 148.035 ;
        RECT 6.515 147.990 6.805 148.035 ;
        RECT 10.095 147.990 10.385 148.035 ;
        RECT 4.680 147.850 10.385 147.990 ;
        RECT 4.680 147.805 4.970 147.850 ;
        RECT 6.515 147.805 6.805 147.850 ;
        RECT 10.095 147.805 10.385 147.850 ;
        RECT 11.100 148.010 11.420 148.050 ;
        RECT 11.100 147.790 11.465 148.010 ;
        RECT 14.320 147.790 14.640 148.050 ;
        RECT 18.090 147.990 18.230 148.190 ;
        RECT 18.475 148.145 18.765 148.375 ;
        RECT 18.920 148.130 19.240 148.390 ;
        RECT 24.070 148.190 25.525 148.330 ;
        RECT 24.070 148.050 24.210 148.190 ;
        RECT 20.760 147.990 21.080 148.050 ;
        RECT 23.075 147.990 23.365 148.035 ;
        RECT 18.090 147.850 23.365 147.990 ;
        RECT 20.760 147.790 21.080 147.850 ;
        RECT 23.075 147.805 23.365 147.850 ;
        RECT 23.980 147.790 24.300 148.050 ;
        RECT 24.915 147.970 25.205 148.035 ;
        RECT 25.385 147.970 25.525 148.190 ;
        RECT 25.910 148.035 26.050 148.530 ;
        RECT 27.200 148.130 27.520 148.390 ;
        RECT 27.750 148.330 27.890 148.530 ;
        RECT 27.750 148.190 32.490 148.330 ;
        RECT 24.915 147.830 25.525 147.970 ;
        RECT 24.915 147.805 25.205 147.830 ;
        RECT 25.835 147.805 26.125 148.035 ;
        RECT 27.290 147.990 27.430 148.130 ;
        RECT 27.750 148.035 27.890 148.190 ;
        RECT 26.830 147.850 27.430 147.990 ;
        RECT 11.175 147.695 11.465 147.790 ;
        RECT 5.595 147.465 5.885 147.695 ;
        RECT 7.875 147.650 8.525 147.695 ;
        RECT 11.175 147.650 11.765 147.695 ;
        RECT 7.875 147.510 11.765 147.650 ;
        RECT 7.875 147.465 8.525 147.510 ;
        RECT 11.475 147.465 11.765 147.510 ;
        RECT 13.860 147.650 14.180 147.710 ;
        RECT 22.600 147.650 22.920 147.710 ;
        RECT 24.440 147.650 24.760 147.710 ;
        RECT 26.830 147.695 26.970 147.850 ;
        RECT 27.675 147.805 27.965 148.035 ;
        RECT 29.040 147.790 29.360 148.050 ;
        RECT 30.420 147.790 30.740 148.050 ;
        RECT 30.880 147.790 31.200 148.050 ;
        RECT 13.860 147.510 20.530 147.650 ;
        RECT 4.660 147.310 4.980 147.370 ;
        RECT 5.670 147.310 5.810 147.465 ;
        RECT 13.860 147.450 14.180 147.510 ;
        RECT 4.660 147.170 5.810 147.310 ;
        RECT 12.940 147.310 13.260 147.370 ;
        RECT 18.015 147.310 18.305 147.355 ;
        RECT 19.380 147.310 19.700 147.370 ;
        RECT 20.390 147.355 20.530 147.510 ;
        RECT 22.600 147.510 26.510 147.650 ;
        RECT 22.600 147.450 22.920 147.510 ;
        RECT 24.440 147.450 24.760 147.510 ;
        RECT 12.940 147.170 19.700 147.310 ;
        RECT 4.660 147.110 4.980 147.170 ;
        RECT 12.940 147.110 13.260 147.170 ;
        RECT 18.015 147.125 18.305 147.170 ;
        RECT 19.380 147.110 19.700 147.170 ;
        RECT 20.315 147.125 20.605 147.355 ;
        RECT 23.520 147.310 23.840 147.370 ;
        RECT 23.995 147.310 24.285 147.355 ;
        RECT 23.520 147.170 24.285 147.310 ;
        RECT 26.370 147.310 26.510 147.510 ;
        RECT 26.755 147.465 27.045 147.695 ;
        RECT 27.195 147.650 27.485 147.695 ;
        RECT 28.120 147.650 28.440 147.710 ;
        RECT 27.195 147.510 28.440 147.650 ;
        RECT 27.195 147.465 27.485 147.510 ;
        RECT 28.120 147.450 28.440 147.510 ;
        RECT 29.975 147.465 30.265 147.695 ;
        RECT 32.350 147.650 32.490 148.190 ;
        RECT 32.810 147.970 32.950 148.530 ;
        RECT 33.180 148.530 34.330 148.670 ;
        RECT 33.180 148.470 33.500 148.530 ;
        RECT 34.190 148.035 34.330 148.530 ;
        RECT 39.160 148.530 40.795 148.670 ;
        RECT 39.160 148.470 39.480 148.530 ;
        RECT 35.480 148.130 35.800 148.390 ;
        RECT 36.400 148.330 36.720 148.390 ;
        RECT 40.655 148.330 40.795 148.530 ;
        RECT 41.000 148.530 42.685 148.670 ;
        RECT 41.000 148.470 41.320 148.530 ;
        RECT 42.395 148.485 42.685 148.530 ;
        RECT 44.220 148.670 44.540 148.730 ;
        RECT 44.220 148.530 46.775 148.670 ;
        RECT 44.220 148.470 44.540 148.530 ;
        RECT 46.060 148.330 46.380 148.390 ;
        RECT 36.400 148.190 39.850 148.330 ;
        RECT 40.655 148.190 41.230 148.330 ;
        RECT 36.400 148.130 36.720 148.190 ;
        RECT 39.710 148.050 39.850 148.190 ;
        RECT 33.655 147.990 33.945 148.035 ;
        RECT 33.270 147.970 33.945 147.990 ;
        RECT 32.810 147.850 33.945 147.970 ;
        RECT 32.810 147.830 33.410 147.850 ;
        RECT 33.655 147.805 33.945 147.850 ;
        RECT 34.115 147.805 34.405 148.035 ;
        RECT 37.780 147.990 38.100 148.050 ;
        RECT 38.485 147.990 38.775 148.035 ;
        RECT 35.110 147.850 38.775 147.990 ;
        RECT 35.110 147.650 35.250 147.850 ;
        RECT 37.780 147.790 38.100 147.850 ;
        RECT 38.485 147.805 38.775 147.850 ;
        RECT 39.620 147.790 39.940 148.050 ;
        RECT 40.080 148.035 40.400 148.050 ;
        RECT 41.090 148.035 41.230 148.190 ;
        RECT 41.550 148.190 43.070 148.330 ;
        RECT 41.550 148.050 41.690 148.190 ;
        RECT 40.080 147.805 40.565 148.035 ;
        RECT 41.015 147.805 41.305 148.035 ;
        RECT 40.080 147.790 40.400 147.805 ;
        RECT 41.460 147.790 41.780 148.050 ;
        RECT 42.395 147.990 42.685 148.035 ;
        RECT 42.010 147.850 42.685 147.990 ;
        RECT 36.415 147.650 36.705 147.695 ;
        RECT 32.350 147.510 35.250 147.650 ;
        RECT 35.570 147.510 36.705 147.650 ;
        RECT 30.050 147.310 30.190 147.465 ;
        RECT 26.370 147.170 30.190 147.310 ;
        RECT 32.720 147.310 33.040 147.370 ;
        RECT 35.570 147.310 35.710 147.510 ;
        RECT 36.415 147.465 36.705 147.510 ;
        RECT 37.320 147.650 37.640 147.710 ;
        RECT 39.175 147.650 39.465 147.695 ;
        RECT 37.320 147.510 39.465 147.650 ;
        RECT 37.320 147.450 37.640 147.510 ;
        RECT 39.175 147.465 39.465 147.510 ;
        RECT 32.720 147.170 35.710 147.310 ;
        RECT 35.940 147.310 36.260 147.370 ;
        RECT 36.875 147.310 37.165 147.355 ;
        RECT 35.940 147.170 37.165 147.310 ;
        RECT 23.520 147.110 23.840 147.170 ;
        RECT 23.995 147.125 24.285 147.170 ;
        RECT 32.720 147.110 33.040 147.170 ;
        RECT 35.940 147.110 36.260 147.170 ;
        RECT 36.875 147.125 37.165 147.170 ;
        RECT 37.780 147.110 38.100 147.370 ;
        RECT 38.240 147.310 38.560 147.370 ;
        RECT 42.010 147.310 42.150 147.850 ;
        RECT 42.395 147.805 42.685 147.850 ;
        RECT 42.930 147.650 43.070 148.190 ;
        RECT 44.310 148.190 46.380 148.330 ;
        RECT 43.760 147.790 44.080 148.050 ;
        RECT 44.310 148.035 44.450 148.190 ;
        RECT 46.060 148.130 46.380 148.190 ;
        RECT 45.140 148.035 45.460 148.050 ;
        RECT 46.635 148.035 46.775 148.530 ;
        RECT 47.070 148.330 47.210 148.870 ;
        RECT 48.375 148.870 51.440 149.010 ;
        RECT 48.375 148.825 48.665 148.870 ;
        RECT 51.120 148.810 51.440 148.870 ;
        RECT 52.055 149.010 52.345 149.055 ;
        RECT 54.800 149.010 55.120 149.070 ;
        RECT 52.055 148.870 55.120 149.010 ;
        RECT 52.055 148.825 52.345 148.870 ;
        RECT 54.800 148.810 55.120 148.870 ;
        RECT 55.720 148.810 56.040 149.070 ;
        RECT 57.575 149.010 57.865 149.055 ;
        RECT 58.020 149.010 58.340 149.070 ;
        RECT 57.575 148.870 79.410 149.010 ;
        RECT 57.575 148.825 57.865 148.870 ;
        RECT 58.020 148.810 58.340 148.870 ;
        RECT 47.455 148.670 47.745 148.715 ;
        RECT 48.820 148.670 49.140 148.730 ;
        RECT 47.455 148.530 49.140 148.670 ;
        RECT 55.810 148.670 55.950 148.810 ;
        RECT 58.480 148.670 58.800 148.730 ;
        RECT 55.810 148.530 58.800 148.670 ;
        RECT 47.455 148.485 47.745 148.530 ;
        RECT 48.820 148.470 49.140 148.530 ;
        RECT 58.480 148.470 58.800 148.530 ;
        RECT 60.435 148.670 60.725 148.715 ;
        RECT 63.555 148.670 63.845 148.715 ;
        RECT 65.445 148.670 65.735 148.715 ;
        RECT 66.760 148.670 67.080 148.730 ;
        RECT 60.435 148.530 65.735 148.670 ;
        RECT 60.435 148.485 60.725 148.530 ;
        RECT 63.555 148.485 63.845 148.530 ;
        RECT 65.445 148.485 65.735 148.530 ;
        RECT 65.930 148.530 67.080 148.670 ;
        RECT 50.660 148.330 50.980 148.390 ;
        RECT 54.355 148.330 54.645 148.375 ;
        RECT 57.100 148.330 57.420 148.390 ;
        RECT 62.160 148.330 62.480 148.390 ;
        RECT 65.930 148.330 66.070 148.530 ;
        RECT 66.760 148.470 67.080 148.530 ;
        RECT 67.695 148.670 67.985 148.715 ;
        RECT 69.945 148.670 70.235 148.715 ;
        RECT 71.835 148.670 72.125 148.715 ;
        RECT 74.955 148.670 75.245 148.715 ;
        RECT 67.695 148.530 68.370 148.670 ;
        RECT 67.695 148.485 67.985 148.530 ;
        RECT 47.070 148.190 54.645 148.330 ;
        RECT 50.660 148.130 50.980 148.190 ;
        RECT 54.355 148.145 54.645 148.190 ;
        RECT 55.350 148.190 57.725 148.330 ;
        RECT 44.235 147.805 44.525 148.035 ;
        RECT 44.975 147.805 45.460 148.035 ;
        RECT 46.560 147.805 46.850 148.035 ;
        RECT 45.140 147.790 45.460 147.805 ;
        RECT 49.280 147.790 49.600 148.050 ;
        RECT 49.740 147.790 50.060 148.050 ;
        RECT 50.200 147.790 50.520 148.050 ;
        RECT 51.120 147.790 51.440 148.050 ;
        RECT 52.960 147.790 53.280 148.050 ;
        RECT 53.420 147.790 53.740 148.050 ;
        RECT 54.800 147.790 55.120 148.050 ;
        RECT 55.350 148.035 55.490 148.190 ;
        RECT 57.100 148.130 57.420 148.190 ;
        RECT 55.275 147.805 55.565 148.035 ;
        RECT 55.735 147.805 56.025 148.035 ;
        RECT 45.615 147.650 45.905 147.695 ;
        RECT 42.930 147.510 45.905 147.650 ;
        RECT 42.930 147.370 43.070 147.510 ;
        RECT 45.615 147.465 45.905 147.510 ;
        RECT 46.075 147.650 46.365 147.695 ;
        RECT 50.290 147.650 50.430 147.790 ;
        RECT 54.340 147.650 54.660 147.710 ;
        RECT 55.810 147.650 55.950 147.805 ;
        RECT 46.075 147.510 49.970 147.650 ;
        RECT 50.290 147.510 55.950 147.650 ;
        RECT 46.075 147.465 46.365 147.510 ;
        RECT 49.830 147.370 49.970 147.510 ;
        RECT 54.340 147.450 54.660 147.510 ;
        RECT 38.240 147.170 42.150 147.310 ;
        RECT 38.240 147.110 38.560 147.170 ;
        RECT 42.840 147.110 43.160 147.370 ;
        RECT 45.140 147.310 45.460 147.370 ;
        RECT 46.520 147.310 46.840 147.370 ;
        RECT 45.140 147.170 46.840 147.310 ;
        RECT 45.140 147.110 45.460 147.170 ;
        RECT 46.520 147.110 46.840 147.170 ;
        RECT 49.740 147.110 50.060 147.370 ;
        RECT 54.800 147.310 55.120 147.370 ;
        RECT 55.720 147.310 56.040 147.370 ;
        RECT 54.800 147.170 56.040 147.310 ;
        RECT 54.800 147.110 55.120 147.170 ;
        RECT 55.720 147.110 56.040 147.170 ;
        RECT 57.100 147.110 57.420 147.370 ;
        RECT 57.585 147.310 57.725 148.190 ;
        RECT 62.160 148.190 66.070 148.330 ;
        RECT 66.315 148.330 66.605 148.375 ;
        RECT 67.220 148.330 67.540 148.390 ;
        RECT 66.315 148.190 67.540 148.330 ;
        RECT 62.160 148.130 62.480 148.190 ;
        RECT 66.315 148.145 66.605 148.190 ;
        RECT 67.220 148.130 67.540 148.190 ;
        RECT 59.355 147.695 59.645 148.010 ;
        RECT 60.435 147.990 60.725 148.035 ;
        RECT 64.015 147.990 64.305 148.035 ;
        RECT 65.850 147.990 66.140 148.035 ;
        RECT 68.230 147.990 68.370 148.530 ;
        RECT 69.945 148.530 75.245 148.670 ;
        RECT 69.945 148.485 70.235 148.530 ;
        RECT 71.835 148.485 72.125 148.530 ;
        RECT 74.955 148.485 75.245 148.530 ;
        RECT 77.800 148.470 78.120 148.730 ;
        RECT 78.735 148.485 79.025 148.715 ;
        RECT 69.060 148.130 69.380 148.390 ;
        RECT 72.280 148.330 72.600 148.390 ;
        RECT 78.810 148.330 78.950 148.485 ;
        RECT 72.280 148.190 78.950 148.330 ;
        RECT 72.280 148.130 72.600 148.190 ;
        RECT 60.435 147.850 66.140 147.990 ;
        RECT 60.435 147.805 60.725 147.850 ;
        RECT 64.015 147.805 64.305 147.850 ;
        RECT 65.850 147.805 66.140 147.850 ;
        RECT 66.390 147.850 68.370 147.990 ;
        RECT 59.055 147.650 59.645 147.695 ;
        RECT 62.295 147.650 62.945 147.695 ;
        RECT 64.460 147.650 64.780 147.710 ;
        RECT 59.055 147.510 64.780 147.650 ;
        RECT 59.055 147.465 59.345 147.510 ;
        RECT 62.295 147.465 62.945 147.510 ;
        RECT 64.460 147.450 64.780 147.510 ;
        RECT 64.935 147.650 65.225 147.695 ;
        RECT 66.390 147.650 66.530 147.850 ;
        RECT 68.615 147.805 68.905 148.035 ;
        RECT 69.540 147.990 69.830 148.035 ;
        RECT 71.375 147.990 71.665 148.035 ;
        RECT 74.955 147.990 75.245 148.035 ;
        RECT 69.540 147.850 75.245 147.990 ;
        RECT 69.540 147.805 69.830 147.850 ;
        RECT 71.375 147.805 71.665 147.850 ;
        RECT 74.955 147.805 75.245 147.850 ;
        RECT 75.960 148.010 76.280 148.050 ;
        RECT 64.935 147.510 66.530 147.650 ;
        RECT 66.760 147.650 67.080 147.710 ;
        RECT 68.690 147.650 68.830 147.805 ;
        RECT 75.960 147.790 76.325 148.010 ;
        RECT 66.760 147.510 68.830 147.650 ;
        RECT 64.935 147.465 65.225 147.510 ;
        RECT 66.760 147.450 67.080 147.510 ;
        RECT 70.440 147.450 70.760 147.710 ;
        RECT 76.035 147.695 76.325 147.790 ;
        RECT 72.735 147.650 73.385 147.695 ;
        RECT 76.035 147.650 76.625 147.695 ;
        RECT 72.735 147.510 76.625 147.650 ;
        RECT 72.735 147.465 73.385 147.510 ;
        RECT 76.335 147.465 76.625 147.510 ;
        RECT 75.500 147.310 75.820 147.370 ;
        RECT 57.585 147.170 75.820 147.310 ;
        RECT 79.270 147.310 79.410 148.870 ;
        RECT 90.220 148.810 90.540 149.070 ;
        RECT 98.040 149.010 98.360 149.070 ;
        RECT 102.195 149.010 102.485 149.055 ;
        RECT 115.980 149.010 116.300 149.070 ;
        RECT 98.040 148.870 116.300 149.010 ;
        RECT 98.040 148.810 98.360 148.870 ;
        RECT 102.195 148.825 102.485 148.870 ;
        RECT 115.980 148.810 116.300 148.870 ;
        RECT 118.280 148.810 118.600 149.070 ;
        RECT 118.740 149.010 119.060 149.070 ;
        RECT 121.960 149.010 122.280 149.070 ;
        RECT 130.255 149.010 130.545 149.055 ;
        RECT 144.960 149.010 145.280 149.070 ;
        RECT 118.740 148.870 122.280 149.010 ;
        RECT 118.740 148.810 119.060 148.870 ;
        RECT 121.960 148.810 122.280 148.870 ;
        RECT 125.735 148.870 130.010 149.010 ;
        RECT 82.400 148.670 82.720 148.730 ;
        RECT 80.650 148.530 82.720 148.670 ;
        RECT 79.640 148.330 79.960 148.390 ;
        RECT 80.650 148.375 80.790 148.530 ;
        RECT 82.400 148.470 82.720 148.530 ;
        RECT 86.095 148.670 86.385 148.715 ;
        RECT 90.310 148.670 90.450 148.810 ;
        RECT 86.095 148.530 90.450 148.670 ;
        RECT 94.325 148.670 94.615 148.715 ;
        RECT 96.215 148.670 96.505 148.715 ;
        RECT 99.335 148.670 99.625 148.715 ;
        RECT 94.325 148.530 99.625 148.670 ;
        RECT 86.095 148.485 86.385 148.530 ;
        RECT 94.325 148.485 94.615 148.530 ;
        RECT 96.215 148.485 96.505 148.530 ;
        RECT 99.335 148.485 99.625 148.530 ;
        RECT 104.020 148.470 104.340 148.730 ;
        RECT 115.060 148.670 115.380 148.730 ;
        RECT 108.250 148.530 115.380 148.670 ;
        RECT 80.575 148.330 80.865 148.375 ;
        RECT 79.640 148.190 80.865 148.330 ;
        RECT 79.640 148.130 79.960 148.190 ;
        RECT 80.575 148.145 80.865 148.190 ;
        RECT 81.480 148.130 81.800 148.390 ;
        RECT 83.335 148.330 83.625 148.375 ;
        RECT 84.240 148.330 84.560 148.390 ;
        RECT 83.335 148.190 84.560 148.330 ;
        RECT 83.335 148.145 83.625 148.190 ;
        RECT 84.240 148.130 84.560 148.190 ;
        RECT 89.300 148.330 89.620 148.390 ;
        RECT 91.155 148.330 91.445 148.375 ;
        RECT 89.300 148.190 91.445 148.330 ;
        RECT 89.300 148.130 89.620 148.190 ;
        RECT 91.155 148.145 91.445 148.190 ;
        RECT 93.440 148.130 93.760 148.390 ;
        RECT 94.820 148.330 95.140 148.390 ;
        RECT 94.820 148.190 103.790 148.330 ;
        RECT 94.820 148.130 95.140 148.190 ;
        RECT 88.380 147.990 88.700 148.050 ;
        RECT 88.855 147.990 89.145 148.035 ;
        RECT 81.110 147.850 89.145 147.990 ;
        RECT 81.110 147.695 81.250 147.850 ;
        RECT 88.380 147.790 88.700 147.850 ;
        RECT 88.855 147.805 89.145 147.850 ;
        RECT 90.680 147.790 91.000 148.050 ;
        RECT 91.600 147.790 91.920 148.050 ;
        RECT 92.075 147.990 92.365 148.035 ;
        RECT 92.520 147.990 92.840 148.050 ;
        RECT 92.075 147.850 92.840 147.990 ;
        RECT 92.075 147.805 92.365 147.850 ;
        RECT 92.520 147.790 92.840 147.850 ;
        RECT 93.920 147.990 94.210 148.035 ;
        RECT 95.755 147.990 96.045 148.035 ;
        RECT 99.335 147.990 99.625 148.035 ;
        RECT 93.920 147.850 99.625 147.990 ;
        RECT 93.920 147.805 94.210 147.850 ;
        RECT 95.755 147.805 96.045 147.850 ;
        RECT 99.335 147.805 99.625 147.850 ;
        RECT 100.340 148.010 100.660 148.050 ;
        RECT 100.340 147.790 100.705 148.010 ;
        RECT 100.415 147.695 100.705 147.790 ;
        RECT 81.035 147.465 81.325 147.695 ;
        RECT 89.775 147.650 90.065 147.695 ;
        RECT 94.835 147.650 95.125 147.695 ;
        RECT 81.570 147.510 88.610 147.650 ;
        RECT 81.570 147.310 81.710 147.510 ;
        RECT 79.270 147.170 81.710 147.310 ;
        RECT 75.500 147.110 75.820 147.170 ;
        RECT 83.780 147.110 84.100 147.370 ;
        RECT 84.255 147.310 84.545 147.355 ;
        RECT 84.700 147.310 85.020 147.370 ;
        RECT 87.935 147.310 88.225 147.355 ;
        RECT 84.255 147.170 88.225 147.310 ;
        RECT 88.470 147.310 88.610 147.510 ;
        RECT 89.775 147.510 95.125 147.650 ;
        RECT 89.775 147.465 90.065 147.510 ;
        RECT 94.835 147.465 95.125 147.510 ;
        RECT 97.115 147.650 97.765 147.695 ;
        RECT 100.415 147.650 101.005 147.695 ;
        RECT 97.115 147.510 101.005 147.650 ;
        RECT 103.650 147.650 103.790 148.190 ;
        RECT 104.110 147.990 104.250 148.470 ;
        RECT 105.875 148.330 106.165 148.375 ;
        RECT 107.700 148.330 108.020 148.390 ;
        RECT 105.875 148.190 108.020 148.330 ;
        RECT 105.875 148.145 106.165 148.190 ;
        RECT 107.700 148.130 108.020 148.190 ;
        RECT 105.415 147.990 105.705 148.035 ;
        RECT 104.110 147.850 105.705 147.990 ;
        RECT 105.415 147.805 105.705 147.850 ;
        RECT 106.320 147.990 106.640 148.050 ;
        RECT 107.255 147.990 107.545 148.035 ;
        RECT 108.250 147.990 108.390 148.530 ;
        RECT 115.060 148.470 115.380 148.530 ;
        RECT 115.535 148.485 115.825 148.715 ;
        RECT 118.370 148.670 118.510 148.810 ;
        RECT 118.370 148.530 120.810 148.670 ;
        RECT 113.235 148.330 113.525 148.375 ;
        RECT 110.320 148.190 113.525 148.330 ;
        RECT 106.320 147.850 108.390 147.990 ;
        RECT 106.320 147.790 106.640 147.850 ;
        RECT 107.255 147.805 107.545 147.850 ;
        RECT 109.540 147.790 109.860 148.050 ;
        RECT 108.160 147.650 108.480 147.710 ;
        RECT 103.650 147.510 108.480 147.650 ;
        RECT 97.115 147.465 97.765 147.510 ;
        RECT 100.715 147.465 101.005 147.510 ;
        RECT 108.160 147.450 108.480 147.510 ;
        RECT 110.320 147.310 110.460 148.190 ;
        RECT 113.235 148.145 113.525 148.190 ;
        RECT 115.610 148.330 115.750 148.485 ;
        RECT 115.610 148.190 118.510 148.330 ;
        RECT 110.935 147.990 111.225 148.035 ;
        RECT 111.380 147.990 111.700 148.050 ;
        RECT 110.935 147.850 111.700 147.990 ;
        RECT 110.935 147.805 111.225 147.850 ;
        RECT 111.380 147.790 111.700 147.850 ;
        RECT 111.855 147.805 112.145 148.035 ;
        RECT 112.300 147.990 112.620 148.050 ;
        RECT 112.775 147.990 113.065 148.035 ;
        RECT 112.300 147.850 113.065 147.990 ;
        RECT 88.470 147.170 110.460 147.310 ;
        RECT 84.255 147.125 84.545 147.170 ;
        RECT 84.700 147.110 85.020 147.170 ;
        RECT 87.935 147.125 88.225 147.170 ;
        RECT 111.380 147.110 111.700 147.370 ;
        RECT 111.930 147.310 112.070 147.805 ;
        RECT 112.300 147.790 112.620 147.850 ;
        RECT 112.775 147.805 113.065 147.850 ;
        RECT 113.220 147.450 113.540 147.710 ;
        RECT 112.760 147.310 113.080 147.370 ;
        RECT 115.610 147.310 115.750 148.190 ;
        RECT 115.980 147.990 116.300 148.050 ;
        RECT 118.370 148.035 118.510 148.190 ;
        RECT 119.290 148.190 120.350 148.330 ;
        RECT 119.290 148.050 119.430 148.190 ;
        RECT 117.375 147.990 117.665 148.035 ;
        RECT 115.980 147.850 117.665 147.990 ;
        RECT 115.980 147.790 116.300 147.850 ;
        RECT 117.375 147.805 117.665 147.850 ;
        RECT 118.295 147.990 118.585 148.035 ;
        RECT 118.740 147.990 119.060 148.050 ;
        RECT 118.295 147.850 119.060 147.990 ;
        RECT 118.295 147.805 118.585 147.850 ;
        RECT 118.740 147.790 119.060 147.850 ;
        RECT 119.200 147.790 119.520 148.050 ;
        RECT 120.210 148.035 120.350 148.190 ;
        RECT 120.670 148.035 120.810 148.530 ;
        RECT 121.040 148.470 121.360 148.730 ;
        RECT 121.130 148.330 121.270 148.470 ;
        RECT 125.735 148.330 125.875 148.870 ;
        RECT 126.115 148.670 126.405 148.715 ;
        RECT 128.860 148.670 129.180 148.730 ;
        RECT 126.115 148.530 129.180 148.670 ;
        RECT 129.870 148.670 130.010 148.870 ;
        RECT 130.255 148.870 145.280 149.010 ;
        RECT 130.255 148.825 130.545 148.870 ;
        RECT 144.960 148.810 145.280 148.870 ;
        RECT 131.620 148.670 131.940 148.730 ;
        RECT 129.870 148.530 131.940 148.670 ;
        RECT 126.115 148.485 126.405 148.530 ;
        RECT 128.860 148.470 129.180 148.530 ;
        RECT 131.620 148.470 131.940 148.530 ;
        RECT 134.805 148.670 135.095 148.715 ;
        RECT 136.695 148.670 136.985 148.715 ;
        RECT 139.815 148.670 140.105 148.715 ;
        RECT 134.805 148.530 140.105 148.670 ;
        RECT 134.805 148.485 135.095 148.530 ;
        RECT 136.695 148.485 136.985 148.530 ;
        RECT 139.815 148.485 140.105 148.530 ;
        RECT 141.280 148.470 141.600 148.730 ;
        RECT 121.130 148.190 125.875 148.330 ;
        RECT 119.675 147.805 119.965 148.035 ;
        RECT 120.135 147.805 120.425 148.035 ;
        RECT 120.670 147.850 120.980 148.035 ;
        RECT 121.130 147.990 121.270 148.190 ;
        RECT 121.515 147.990 121.805 148.035 ;
        RECT 122.895 147.990 123.185 148.035 ;
        RECT 121.130 147.850 121.805 147.990 ;
        RECT 120.690 147.805 120.980 147.850 ;
        RECT 121.515 147.805 121.805 147.850 ;
        RECT 122.050 147.850 123.185 147.990 ;
        RECT 119.750 147.650 119.890 147.805 ;
        RECT 122.050 147.650 122.190 147.850 ;
        RECT 122.895 147.805 123.185 147.850 ;
        RECT 123.340 147.990 123.660 148.050 ;
        RECT 124.350 148.035 124.490 148.190 ;
        RECT 127.480 148.130 127.800 148.390 ;
        RECT 132.540 148.330 132.860 148.390 ;
        RECT 133.920 148.330 134.240 148.390 ;
        RECT 132.540 148.190 134.240 148.330 ;
        RECT 132.540 148.130 132.860 148.190 ;
        RECT 133.920 148.130 134.240 148.190 ;
        RECT 123.815 147.990 124.105 148.035 ;
        RECT 123.340 147.850 124.105 147.990 ;
        RECT 123.340 147.790 123.660 147.850 ;
        RECT 123.815 147.805 124.105 147.850 ;
        RECT 124.275 147.805 124.565 148.035 ;
        RECT 124.720 147.790 125.040 148.050 ;
        RECT 131.160 147.990 131.480 148.050 ;
        RECT 131.635 147.990 131.925 148.035 ;
        RECT 127.595 147.850 131.925 147.990 ;
        RECT 117.450 147.510 122.190 147.650 ;
        RECT 117.450 147.370 117.590 147.510 ;
        RECT 111.930 147.170 115.750 147.310 ;
        RECT 112.760 147.110 113.080 147.170 ;
        RECT 117.360 147.110 117.680 147.370 ;
        RECT 117.835 147.310 118.125 147.355 ;
        RECT 120.580 147.310 120.900 147.370 ;
        RECT 117.835 147.170 120.900 147.310 ;
        RECT 122.050 147.310 122.190 147.510 ;
        RECT 122.435 147.650 122.725 147.695 ;
        RECT 126.560 147.650 126.880 147.710 ;
        RECT 122.435 147.510 126.880 147.650 ;
        RECT 122.435 147.465 122.725 147.510 ;
        RECT 126.560 147.450 126.880 147.510 ;
        RECT 126.100 147.310 126.420 147.370 ;
        RECT 127.595 147.310 127.735 147.850 ;
        RECT 131.160 147.790 131.480 147.850 ;
        RECT 131.635 147.805 131.925 147.850 ;
        RECT 132.095 147.990 132.385 148.035 ;
        RECT 134.400 147.990 134.690 148.035 ;
        RECT 136.235 147.990 136.525 148.035 ;
        RECT 139.815 147.990 140.105 148.035 ;
        RECT 132.095 147.850 133.690 147.990 ;
        RECT 132.095 147.805 132.385 147.850 ;
        RECT 133.550 147.710 133.690 147.850 ;
        RECT 134.400 147.850 140.105 147.990 ;
        RECT 134.400 147.805 134.690 147.850 ;
        RECT 136.235 147.805 136.525 147.850 ;
        RECT 139.815 147.805 140.105 147.850 ;
        RECT 140.895 147.990 141.185 148.010 ;
        RECT 141.370 147.990 141.510 148.470 ;
        RECT 140.895 147.850 141.510 147.990 ;
        RECT 133.015 147.650 133.305 147.695 ;
        RECT 130.790 147.510 133.305 147.650 ;
        RECT 130.790 147.370 130.930 147.510 ;
        RECT 133.015 147.465 133.305 147.510 ;
        RECT 133.460 147.450 133.780 147.710 ;
        RECT 140.895 147.695 141.185 147.850 ;
        RECT 135.315 147.465 135.605 147.695 ;
        RECT 137.595 147.650 138.245 147.695 ;
        RECT 140.895 147.650 141.485 147.695 ;
        RECT 137.595 147.510 141.485 147.650 ;
        RECT 137.595 147.465 138.245 147.510 ;
        RECT 141.195 147.465 141.485 147.510 ;
        RECT 122.050 147.170 127.735 147.310 ;
        RECT 117.835 147.125 118.125 147.170 ;
        RECT 120.580 147.110 120.900 147.170 ;
        RECT 126.100 147.110 126.420 147.170 ;
        RECT 127.940 147.110 128.260 147.370 ;
        RECT 128.400 147.110 128.720 147.370 ;
        RECT 130.700 147.110 131.020 147.370 ;
        RECT 132.555 147.310 132.845 147.355 ;
        RECT 134.380 147.310 134.700 147.370 ;
        RECT 132.555 147.170 134.700 147.310 ;
        RECT 135.390 147.310 135.530 147.465 ;
        RECT 144.040 147.450 144.360 147.710 ;
        RECT 139.900 147.310 140.220 147.370 ;
        RECT 135.390 147.170 140.220 147.310 ;
        RECT 132.555 147.125 132.845 147.170 ;
        RECT 134.380 147.110 134.700 147.170 ;
        RECT 139.900 147.110 140.220 147.170 ;
        RECT 2.750 146.490 159.030 146.970 ;
        RECT 8.340 146.290 8.660 146.350 ;
        RECT 17.080 146.290 17.400 146.350 ;
        RECT 19.840 146.290 20.160 146.350 ;
        RECT 23.075 146.290 23.365 146.335 ;
        RECT 26.280 146.290 26.600 146.350 ;
        RECT 8.340 146.150 17.770 146.290 ;
        RECT 8.340 146.090 8.660 146.150 ;
        RECT 17.080 146.090 17.400 146.150 ;
        RECT 8.430 145.950 8.570 146.090 ;
        RECT 6.130 145.810 8.570 145.950 ;
        RECT 10.195 145.950 10.485 145.995 ;
        RECT 12.480 145.950 12.800 146.010 ;
        RECT 10.195 145.810 12.800 145.950 ;
        RECT 5.120 145.410 5.440 145.670 ;
        RECT 6.130 145.655 6.270 145.810 ;
        RECT 10.195 145.765 10.485 145.810 ;
        RECT 12.480 145.750 12.800 145.810 ;
        RECT 17.630 145.730 17.770 146.150 ;
        RECT 19.840 146.150 22.830 146.290 ;
        RECT 19.840 146.090 20.160 146.150 ;
        RECT 22.690 145.950 22.830 146.150 ;
        RECT 23.075 146.150 26.600 146.290 ;
        RECT 23.075 146.105 23.365 146.150 ;
        RECT 26.280 146.090 26.600 146.150 ;
        RECT 27.660 146.290 27.980 146.350 ;
        RECT 32.720 146.290 33.040 146.350 ;
        RECT 27.660 146.150 33.040 146.290 ;
        RECT 27.660 146.090 27.980 146.150 ;
        RECT 32.720 146.090 33.040 146.150 ;
        RECT 36.400 146.290 36.720 146.350 ;
        RECT 37.320 146.290 37.640 146.350 ;
        RECT 36.400 146.150 37.640 146.290 ;
        RECT 36.400 146.090 36.720 146.150 ;
        RECT 37.320 146.090 37.640 146.150 ;
        RECT 37.780 146.290 38.100 146.350 ;
        RECT 50.200 146.290 50.520 146.350 ;
        RECT 37.780 146.150 50.520 146.290 ;
        RECT 37.780 146.090 38.100 146.150 ;
        RECT 50.200 146.090 50.520 146.150 ;
        RECT 52.040 146.090 52.360 146.350 ;
        RECT 56.180 146.090 56.500 146.350 ;
        RECT 57.100 146.090 57.420 146.350 ;
        RECT 58.020 146.090 58.340 146.350 ;
        RECT 58.495 146.290 58.785 146.335 ;
        RECT 58.940 146.290 59.260 146.350 ;
        RECT 59.860 146.290 60.180 146.350 ;
        RECT 58.495 146.150 60.180 146.290 ;
        RECT 58.495 146.105 58.785 146.150 ;
        RECT 58.940 146.090 59.260 146.150 ;
        RECT 59.860 146.090 60.180 146.150 ;
        RECT 60.335 146.290 60.625 146.335 ;
        RECT 62.160 146.290 62.480 146.350 ;
        RECT 67.220 146.290 67.540 146.350 ;
        RECT 60.335 146.150 62.480 146.290 ;
        RECT 60.335 146.105 60.625 146.150 ;
        RECT 62.160 146.090 62.480 146.150 ;
        RECT 62.710 146.150 67.540 146.290 ;
        RECT 29.040 145.950 29.360 146.010 ;
        RECT 40.095 145.950 40.385 145.995 ;
        RECT 40.540 145.950 40.860 146.010 ;
        RECT 22.690 145.810 26.970 145.950 ;
        RECT 6.055 145.425 6.345 145.655 ;
        RECT 6.515 145.610 6.805 145.655 ;
        RECT 6.960 145.610 7.280 145.670 ;
        RECT 6.515 145.470 7.280 145.610 ;
        RECT 6.515 145.425 6.805 145.470 ;
        RECT 6.960 145.410 7.280 145.470 ;
        RECT 7.420 145.410 7.740 145.670 ;
        RECT 7.880 145.410 8.200 145.670 ;
        RECT 10.655 145.610 10.945 145.655 ;
        RECT 13.860 145.610 14.180 145.670 ;
        RECT 10.655 145.470 14.180 145.610 ;
        RECT 10.655 145.425 10.945 145.470 ;
        RECT 13.860 145.410 14.180 145.470 ;
        RECT 14.320 145.410 14.640 145.670 ;
        RECT 17.080 145.410 17.400 145.670 ;
        RECT 17.630 145.655 18.230 145.730 ;
        RECT 17.630 145.590 18.305 145.655 ;
        RECT 18.015 145.425 18.305 145.590 ;
        RECT 18.475 145.425 18.765 145.655 ;
        RECT 18.935 145.425 19.225 145.655 ;
        RECT 20.315 145.610 20.605 145.655 ;
        RECT 19.470 145.470 20.605 145.610 ;
        RECT 7.510 145.270 7.650 145.410 ;
        RECT 7.510 145.130 11.330 145.270 ;
        RECT 8.340 144.730 8.660 144.990 ;
        RECT 11.190 144.930 11.330 145.130 ;
        RECT 11.560 145.070 11.880 145.330 ;
        RECT 14.780 145.070 15.100 145.330 ;
        RECT 15.240 145.070 15.560 145.330 ;
        RECT 15.700 145.270 16.020 145.330 ;
        RECT 18.550 145.270 18.690 145.425 ;
        RECT 15.700 145.130 18.690 145.270 ;
        RECT 15.700 145.070 16.020 145.130 ;
        RECT 18.000 144.930 18.320 144.990 ;
        RECT 19.010 144.930 19.150 145.425 ;
        RECT 11.190 144.790 17.770 144.930 ;
        RECT 5.120 144.590 5.440 144.650 ;
        RECT 12.495 144.590 12.785 144.635 ;
        RECT 5.120 144.450 12.785 144.590 ;
        RECT 17.630 144.590 17.770 144.790 ;
        RECT 18.000 144.790 19.150 144.930 ;
        RECT 18.000 144.730 18.320 144.790 ;
        RECT 19.470 144.590 19.610 145.470 ;
        RECT 20.315 145.425 20.605 145.470 ;
        RECT 20.775 145.425 21.065 145.655 ;
        RECT 21.695 145.425 21.985 145.655 ;
        RECT 22.155 145.610 22.445 145.655 ;
        RECT 22.155 145.470 22.830 145.610 ;
        RECT 22.155 145.425 22.445 145.470 ;
        RECT 20.850 145.270 20.990 145.425 ;
        RECT 19.930 145.130 20.990 145.270 ;
        RECT 19.930 144.975 20.070 145.130 ;
        RECT 19.855 144.745 20.145 144.975 ;
        RECT 21.770 144.930 21.910 145.425 ;
        RECT 22.690 145.330 22.830 145.470 ;
        RECT 23.535 145.425 23.825 145.655 ;
        RECT 24.900 145.610 25.220 145.670 ;
        RECT 25.375 145.610 25.665 145.655 ;
        RECT 24.900 145.470 25.665 145.610 ;
        RECT 22.600 145.070 22.920 145.330 ;
        RECT 23.610 145.270 23.750 145.425 ;
        RECT 24.900 145.410 25.220 145.470 ;
        RECT 25.375 145.425 25.665 145.470 ;
        RECT 26.280 145.410 26.600 145.670 ;
        RECT 26.830 145.655 26.970 145.810 ;
        RECT 29.040 145.810 31.570 145.950 ;
        RECT 29.040 145.750 29.360 145.810 ;
        RECT 26.755 145.425 27.045 145.655 ;
        RECT 30.895 145.425 31.185 145.655 ;
        RECT 31.430 145.610 31.570 145.810 ;
        RECT 40.095 145.810 40.860 145.950 ;
        RECT 40.095 145.765 40.385 145.810 ;
        RECT 40.540 145.750 40.860 145.810 ;
        RECT 42.375 145.950 43.025 145.995 ;
        RECT 45.975 145.950 46.265 145.995 ;
        RECT 52.130 145.950 52.270 146.090 ;
        RECT 56.270 145.950 56.410 146.090 ;
        RECT 42.375 145.810 46.265 145.950 ;
        RECT 42.375 145.765 43.025 145.810 ;
        RECT 45.675 145.765 46.265 145.810 ;
        RECT 48.220 145.810 52.270 145.950 ;
        RECT 54.430 145.810 56.410 145.950 ;
        RECT 57.190 145.950 57.330 146.090 ;
        RECT 57.190 145.810 61.010 145.950 ;
        RECT 45.675 145.670 45.965 145.765 ;
        RECT 38.715 145.610 39.005 145.655 ;
        RECT 31.430 145.470 34.330 145.610 ;
        RECT 27.660 145.270 27.980 145.330 ;
        RECT 23.610 145.130 27.980 145.270 ;
        RECT 27.660 145.070 27.980 145.130 ;
        RECT 28.135 145.270 28.425 145.315 ;
        RECT 29.040 145.270 29.360 145.330 ;
        RECT 28.135 145.130 29.360 145.270 ;
        RECT 28.135 145.085 28.425 145.130 ;
        RECT 29.040 145.070 29.360 145.130 ;
        RECT 23.980 144.930 24.300 144.990 ;
        RECT 21.770 144.790 24.300 144.930 ;
        RECT 23.980 144.730 24.300 144.790 ;
        RECT 24.455 144.930 24.745 144.975 ;
        RECT 27.200 144.930 27.520 144.990 ;
        RECT 24.455 144.790 27.520 144.930 ;
        RECT 24.455 144.745 24.745 144.790 ;
        RECT 27.200 144.730 27.520 144.790 ;
        RECT 28.580 144.730 28.900 144.990 ;
        RECT 30.970 144.930 31.110 145.425 ;
        RECT 34.190 145.330 34.330 145.470 ;
        RECT 35.110 145.470 39.005 145.610 ;
        RECT 34.100 145.070 34.420 145.330 ;
        RECT 34.560 145.270 34.880 145.330 ;
        RECT 35.110 145.270 35.250 145.470 ;
        RECT 38.715 145.425 39.005 145.470 ;
        RECT 39.180 145.610 39.470 145.655 ;
        RECT 41.015 145.610 41.305 145.655 ;
        RECT 44.595 145.610 44.885 145.655 ;
        RECT 39.180 145.470 44.885 145.610 ;
        RECT 39.180 145.425 39.470 145.470 ;
        RECT 41.015 145.425 41.305 145.470 ;
        RECT 44.595 145.425 44.885 145.470 ;
        RECT 45.600 145.450 45.965 145.670 ;
        RECT 48.220 145.610 48.360 145.810 ;
        RECT 46.150 145.470 48.360 145.610 ;
        RECT 48.820 145.610 49.140 145.670 ;
        RECT 49.755 145.610 50.045 145.655 ;
        RECT 48.820 145.470 50.045 145.610 ;
        RECT 45.600 145.410 45.920 145.450 ;
        RECT 34.560 145.130 35.250 145.270 ;
        RECT 35.495 145.270 35.785 145.315 ;
        RECT 37.780 145.270 38.100 145.330 ;
        RECT 43.760 145.270 44.080 145.330 ;
        RECT 35.495 145.130 38.100 145.270 ;
        RECT 34.560 145.070 34.880 145.130 ;
        RECT 35.495 145.085 35.785 145.130 ;
        RECT 37.780 145.070 38.100 145.130 ;
        RECT 39.250 145.130 44.080 145.270 ;
        RECT 39.250 144.930 39.390 145.130 ;
        RECT 43.760 145.070 44.080 145.130 ;
        RECT 45.140 145.270 45.460 145.330 ;
        RECT 46.150 145.270 46.290 145.470 ;
        RECT 48.820 145.410 49.140 145.470 ;
        RECT 49.755 145.425 50.045 145.470 ;
        RECT 50.200 145.410 50.520 145.670 ;
        RECT 52.975 145.610 53.265 145.655 ;
        RECT 54.430 145.610 54.570 145.810 ;
        RECT 51.210 145.470 52.270 145.610 ;
        RECT 45.140 145.130 46.290 145.270 ;
        RECT 47.455 145.270 47.745 145.315 ;
        RECT 48.360 145.270 48.680 145.330 ;
        RECT 47.455 145.130 48.680 145.270 ;
        RECT 45.140 145.070 45.460 145.130 ;
        RECT 47.455 145.085 47.745 145.130 ;
        RECT 48.360 145.070 48.680 145.130 ;
        RECT 30.970 144.790 39.390 144.930 ;
        RECT 39.585 144.930 39.875 144.975 ;
        RECT 41.475 144.930 41.765 144.975 ;
        RECT 44.595 144.930 44.885 144.975 ;
        RECT 51.210 144.930 51.350 145.470 ;
        RECT 51.595 145.085 51.885 145.315 ;
        RECT 52.130 145.270 52.270 145.470 ;
        RECT 52.975 145.470 54.570 145.610 ;
        RECT 52.975 145.425 53.265 145.470 ;
        RECT 54.800 145.410 55.120 145.670 ;
        RECT 60.870 145.655 61.010 145.810 ;
        RECT 62.710 145.670 62.850 146.150 ;
        RECT 67.220 146.090 67.540 146.150 ;
        RECT 68.140 146.290 68.460 146.350 ;
        RECT 73.675 146.290 73.965 146.335 ;
        RECT 82.415 146.290 82.705 146.335 ;
        RECT 97.120 146.290 97.440 146.350 ;
        RECT 68.140 146.150 73.965 146.290 ;
        RECT 68.140 146.090 68.460 146.150 ;
        RECT 73.675 146.105 73.965 146.150 ;
        RECT 74.210 146.150 82.705 146.290 ;
        RECT 66.295 145.950 66.945 145.995 ;
        RECT 69.895 145.950 70.185 145.995 ;
        RECT 66.295 145.810 70.185 145.950 ;
        RECT 66.295 145.765 66.945 145.810 ;
        RECT 69.595 145.765 70.185 145.810 ;
        RECT 70.900 145.950 71.220 146.010 ;
        RECT 74.210 145.950 74.350 146.150 ;
        RECT 82.415 146.105 82.705 146.150 ;
        RECT 82.950 146.150 97.440 146.290 ;
        RECT 70.900 145.810 74.350 145.950 ;
        RECT 75.500 145.950 75.820 146.010 ;
        RECT 76.895 145.950 77.185 145.995 ;
        RECT 82.950 145.950 83.090 146.150 ;
        RECT 97.120 146.090 97.440 146.150 ;
        RECT 101.260 146.290 101.580 146.350 ;
        RECT 104.035 146.290 104.325 146.335 ;
        RECT 127.940 146.290 128.260 146.350 ;
        RECT 101.260 146.150 104.325 146.290 ;
        RECT 101.260 146.090 101.580 146.150 ;
        RECT 104.035 146.105 104.325 146.150 ;
        RECT 111.470 146.150 128.260 146.290 ;
        RECT 87.460 145.950 87.780 146.010 ;
        RECT 75.500 145.810 83.090 145.950 ;
        RECT 86.170 145.810 87.780 145.950 ;
        RECT 55.735 145.610 56.025 145.655 ;
        RECT 55.735 145.470 58.250 145.610 ;
        RECT 55.735 145.425 56.025 145.470 ;
        RECT 55.275 145.270 55.565 145.315 ;
        RECT 52.130 145.130 55.565 145.270 ;
        RECT 55.275 145.085 55.565 145.130 ;
        RECT 39.585 144.790 44.885 144.930 ;
        RECT 39.585 144.745 39.875 144.790 ;
        RECT 41.475 144.745 41.765 144.790 ;
        RECT 44.595 144.745 44.885 144.790 ;
        RECT 47.530 144.790 51.350 144.930 ;
        RECT 20.300 144.590 20.620 144.650 ;
        RECT 17.630 144.450 20.620 144.590 ;
        RECT 5.120 144.390 5.440 144.450 ;
        RECT 12.495 144.405 12.785 144.450 ;
        RECT 20.300 144.390 20.620 144.450 ;
        RECT 25.360 144.590 25.680 144.650 ;
        RECT 26.280 144.590 26.600 144.650 ;
        RECT 25.360 144.450 26.600 144.590 ;
        RECT 25.360 144.390 25.680 144.450 ;
        RECT 26.280 144.390 26.600 144.450 ;
        RECT 27.675 144.590 27.965 144.635 ;
        RECT 28.670 144.590 28.810 144.730 ;
        RECT 47.530 144.650 47.670 144.790 ;
        RECT 27.675 144.450 28.810 144.590 ;
        RECT 27.675 144.405 27.965 144.450 ;
        RECT 30.420 144.390 30.740 144.650 ;
        RECT 31.340 144.390 31.660 144.650 ;
        RECT 38.255 144.590 38.545 144.635 ;
        RECT 38.700 144.590 39.020 144.650 ;
        RECT 38.255 144.450 39.020 144.590 ;
        RECT 38.255 144.405 38.545 144.450 ;
        RECT 38.700 144.390 39.020 144.450 ;
        RECT 47.440 144.390 47.760 144.650 ;
        RECT 48.820 144.390 49.140 144.650 ;
        RECT 50.660 144.590 50.980 144.650 ;
        RECT 51.135 144.590 51.425 144.635 ;
        RECT 50.660 144.450 51.425 144.590 ;
        RECT 51.670 144.590 51.810 145.085 ;
        RECT 56.640 145.070 56.960 145.330 ;
        RECT 57.575 145.085 57.865 145.315 ;
        RECT 58.110 145.270 58.250 145.470 ;
        RECT 60.795 145.425 61.085 145.655 ;
        RECT 62.620 145.410 62.940 145.670 ;
        RECT 63.100 145.610 63.390 145.655 ;
        RECT 64.935 145.610 65.225 145.655 ;
        RECT 68.515 145.610 68.805 145.655 ;
        RECT 63.100 145.470 68.805 145.610 ;
        RECT 63.100 145.425 63.390 145.470 ;
        RECT 64.935 145.425 65.225 145.470 ;
        RECT 68.515 145.425 68.805 145.470 ;
        RECT 69.595 145.450 69.885 145.765 ;
        RECT 70.900 145.750 71.220 145.810 ;
        RECT 75.500 145.750 75.820 145.810 ;
        RECT 76.895 145.765 77.185 145.810 ;
        RECT 76.435 145.610 76.725 145.655 ;
        RECT 86.170 145.610 86.310 145.810 ;
        RECT 87.460 145.750 87.780 145.810 ;
        RECT 91.600 145.950 91.920 146.010 ;
        RECT 92.075 145.950 92.365 145.995 ;
        RECT 109.540 145.950 109.860 146.010 ;
        RECT 91.600 145.810 92.365 145.950 ;
        RECT 91.600 145.750 91.920 145.810 ;
        RECT 92.075 145.765 92.365 145.810 ;
        RECT 102.730 145.810 111.150 145.950 ;
        RECT 102.730 145.670 102.870 145.810 ;
        RECT 109.540 145.750 109.860 145.810 ;
        RECT 87.015 145.610 87.305 145.655 ;
        RECT 74.210 145.470 86.310 145.610 ;
        RECT 86.630 145.470 87.305 145.610 ;
        RECT 58.480 145.270 58.800 145.330 ;
        RECT 62.160 145.270 62.480 145.330 ;
        RECT 58.110 145.130 62.480 145.270 ;
        RECT 53.895 144.930 54.185 144.975 ;
        RECT 56.730 144.930 56.870 145.070 ;
        RECT 53.895 144.790 56.870 144.930 ;
        RECT 53.895 144.745 54.185 144.790 ;
        RECT 57.650 144.650 57.790 145.085 ;
        RECT 58.480 145.070 58.800 145.130 ;
        RECT 62.160 145.070 62.480 145.130 ;
        RECT 64.000 145.070 64.320 145.330 ;
        RECT 64.460 145.270 64.780 145.330 ;
        RECT 69.610 145.270 69.750 145.450 ;
        RECT 64.460 145.130 72.050 145.270 ;
        RECT 64.460 145.070 64.780 145.130 ;
        RECT 63.505 144.930 63.795 144.975 ;
        RECT 65.395 144.930 65.685 144.975 ;
        RECT 68.515 144.930 68.805 144.975 ;
        RECT 63.505 144.790 68.805 144.930 ;
        RECT 63.505 144.745 63.795 144.790 ;
        RECT 65.395 144.745 65.685 144.790 ;
        RECT 68.515 144.745 68.805 144.790 ;
        RECT 57.100 144.590 57.420 144.650 ;
        RECT 51.670 144.450 57.420 144.590 ;
        RECT 50.660 144.390 50.980 144.450 ;
        RECT 51.135 144.405 51.425 144.450 ;
        RECT 57.100 144.390 57.420 144.450 ;
        RECT 57.560 144.590 57.880 144.650 ;
        RECT 61.715 144.590 62.005 144.635 ;
        RECT 63.080 144.590 63.400 144.650 ;
        RECT 57.560 144.450 63.400 144.590 ;
        RECT 57.560 144.390 57.880 144.450 ;
        RECT 61.715 144.405 62.005 144.450 ;
        RECT 63.080 144.390 63.400 144.450 ;
        RECT 67.220 144.590 67.540 144.650 ;
        RECT 70.900 144.590 71.220 144.650 ;
        RECT 67.220 144.450 71.220 144.590 ;
        RECT 67.220 144.390 67.540 144.450 ;
        RECT 70.900 144.390 71.220 144.450 ;
        RECT 71.360 144.390 71.680 144.650 ;
        RECT 71.910 144.590 72.050 145.130 ;
        RECT 72.295 145.085 72.585 145.315 ;
        RECT 72.740 145.270 73.060 145.330 ;
        RECT 73.215 145.270 73.505 145.315 ;
        RECT 72.740 145.130 73.505 145.270 ;
        RECT 72.370 144.930 72.510 145.085 ;
        RECT 72.740 145.070 73.060 145.130 ;
        RECT 73.215 145.085 73.505 145.130 ;
        RECT 74.210 144.930 74.350 145.470 ;
        RECT 76.435 145.425 76.725 145.470 ;
        RECT 74.580 145.270 74.900 145.330 ;
        RECT 81.110 145.315 81.250 145.470 ;
        RECT 76.895 145.270 77.185 145.315 ;
        RECT 74.580 145.130 77.185 145.270 ;
        RECT 74.580 145.070 74.900 145.130 ;
        RECT 76.895 145.085 77.185 145.130 ;
        RECT 81.035 145.085 81.325 145.315 ;
        RECT 81.955 145.270 82.245 145.315 ;
        RECT 82.400 145.270 82.720 145.330 ;
        RECT 81.955 145.130 82.720 145.270 ;
        RECT 81.955 145.085 82.245 145.130 ;
        RECT 82.400 145.070 82.720 145.130 ;
        RECT 75.040 144.930 75.360 144.990 ;
        RECT 72.370 144.790 75.360 144.930 ;
        RECT 75.040 144.730 75.360 144.790 ;
        RECT 75.515 144.930 75.805 144.975 ;
        RECT 86.630 144.930 86.770 145.470 ;
        RECT 87.015 145.425 87.305 145.470 ;
        RECT 87.935 145.425 88.225 145.655 ;
        RECT 88.380 145.610 88.700 145.670 ;
        RECT 89.775 145.610 90.065 145.655 ;
        RECT 88.380 145.470 90.065 145.610 ;
        RECT 88.010 145.270 88.150 145.425 ;
        RECT 88.380 145.410 88.700 145.470 ;
        RECT 89.775 145.425 90.065 145.470 ;
        RECT 90.220 145.410 90.540 145.670 ;
        RECT 93.915 145.610 94.205 145.655 ;
        RECT 98.960 145.610 99.280 145.670 ;
        RECT 99.435 145.610 99.725 145.655 ;
        RECT 93.915 145.470 96.660 145.610 ;
        RECT 93.915 145.425 94.205 145.470 ;
        RECT 90.680 145.270 91.000 145.330 ;
        RECT 88.010 145.130 91.000 145.270 ;
        RECT 90.680 145.070 91.000 145.130 ;
        RECT 91.140 145.070 91.460 145.330 ;
        RECT 91.615 145.270 91.905 145.315 ;
        RECT 92.060 145.270 92.380 145.330 ;
        RECT 91.615 145.130 92.380 145.270 ;
        RECT 91.615 145.085 91.905 145.130 ;
        RECT 92.060 145.070 92.380 145.130 ;
        RECT 95.295 145.085 95.585 145.315 ;
        RECT 96.520 145.270 96.660 145.470 ;
        RECT 98.960 145.470 99.725 145.610 ;
        RECT 98.960 145.410 99.280 145.470 ;
        RECT 99.435 145.425 99.725 145.470 ;
        RECT 100.355 145.610 100.645 145.655 ;
        RECT 100.800 145.610 101.120 145.670 ;
        RECT 100.355 145.470 101.120 145.610 ;
        RECT 100.355 145.425 100.645 145.470 ;
        RECT 100.800 145.410 101.120 145.470 ;
        RECT 101.260 145.610 101.580 145.670 ;
        RECT 101.735 145.610 102.025 145.655 ;
        RECT 101.260 145.470 102.025 145.610 ;
        RECT 101.260 145.410 101.580 145.470 ;
        RECT 101.735 145.425 102.025 145.470 ;
        RECT 102.640 145.410 102.960 145.670 ;
        RECT 107.255 145.425 107.545 145.655 ;
        RECT 108.160 145.610 108.480 145.670 ;
        RECT 111.010 145.655 111.150 145.810 ;
        RECT 109.095 145.610 109.385 145.655 ;
        RECT 108.160 145.470 109.385 145.610 ;
        RECT 98.515 145.270 98.805 145.315 ;
        RECT 107.330 145.270 107.470 145.425 ;
        RECT 108.160 145.410 108.480 145.470 ;
        RECT 109.095 145.425 109.385 145.470 ;
        RECT 110.935 145.425 111.225 145.655 ;
        RECT 96.520 145.130 107.470 145.270 ;
        RECT 109.170 145.270 109.310 145.425 ;
        RECT 111.470 145.270 111.610 146.150 ;
        RECT 127.940 146.090 128.260 146.150 ;
        RECT 129.335 146.290 129.625 146.335 ;
        RECT 131.620 146.290 131.940 146.350 ;
        RECT 133.160 146.335 133.480 146.350 ;
        RECT 129.335 146.150 131.940 146.290 ;
        RECT 129.335 146.105 129.625 146.150 ;
        RECT 112.300 145.950 112.620 146.010 ;
        RECT 112.775 145.950 113.065 145.995 ;
        RECT 112.300 145.810 113.065 145.950 ;
        RECT 112.300 145.750 112.620 145.810 ;
        RECT 112.775 145.765 113.065 145.810 ;
        RECT 113.235 145.765 113.525 145.995 ;
        RECT 114.600 145.950 114.920 146.010 ;
        RECT 116.440 145.950 116.760 146.010 ;
        RECT 124.720 145.950 125.040 146.010 ;
        RECT 127.020 145.950 127.340 146.010 ;
        RECT 129.410 145.950 129.550 146.105 ;
        RECT 131.620 146.090 131.940 146.150 ;
        RECT 133.015 146.105 133.480 146.335 ;
        RECT 133.160 146.090 133.480 146.105 ;
        RECT 140.360 146.290 140.680 146.350 ;
        RECT 143.595 146.290 143.885 146.335 ;
        RECT 140.360 146.150 143.885 146.290 ;
        RECT 140.360 146.090 140.680 146.150 ;
        RECT 143.595 146.105 143.885 146.150 ;
        RECT 144.960 146.090 145.280 146.350 ;
        RECT 138.055 145.950 138.705 145.995 ;
        RECT 141.655 145.950 141.945 145.995 ;
        RECT 114.600 145.810 125.410 145.950 ;
        RECT 113.310 145.610 113.450 145.765 ;
        RECT 114.600 145.750 114.920 145.810 ;
        RECT 116.440 145.750 116.760 145.810 ;
        RECT 124.720 145.750 125.040 145.810 ;
        RECT 109.170 145.130 111.610 145.270 ;
        RECT 111.930 145.470 113.450 145.610 ;
        RECT 98.515 145.085 98.805 145.130 ;
        RECT 89.760 144.930 90.080 144.990 ;
        RECT 75.515 144.790 90.080 144.930 ;
        RECT 91.230 144.930 91.370 145.070 ;
        RECT 94.360 144.930 94.680 144.990 ;
        RECT 91.230 144.790 94.680 144.930 ;
        RECT 75.515 144.745 75.805 144.790 ;
        RECT 89.760 144.730 90.080 144.790 ;
        RECT 94.360 144.730 94.680 144.790 ;
        RECT 94.820 144.730 95.140 144.990 ;
        RECT 95.370 144.930 95.510 145.085 ;
        RECT 102.180 144.930 102.500 144.990 ;
        RECT 95.370 144.790 102.500 144.930 ;
        RECT 102.180 144.730 102.500 144.790 ;
        RECT 102.655 144.930 102.945 144.975 ;
        RECT 105.860 144.930 106.180 144.990 ;
        RECT 102.655 144.790 106.180 144.930 ;
        RECT 102.655 144.745 102.945 144.790 ;
        RECT 105.860 144.730 106.180 144.790 ;
        RECT 107.255 144.745 107.545 144.975 ;
        RECT 110.920 144.930 111.240 144.990 ;
        RECT 111.930 144.930 112.070 145.470 ;
        RECT 117.820 145.410 118.140 145.670 ;
        RECT 120.580 145.410 120.900 145.670 ;
        RECT 121.040 145.410 121.360 145.670 ;
        RECT 121.500 145.610 121.820 145.670 ;
        RECT 122.420 145.610 122.740 145.670 ;
        RECT 125.270 145.655 125.410 145.810 ;
        RECT 127.020 145.810 129.550 145.950 ;
        RECT 130.790 145.810 133.690 145.950 ;
        RECT 127.020 145.750 127.340 145.810 ;
        RECT 130.790 145.670 130.930 145.810 ;
        RECT 123.355 145.610 123.645 145.655 ;
        RECT 121.500 145.470 123.645 145.610 ;
        RECT 121.500 145.410 121.820 145.470 ;
        RECT 122.420 145.410 122.740 145.470 ;
        RECT 123.355 145.425 123.645 145.470 ;
        RECT 125.195 145.425 125.485 145.655 ;
        RECT 130.700 145.610 131.020 145.670 ;
        RECT 125.730 145.470 131.020 145.610 ;
        RECT 113.220 145.070 113.540 145.330 ;
        RECT 110.920 144.790 112.070 144.930 ;
        RECT 115.535 144.930 115.825 144.975 ;
        RECT 117.360 144.930 117.680 144.990 ;
        RECT 115.535 144.790 117.680 144.930 ;
        RECT 120.670 144.930 120.810 145.410 ;
        RECT 125.730 145.330 125.870 145.470 ;
        RECT 130.700 145.410 131.020 145.470 ;
        RECT 131.160 145.610 131.480 145.670 ;
        RECT 133.550 145.655 133.690 145.810 ;
        RECT 138.055 145.810 141.945 145.950 ;
        RECT 138.055 145.765 138.705 145.810 ;
        RECT 141.355 145.765 141.945 145.810 ;
        RECT 141.355 145.670 141.645 145.765 ;
        RECT 142.660 145.750 142.980 146.010 ;
        RECT 132.095 145.610 132.385 145.655 ;
        RECT 131.160 145.470 132.385 145.610 ;
        RECT 131.160 145.410 131.480 145.470 ;
        RECT 132.095 145.425 132.385 145.470 ;
        RECT 133.475 145.425 133.765 145.655 ;
        RECT 133.920 145.610 134.240 145.670 ;
        RECT 134.395 145.610 134.685 145.655 ;
        RECT 133.920 145.470 134.685 145.610 ;
        RECT 133.920 145.410 134.240 145.470 ;
        RECT 134.395 145.425 134.685 145.470 ;
        RECT 134.860 145.610 135.150 145.655 ;
        RECT 136.695 145.610 136.985 145.655 ;
        RECT 140.275 145.610 140.565 145.655 ;
        RECT 134.860 145.470 140.565 145.610 ;
        RECT 134.860 145.425 135.150 145.470 ;
        RECT 136.695 145.425 136.985 145.470 ;
        RECT 140.275 145.425 140.565 145.470 ;
        RECT 141.280 145.450 141.645 145.670 ;
        RECT 142.750 145.610 142.890 145.750 ;
        RECT 144.515 145.610 144.805 145.655 ;
        RECT 142.750 145.470 144.805 145.610 ;
        RECT 145.050 145.610 145.190 146.090 ;
        RECT 145.895 145.610 146.185 145.655 ;
        RECT 145.050 145.470 146.185 145.610 ;
        RECT 141.280 145.410 141.600 145.450 ;
        RECT 144.515 145.425 144.805 145.470 ;
        RECT 145.895 145.425 146.185 145.470 ;
        RECT 122.895 145.270 123.185 145.315 ;
        RECT 125.640 145.270 125.960 145.330 ;
        RECT 122.895 145.130 125.960 145.270 ;
        RECT 122.895 145.085 123.185 145.130 ;
        RECT 125.640 145.070 125.960 145.130 ;
        RECT 127.480 145.270 127.800 145.330 ;
        RECT 127.955 145.270 128.245 145.315 ;
        RECT 127.480 145.130 128.245 145.270 ;
        RECT 127.480 145.070 127.800 145.130 ;
        RECT 127.955 145.085 128.245 145.130 ;
        RECT 128.875 145.270 129.165 145.315 ;
        RECT 129.320 145.270 129.640 145.330 ;
        RECT 128.875 145.130 129.640 145.270 ;
        RECT 128.875 145.085 129.165 145.130 ;
        RECT 129.320 145.070 129.640 145.130 ;
        RECT 131.620 145.070 131.940 145.330 ;
        RECT 135.775 145.270 136.065 145.315 ;
        RECT 135.775 145.130 141.050 145.270 ;
        RECT 135.775 145.085 136.065 145.130 ;
        RECT 123.800 144.930 124.120 144.990 ;
        RECT 120.670 144.790 124.120 144.930 ;
        RECT 131.710 144.930 131.850 145.070 ;
        RECT 135.265 144.930 135.555 144.975 ;
        RECT 137.155 144.930 137.445 144.975 ;
        RECT 140.275 144.930 140.565 144.975 ;
        RECT 131.710 144.790 132.745 144.930 ;
        RECT 75.960 144.590 76.280 144.650 ;
        RECT 71.910 144.450 76.280 144.590 ;
        RECT 75.960 144.390 76.280 144.450 ;
        RECT 79.180 144.390 79.500 144.650 ;
        RECT 84.240 144.390 84.560 144.650 ;
        RECT 88.840 144.390 89.160 144.650 ;
        RECT 92.980 144.390 93.300 144.650 ;
        RECT 96.660 144.590 96.980 144.650 ;
        RECT 98.960 144.590 99.280 144.650 ;
        RECT 96.660 144.450 99.280 144.590 ;
        RECT 96.660 144.390 96.980 144.450 ;
        RECT 98.960 144.390 99.280 144.450 ;
        RECT 100.800 144.590 101.120 144.650 ;
        RECT 107.330 144.590 107.470 144.745 ;
        RECT 110.920 144.730 111.240 144.790 ;
        RECT 115.535 144.745 115.825 144.790 ;
        RECT 117.360 144.730 117.680 144.790 ;
        RECT 123.800 144.730 124.120 144.790 ;
        RECT 100.800 144.450 107.470 144.590 ;
        RECT 123.340 144.590 123.660 144.650 ;
        RECT 130.700 144.590 131.020 144.650 ;
        RECT 123.340 144.450 131.020 144.590 ;
        RECT 100.800 144.390 101.120 144.450 ;
        RECT 123.340 144.390 123.660 144.450 ;
        RECT 130.700 144.390 131.020 144.450 ;
        RECT 131.160 144.390 131.480 144.650 ;
        RECT 131.620 144.590 131.940 144.650 ;
        RECT 132.095 144.590 132.385 144.635 ;
        RECT 131.620 144.450 132.385 144.590 ;
        RECT 132.605 144.590 132.745 144.790 ;
        RECT 135.265 144.790 140.565 144.930 ;
        RECT 140.910 144.930 141.050 145.130 ;
        RECT 144.975 144.930 145.265 144.975 ;
        RECT 140.910 144.790 145.265 144.930 ;
        RECT 135.265 144.745 135.555 144.790 ;
        RECT 137.155 144.745 137.445 144.790 ;
        RECT 140.275 144.745 140.565 144.790 ;
        RECT 144.975 144.745 145.265 144.790 ;
        RECT 135.760 144.590 136.080 144.650 ;
        RECT 132.605 144.450 136.080 144.590 ;
        RECT 131.620 144.390 131.940 144.450 ;
        RECT 132.095 144.405 132.385 144.450 ;
        RECT 135.760 144.390 136.080 144.450 ;
        RECT 143.120 144.390 143.440 144.650 ;
        RECT 2.750 143.770 158.230 144.250 ;
        RECT 6.960 143.570 7.280 143.630 ;
        RECT 13.185 143.570 13.475 143.615 ;
        RECT 14.780 143.570 15.100 143.630 ;
        RECT 21.220 143.570 21.540 143.630 ;
        RECT 6.960 143.430 10.410 143.570 ;
        RECT 6.960 143.370 7.280 143.430 ;
        RECT 4.680 143.230 4.970 143.275 ;
        RECT 6.540 143.230 6.830 143.275 ;
        RECT 9.320 143.230 9.610 143.275 ;
        RECT 4.680 143.090 9.610 143.230 ;
        RECT 10.270 143.230 10.410 143.430 ;
        RECT 13.185 143.430 15.100 143.570 ;
        RECT 13.185 143.385 13.475 143.430 ;
        RECT 14.780 143.370 15.100 143.430 ;
        RECT 15.790 143.430 21.540 143.570 ;
        RECT 15.790 143.230 15.930 143.430 ;
        RECT 21.220 143.370 21.540 143.430 ;
        RECT 23.535 143.570 23.825 143.615 ;
        RECT 26.740 143.570 27.060 143.630 ;
        RECT 23.535 143.430 27.060 143.570 ;
        RECT 23.535 143.385 23.825 143.430 ;
        RECT 26.740 143.370 27.060 143.430 ;
        RECT 27.660 143.570 27.980 143.630 ;
        RECT 36.400 143.570 36.720 143.630 ;
        RECT 38.255 143.570 38.545 143.615 ;
        RECT 27.660 143.430 36.170 143.570 ;
        RECT 27.660 143.370 27.980 143.430 ;
        RECT 10.270 143.090 15.930 143.230 ;
        RECT 4.680 143.045 4.970 143.090 ;
        RECT 6.540 143.045 6.830 143.090 ;
        RECT 9.320 143.045 9.610 143.090 ;
        RECT 16.175 143.045 16.465 143.275 ;
        RECT 4.200 142.890 4.520 142.950 ;
        RECT 16.250 142.890 16.390 143.045 ;
        RECT 20.300 143.030 20.620 143.290 ;
        RECT 30.385 143.230 30.675 143.275 ;
        RECT 32.275 143.230 32.565 143.275 ;
        RECT 35.395 143.230 35.685 143.275 ;
        RECT 30.385 143.090 35.685 143.230 ;
        RECT 36.030 143.230 36.170 143.430 ;
        RECT 36.400 143.430 38.545 143.570 ;
        RECT 36.400 143.370 36.720 143.430 ;
        RECT 38.255 143.385 38.545 143.430 ;
        RECT 41.015 143.570 41.305 143.615 ;
        RECT 42.380 143.570 42.700 143.630 ;
        RECT 41.015 143.430 42.700 143.570 ;
        RECT 41.015 143.385 41.305 143.430 ;
        RECT 42.380 143.370 42.700 143.430 ;
        RECT 42.840 143.570 43.160 143.630 ;
        RECT 47.440 143.570 47.760 143.630 ;
        RECT 42.840 143.430 47.760 143.570 ;
        RECT 42.840 143.370 43.160 143.430 ;
        RECT 47.440 143.370 47.760 143.430 ;
        RECT 49.280 143.570 49.600 143.630 ;
        RECT 52.975 143.570 53.265 143.615 ;
        RECT 57.560 143.570 57.880 143.630 ;
        RECT 49.280 143.430 53.265 143.570 ;
        RECT 49.280 143.370 49.600 143.430 ;
        RECT 52.975 143.385 53.265 143.430 ;
        RECT 54.430 143.430 57.880 143.570 ;
        RECT 41.935 143.230 42.225 143.275 ;
        RECT 36.030 143.090 42.225 143.230 ;
        RECT 30.385 143.045 30.675 143.090 ;
        RECT 32.275 143.045 32.565 143.090 ;
        RECT 35.395 143.045 35.685 143.090 ;
        RECT 41.935 143.045 42.225 143.090 ;
        RECT 44.220 143.230 44.540 143.290 ;
        RECT 44.220 143.090 50.890 143.230 ;
        RECT 44.220 143.030 44.540 143.090 ;
        RECT 4.200 142.750 10.410 142.890 ;
        RECT 4.200 142.690 4.520 142.750 ;
        RECT 10.270 142.610 10.410 142.750 ;
        RECT 15.790 142.750 16.390 142.890 ;
        RECT 6.040 142.350 6.360 142.610 ;
        RECT 9.320 142.550 9.610 142.595 ;
        RECT 7.075 142.410 9.610 142.550 ;
        RECT 7.075 142.255 7.290 142.410 ;
        RECT 9.320 142.365 9.610 142.410 ;
        RECT 10.180 142.350 10.500 142.610 ;
        RECT 14.795 142.550 15.085 142.595 ;
        RECT 15.790 142.550 15.930 142.750 ;
        RECT 18.460 142.690 18.780 142.950 ;
        RECT 19.380 142.690 19.700 142.950 ;
        RECT 14.795 142.410 15.930 142.550 ;
        RECT 20.390 142.550 20.530 143.030 ;
        RECT 29.515 142.890 29.805 142.935 ;
        RECT 34.560 142.890 34.880 142.950 ;
        RECT 37.780 142.890 38.100 142.950 ;
        RECT 42.840 142.890 43.160 142.950 ;
        RECT 45.140 142.890 45.460 142.950 ;
        RECT 21.310 142.750 23.290 142.890 ;
        RECT 21.310 142.595 21.450 142.750 ;
        RECT 23.150 142.610 23.290 142.750 ;
        RECT 29.515 142.750 37.550 142.890 ;
        RECT 29.515 142.705 29.805 142.750 ;
        RECT 34.560 142.690 34.880 142.750 ;
        RECT 20.775 142.550 21.065 142.595 ;
        RECT 20.390 142.410 21.065 142.550 ;
        RECT 14.795 142.365 15.085 142.410 ;
        RECT 20.775 142.365 21.065 142.410 ;
        RECT 21.235 142.365 21.525 142.595 ;
        RECT 22.155 142.365 22.445 142.595 ;
        RECT 22.615 142.365 22.905 142.595 ;
        RECT 11.100 142.255 11.420 142.270 ;
        RECT 5.140 142.210 5.430 142.255 ;
        RECT 7.000 142.210 7.290 142.255 ;
        RECT 5.140 142.070 7.290 142.210 ;
        RECT 5.140 142.025 5.430 142.070 ;
        RECT 7.000 142.025 7.290 142.070 ;
        RECT 7.920 142.210 8.210 142.255 ;
        RECT 11.100 142.210 11.470 142.255 ;
        RECT 7.920 142.070 11.470 142.210 ;
        RECT 7.920 142.025 8.210 142.070 ;
        RECT 11.100 142.025 11.470 142.070 ;
        RECT 18.015 142.210 18.305 142.255 ;
        RECT 19.840 142.210 20.160 142.270 ;
        RECT 22.230 142.210 22.370 142.365 ;
        RECT 18.015 142.070 20.160 142.210 ;
        RECT 18.015 142.025 18.305 142.070 ;
        RECT 11.100 142.010 11.420 142.025 ;
        RECT 13.860 141.670 14.180 141.930 ;
        RECT 14.320 141.870 14.640 141.930 ;
        RECT 18.090 141.870 18.230 142.025 ;
        RECT 19.840 142.010 20.160 142.070 ;
        RECT 20.850 142.070 22.370 142.210 ;
        RECT 22.690 142.210 22.830 142.365 ;
        RECT 23.060 142.350 23.380 142.610 ;
        RECT 23.980 142.350 24.300 142.610 ;
        RECT 25.820 142.550 26.140 142.610 ;
        RECT 24.530 142.410 26.140 142.550 ;
        RECT 24.530 142.210 24.670 142.410 ;
        RECT 25.820 142.350 26.140 142.410 ;
        RECT 28.120 142.550 28.440 142.610 ;
        RECT 28.595 142.550 28.885 142.595 ;
        RECT 28.120 142.410 28.885 142.550 ;
        RECT 28.120 142.350 28.440 142.410 ;
        RECT 28.595 142.365 28.885 142.410 ;
        RECT 29.980 142.550 30.270 142.595 ;
        RECT 31.815 142.550 32.105 142.595 ;
        RECT 35.395 142.550 35.685 142.595 ;
        RECT 29.980 142.410 35.685 142.550 ;
        RECT 29.980 142.365 30.270 142.410 ;
        RECT 31.815 142.365 32.105 142.410 ;
        RECT 35.395 142.365 35.685 142.410 ;
        RECT 35.940 142.550 36.260 142.610 ;
        RECT 36.475 142.550 36.765 142.570 ;
        RECT 35.940 142.410 36.765 142.550 ;
        RECT 35.940 142.350 36.260 142.410 ;
        RECT 36.475 142.255 36.765 142.410 ;
        RECT 30.895 142.210 31.185 142.255 ;
        RECT 22.690 142.070 24.670 142.210 ;
        RECT 24.990 142.070 31.185 142.210 ;
        RECT 20.850 141.930 20.990 142.070 ;
        RECT 14.320 141.730 18.230 141.870 ;
        RECT 14.320 141.670 14.640 141.730 ;
        RECT 20.760 141.670 21.080 141.930 ;
        RECT 24.990 141.915 25.130 142.070 ;
        RECT 30.895 142.025 31.185 142.070 ;
        RECT 33.175 142.210 33.825 142.255 ;
        RECT 36.475 142.210 37.065 142.255 ;
        RECT 33.175 142.070 37.065 142.210 ;
        RECT 33.175 142.025 33.825 142.070 ;
        RECT 36.775 142.025 37.065 142.070 ;
        RECT 24.915 141.685 25.205 141.915 ;
        RECT 25.820 141.670 26.140 141.930 ;
        RECT 37.410 141.870 37.550 142.750 ;
        RECT 37.780 142.750 40.770 142.890 ;
        RECT 37.780 142.690 38.100 142.750 ;
        RECT 38.700 142.350 39.020 142.610 ;
        RECT 39.160 142.350 39.480 142.610 ;
        RECT 40.080 142.350 40.400 142.610 ;
        RECT 40.630 142.210 40.770 142.750 ;
        RECT 42.840 142.750 45.460 142.890 ;
        RECT 42.840 142.690 43.160 142.750 ;
        RECT 45.140 142.690 45.460 142.750 ;
        RECT 48.360 142.890 48.680 142.950 ;
        RECT 48.835 142.890 49.125 142.935 ;
        RECT 48.360 142.750 49.125 142.890 ;
        RECT 48.360 142.690 48.680 142.750 ;
        RECT 48.835 142.705 49.125 142.750 ;
        RECT 46.060 142.550 46.380 142.610 ;
        RECT 49.755 142.550 50.045 142.595 ;
        RECT 46.060 142.410 50.045 142.550 ;
        RECT 46.060 142.350 46.380 142.410 ;
        RECT 49.755 142.365 50.045 142.410 ;
        RECT 50.220 142.365 50.510 142.595 ;
        RECT 50.750 142.550 50.890 143.090 ;
        RECT 51.120 142.890 51.440 142.950 ;
        RECT 54.430 142.935 54.570 143.430 ;
        RECT 57.560 143.370 57.880 143.430 ;
        RECT 59.860 143.570 60.180 143.630 ;
        RECT 64.920 143.570 65.240 143.630 ;
        RECT 59.860 143.430 65.240 143.570 ;
        RECT 59.860 143.370 60.180 143.430 ;
        RECT 64.920 143.370 65.240 143.430 ;
        RECT 69.995 143.570 70.285 143.615 ;
        RECT 70.440 143.570 70.760 143.630 ;
        RECT 69.995 143.430 70.760 143.570 ;
        RECT 69.995 143.385 70.285 143.430 ;
        RECT 70.440 143.370 70.760 143.430 ;
        RECT 71.820 143.570 72.140 143.630 ;
        RECT 73.660 143.570 73.980 143.630 ;
        RECT 71.820 143.430 73.980 143.570 ;
        RECT 71.820 143.370 72.140 143.430 ;
        RECT 73.660 143.370 73.980 143.430 ;
        RECT 78.720 143.370 79.040 143.630 ;
        RECT 82.875 143.385 83.165 143.615 ;
        RECT 83.795 143.570 84.085 143.615 ;
        RECT 88.380 143.570 88.700 143.630 ;
        RECT 83.795 143.430 88.700 143.570 ;
        RECT 83.795 143.385 84.085 143.430 ;
        RECT 57.115 143.230 57.405 143.275 ;
        RECT 59.400 143.230 59.720 143.290 ;
        RECT 57.115 143.090 59.720 143.230 ;
        RECT 57.115 143.045 57.405 143.090 ;
        RECT 59.400 143.030 59.720 143.090 ;
        RECT 61.670 143.230 61.960 143.275 ;
        RECT 64.450 143.230 64.740 143.275 ;
        RECT 66.310 143.230 66.600 143.275 ;
        RECT 61.670 143.090 66.600 143.230 ;
        RECT 61.670 143.045 61.960 143.090 ;
        RECT 64.450 143.045 64.740 143.090 ;
        RECT 66.310 143.045 66.600 143.090 ;
        RECT 69.535 143.230 69.825 143.275 ;
        RECT 78.810 143.230 78.950 143.370 ;
        RECT 69.535 143.090 78.950 143.230 ;
        RECT 69.535 143.045 69.825 143.090 ;
        RECT 79.195 143.045 79.485 143.275 ;
        RECT 82.950 143.230 83.090 143.385 ;
        RECT 88.380 143.370 88.700 143.430 ;
        RECT 88.840 143.370 89.160 143.630 ;
        RECT 89.300 143.370 89.620 143.630 ;
        RECT 90.220 143.370 90.540 143.630 ;
        RECT 92.980 143.570 93.300 143.630 ;
        RECT 105.860 143.570 106.180 143.630 ;
        RECT 116.915 143.570 117.205 143.615 ;
        RECT 129.320 143.570 129.640 143.630 ;
        RECT 92.980 143.430 105.630 143.570 ;
        RECT 92.980 143.370 93.300 143.430 ;
        RECT 82.950 143.090 85.390 143.230 ;
        RECT 54.355 142.890 54.645 142.935 ;
        RECT 51.120 142.750 54.645 142.890 ;
        RECT 51.120 142.690 51.440 142.750 ;
        RECT 54.355 142.705 54.645 142.750 ;
        RECT 54.815 142.890 55.105 142.935 ;
        RECT 56.180 142.890 56.500 142.950 ;
        RECT 57.805 142.890 58.095 142.935 ;
        RECT 54.815 142.750 58.095 142.890 ;
        RECT 54.815 142.705 55.105 142.750 ;
        RECT 56.180 142.690 56.500 142.750 ;
        RECT 57.805 142.705 58.095 142.750 ;
        RECT 66.760 142.690 67.080 142.950 ;
        RECT 68.525 142.890 68.815 142.935 ;
        RECT 70.900 142.890 71.220 142.950 ;
        RECT 68.525 142.750 71.220 142.890 ;
        RECT 68.525 142.705 68.815 142.750 ;
        RECT 70.900 142.690 71.220 142.750 ;
        RECT 72.740 142.890 73.060 142.950 ;
        RECT 73.215 142.890 73.505 142.935 ;
        RECT 75.040 142.890 75.360 142.950 ;
        RECT 76.435 142.890 76.725 142.935 ;
        RECT 72.740 142.750 76.725 142.890 ;
        RECT 79.270 142.890 79.410 143.045 ;
        RECT 83.320 142.890 83.640 142.950 ;
        RECT 79.270 142.750 83.640 142.890 ;
        RECT 72.740 142.690 73.060 142.750 ;
        RECT 73.215 142.705 73.505 142.750 ;
        RECT 75.040 142.690 75.360 142.750 ;
        RECT 76.435 142.705 76.725 142.750 ;
        RECT 83.320 142.690 83.640 142.750 ;
        RECT 52.080 142.550 52.370 142.595 ;
        RECT 61.670 142.550 61.960 142.595 ;
        RECT 64.935 142.550 65.225 142.595 ;
        RECT 65.380 142.550 65.700 142.610 ;
        RECT 50.750 142.410 52.370 142.550 ;
        RECT 52.080 142.365 52.370 142.410 ;
        RECT 53.050 142.410 56.870 142.550 ;
        RECT 50.290 142.210 50.430 142.365 ;
        RECT 40.630 142.070 50.430 142.210 ;
        RECT 51.135 142.025 51.425 142.255 ;
        RECT 51.595 142.210 51.885 142.255 ;
        RECT 53.050 142.210 53.190 142.410 ;
        RECT 56.730 142.270 56.870 142.410 ;
        RECT 61.670 142.410 64.205 142.550 ;
        RECT 61.670 142.365 61.960 142.410 ;
        RECT 51.595 142.070 53.190 142.210 ;
        RECT 53.420 142.210 53.740 142.270 ;
        RECT 55.275 142.210 55.565 142.255 ;
        RECT 53.420 142.070 55.565 142.210 ;
        RECT 51.595 142.025 51.885 142.070 ;
        RECT 40.080 141.870 40.400 141.930 ;
        RECT 37.410 141.730 40.400 141.870 ;
        RECT 40.080 141.670 40.400 141.730 ;
        RECT 43.760 141.670 44.080 141.930 ;
        RECT 44.235 141.870 44.525 141.915 ;
        RECT 46.075 141.870 46.365 141.915 ;
        RECT 44.235 141.730 46.365 141.870 ;
        RECT 44.235 141.685 44.525 141.730 ;
        RECT 46.075 141.685 46.365 141.730 ;
        RECT 47.440 141.870 47.760 141.930 ;
        RECT 51.210 141.870 51.350 142.025 ;
        RECT 53.420 142.010 53.740 142.070 ;
        RECT 55.275 142.025 55.565 142.070 ;
        RECT 47.440 141.730 51.350 141.870 ;
        RECT 55.350 141.870 55.490 142.025 ;
        RECT 56.640 142.010 56.960 142.270 ;
        RECT 63.080 142.255 63.400 142.270 ;
        RECT 59.810 142.210 60.100 142.255 ;
        RECT 63.070 142.210 63.400 142.255 ;
        RECT 59.810 142.070 63.400 142.210 ;
        RECT 59.810 142.025 60.100 142.070 ;
        RECT 63.070 142.025 63.400 142.070 ;
        RECT 63.990 142.255 64.205 142.410 ;
        RECT 64.935 142.410 65.700 142.550 ;
        RECT 64.935 142.365 65.225 142.410 ;
        RECT 65.380 142.350 65.700 142.410 ;
        RECT 67.680 142.350 68.000 142.610 ;
        RECT 69.075 142.550 69.365 142.595 ;
        RECT 68.230 142.410 69.365 142.550 ;
        RECT 63.990 142.210 64.280 142.255 ;
        RECT 65.850 142.210 66.140 142.255 ;
        RECT 63.990 142.070 66.140 142.210 ;
        RECT 63.990 142.025 64.280 142.070 ;
        RECT 65.850 142.025 66.140 142.070 ;
        RECT 63.080 142.010 63.400 142.025 ;
        RECT 68.230 141.930 68.370 142.410 ;
        RECT 69.075 142.365 69.365 142.410 ;
        RECT 69.980 142.550 70.300 142.610 ;
        RECT 70.455 142.550 70.745 142.595 ;
        RECT 69.980 142.410 70.745 142.550 ;
        RECT 69.980 142.350 70.300 142.410 ;
        RECT 70.455 142.365 70.745 142.410 ;
        RECT 71.360 142.550 71.680 142.610 ;
        RECT 71.835 142.550 72.125 142.595 ;
        RECT 75.500 142.550 75.820 142.610 ;
        RECT 71.360 142.535 72.125 142.550 ;
        RECT 72.825 142.535 75.820 142.550 ;
        RECT 71.360 142.410 75.820 142.535 ;
        RECT 71.360 142.350 71.680 142.410 ;
        RECT 71.835 142.395 72.965 142.410 ;
        RECT 71.835 142.365 72.125 142.395 ;
        RECT 75.500 142.350 75.820 142.410 ;
        RECT 81.495 142.365 81.785 142.595 ;
        RECT 76.880 142.010 77.200 142.270 ;
        RECT 77.800 142.010 78.120 142.270 ;
        RECT 81.570 141.930 81.710 142.365 ;
        RECT 85.250 142.270 85.390 143.090 ;
        RECT 88.930 142.890 89.070 143.370 ;
        RECT 90.310 142.890 90.450 143.370 ;
        RECT 90.680 143.230 91.000 143.290 ;
        RECT 98.500 143.230 98.820 143.290 ;
        RECT 105.490 143.230 105.630 143.430 ;
        RECT 105.860 143.430 115.290 143.570 ;
        RECT 105.860 143.370 106.180 143.430 ;
        RECT 106.320 143.230 106.640 143.290 ;
        RECT 90.680 143.090 100.110 143.230 ;
        RECT 105.490 143.090 106.640 143.230 ;
        RECT 90.680 143.030 91.000 143.090 ;
        RECT 98.500 143.030 98.820 143.090 ;
        RECT 99.970 142.890 100.110 143.090 ;
        RECT 106.320 143.030 106.640 143.090 ;
        RECT 106.780 143.230 107.100 143.290 ;
        RECT 115.150 143.230 115.290 143.430 ;
        RECT 116.915 143.430 129.640 143.570 ;
        RECT 116.915 143.385 117.205 143.430 ;
        RECT 129.320 143.370 129.640 143.430 ;
        RECT 131.160 143.570 131.480 143.630 ;
        RECT 140.820 143.570 141.140 143.630 ;
        RECT 131.160 143.430 141.140 143.570 ;
        RECT 131.160 143.370 131.480 143.430 ;
        RECT 140.820 143.370 141.140 143.430 ;
        RECT 141.740 143.370 142.060 143.630 ;
        RECT 143.120 143.370 143.440 143.630 ;
        RECT 125.640 143.230 125.960 143.290 ;
        RECT 129.780 143.230 130.100 143.290 ;
        RECT 141.830 143.230 141.970 143.370 ;
        RECT 106.780 143.090 114.830 143.230 ;
        RECT 115.150 143.090 120.325 143.230 ;
        RECT 106.780 143.030 107.100 143.090 ;
        RECT 100.355 142.890 100.645 142.935 ;
        RECT 101.260 142.890 101.580 142.950 ;
        RECT 88.010 142.750 89.070 142.890 ;
        RECT 89.850 142.750 99.650 142.890 ;
        RECT 99.970 142.750 101.950 142.890 ;
        RECT 88.010 142.595 88.150 142.750 ;
        RECT 87.935 142.365 88.225 142.595 ;
        RECT 88.855 142.550 89.145 142.595 ;
        RECT 89.850 142.550 89.990 142.750 ;
        RECT 88.855 142.410 89.990 142.550 ;
        RECT 88.855 142.365 89.145 142.410 ;
        RECT 90.235 142.365 90.525 142.595 ;
        RECT 90.695 142.550 90.985 142.595 ;
        RECT 90.695 142.410 91.830 142.550 ;
        RECT 90.695 142.365 90.985 142.410 ;
        RECT 85.160 142.210 85.480 142.270 ;
        RECT 87.015 142.210 87.305 142.255 ;
        RECT 85.160 142.070 87.305 142.210 ;
        RECT 85.160 142.010 85.480 142.070 ;
        RECT 87.015 142.025 87.305 142.070 ;
        RECT 68.140 141.870 68.460 141.930 ;
        RECT 55.350 141.730 68.460 141.870 ;
        RECT 47.440 141.670 47.760 141.730 ;
        RECT 68.140 141.670 68.460 141.730 ;
        RECT 74.580 141.670 74.900 141.930 ;
        RECT 81.480 141.670 81.800 141.930 ;
        RECT 82.400 141.870 82.720 141.930 ;
        RECT 90.310 141.870 90.450 142.365 ;
        RECT 91.690 142.270 91.830 142.410 ;
        RECT 92.060 142.350 92.380 142.610 ;
        RECT 92.520 142.550 92.840 142.610 ;
        RECT 92.520 142.410 98.730 142.550 ;
        RECT 92.520 142.350 92.840 142.410 ;
        RECT 91.140 142.010 91.460 142.270 ;
        RECT 91.600 142.210 91.920 142.270 ;
        RECT 96.200 142.210 96.520 142.270 ;
        RECT 91.600 142.070 96.520 142.210 ;
        RECT 91.600 142.010 91.920 142.070 ;
        RECT 96.200 142.010 96.520 142.070 ;
        RECT 82.400 141.730 90.450 141.870 ;
        RECT 82.400 141.670 82.720 141.730 ;
        RECT 98.040 141.670 98.360 141.930 ;
        RECT 98.590 141.870 98.730 142.410 ;
        RECT 98.960 142.350 99.280 142.610 ;
        RECT 99.510 142.210 99.650 142.750 ;
        RECT 100.355 142.705 100.645 142.750 ;
        RECT 101.260 142.690 101.580 142.750 ;
        RECT 99.880 142.550 100.200 142.610 ;
        RECT 101.810 142.595 101.950 142.750 ;
        RECT 108.620 142.690 108.940 142.950 ;
        RECT 112.300 142.890 112.620 142.950 ;
        RECT 114.690 142.935 114.830 143.090 ;
        RECT 114.155 142.890 114.445 142.935 ;
        RECT 112.300 142.750 114.445 142.890 ;
        RECT 112.300 142.690 112.620 142.750 ;
        RECT 114.155 142.705 114.445 142.750 ;
        RECT 114.615 142.705 114.905 142.935 ;
        RECT 100.815 142.550 101.105 142.595 ;
        RECT 99.880 142.410 101.105 142.550 ;
        RECT 99.880 142.350 100.200 142.410 ;
        RECT 100.815 142.365 101.105 142.410 ;
        RECT 101.735 142.365 102.025 142.595 ;
        RECT 104.955 142.550 105.245 142.595 ;
        RECT 105.400 142.550 105.720 142.610 ;
        RECT 104.955 142.410 105.720 142.550 ;
        RECT 104.955 142.365 105.245 142.410 ;
        RECT 105.400 142.350 105.720 142.410 ;
        RECT 105.875 142.365 106.165 142.595 ;
        RECT 106.335 142.550 106.625 142.595 ;
        RECT 106.795 142.550 107.085 142.595 ;
        RECT 108.710 142.550 108.850 142.690 ;
        RECT 120.185 142.610 120.325 143.090 ;
        RECT 125.640 143.090 130.100 143.230 ;
        RECT 125.640 143.030 125.960 143.090 ;
        RECT 129.780 143.030 130.100 143.090 ;
        RECT 137.230 143.090 141.970 143.230 ;
        RECT 122.895 142.890 123.185 142.935 ;
        RECT 122.510 142.750 123.185 142.890 ;
        RECT 106.335 142.410 108.850 142.550 ;
        RECT 106.335 142.365 106.625 142.410 ;
        RECT 106.795 142.365 107.085 142.410 ;
        RECT 100.340 142.210 100.660 142.270 ;
        RECT 101.275 142.210 101.565 142.255 ;
        RECT 102.640 142.210 102.960 142.270 ;
        RECT 105.950 142.210 106.090 142.365 ;
        RECT 109.080 142.350 109.400 142.610 ;
        RECT 110.000 142.350 110.320 142.610 ;
        RECT 110.460 142.550 110.780 142.610 ;
        RECT 120.120 142.595 120.440 142.610 ;
        RECT 120.110 142.550 120.440 142.595 ;
        RECT 121.960 142.550 122.280 142.610 ;
        RECT 122.510 142.595 122.650 142.750 ;
        RECT 122.895 142.705 123.185 142.750 ;
        RECT 123.800 142.890 124.120 142.950 ;
        RECT 123.800 142.750 132.310 142.890 ;
        RECT 123.800 142.690 124.120 142.750 ;
        RECT 110.460 142.410 119.430 142.550 ;
        RECT 119.925 142.410 120.440 142.550 ;
        RECT 121.765 142.410 122.280 142.550 ;
        RECT 110.460 142.350 110.780 142.410 ;
        RECT 108.160 142.210 108.480 142.270 ;
        RECT 110.090 142.210 110.230 142.350 ;
        RECT 99.510 142.070 102.960 142.210 ;
        RECT 100.340 142.010 100.660 142.070 ;
        RECT 101.275 142.025 101.565 142.070 ;
        RECT 102.640 142.010 102.960 142.070 ;
        RECT 103.650 142.070 110.230 142.210 ;
        RECT 114.140 142.210 114.460 142.270 ;
        RECT 114.615 142.210 114.905 142.255 ;
        RECT 114.140 142.070 114.905 142.210 ;
        RECT 103.650 141.870 103.790 142.070 ;
        RECT 108.160 142.010 108.480 142.070 ;
        RECT 114.140 142.010 114.460 142.070 ;
        RECT 114.615 142.025 114.905 142.070 ;
        RECT 98.590 141.730 103.790 141.870 ;
        RECT 104.035 141.870 104.325 141.915 ;
        RECT 110.920 141.870 111.240 141.930 ;
        RECT 104.035 141.730 111.240 141.870 ;
        RECT 104.035 141.685 104.325 141.730 ;
        RECT 110.920 141.670 111.240 141.730 ;
        RECT 112.300 141.870 112.620 141.930 ;
        RECT 119.290 141.915 119.430 142.410 ;
        RECT 120.110 142.365 120.440 142.410 ;
        RECT 120.120 142.350 120.440 142.365 ;
        RECT 121.960 142.350 122.280 142.410 ;
        RECT 122.435 142.365 122.725 142.595 ;
        RECT 123.340 142.550 123.660 142.610 ;
        RECT 124.275 142.550 124.565 142.595 ;
        RECT 123.340 142.410 124.565 142.550 ;
        RECT 123.340 142.350 123.660 142.410 ;
        RECT 124.275 142.365 124.565 142.410 ;
        RECT 124.720 142.350 125.040 142.610 ;
        RECT 125.195 142.365 125.485 142.595 ;
        RECT 125.640 142.550 125.960 142.610 ;
        RECT 126.115 142.550 126.405 142.595 ;
        RECT 125.640 142.410 126.405 142.550 ;
        RECT 120.580 142.010 120.900 142.270 ;
        RECT 121.055 142.025 121.345 142.255 ;
        RECT 125.270 142.210 125.410 142.365 ;
        RECT 125.640 142.350 125.960 142.410 ;
        RECT 126.115 142.365 126.405 142.410 ;
        RECT 126.560 142.550 126.880 142.610 ;
        RECT 127.495 142.550 127.785 142.595 ;
        RECT 126.560 142.410 127.785 142.550 ;
        RECT 126.560 142.350 126.880 142.410 ;
        RECT 127.495 142.365 127.785 142.410 ;
        RECT 127.940 142.350 128.260 142.610 ;
        RECT 128.400 142.350 128.720 142.610 ;
        RECT 128.860 142.350 129.180 142.610 ;
        RECT 132.170 142.595 132.310 142.750 ;
        RECT 130.715 142.365 131.005 142.595 ;
        RECT 132.095 142.365 132.385 142.595 ;
        RECT 129.795 142.210 130.085 142.255 ;
        RECT 125.270 142.070 130.085 142.210 ;
        RECT 129.795 142.025 130.085 142.070 ;
        RECT 113.235 141.870 113.525 141.915 ;
        RECT 112.300 141.730 113.525 141.870 ;
        RECT 112.300 141.670 112.620 141.730 ;
        RECT 113.235 141.685 113.525 141.730 ;
        RECT 119.215 141.685 119.505 141.915 ;
        RECT 121.130 141.870 121.270 142.025 ;
        RECT 125.640 141.870 125.960 141.930 ;
        RECT 121.130 141.730 125.960 141.870 ;
        RECT 125.640 141.670 125.960 141.730 ;
        RECT 126.560 141.670 126.880 141.930 ;
        RECT 127.940 141.870 128.260 141.930 ;
        RECT 130.790 141.870 130.930 142.365 ;
        RECT 133.460 142.350 133.780 142.610 ;
        RECT 135.760 142.350 136.080 142.610 ;
        RECT 136.680 142.550 137.000 142.610 ;
        RECT 137.230 142.595 137.370 143.090 ;
        RECT 143.210 142.890 143.350 143.370 ;
        RECT 137.690 142.750 141.970 142.890 ;
        RECT 143.210 142.750 144.270 142.890 ;
        RECT 137.155 142.550 137.445 142.595 ;
        RECT 136.680 142.410 137.445 142.550 ;
        RECT 136.680 142.350 137.000 142.410 ;
        RECT 137.155 142.365 137.445 142.410 ;
        RECT 135.850 142.210 135.990 142.350 ;
        RECT 137.690 142.210 137.830 142.750 ;
        RECT 140.360 142.350 140.680 142.610 ;
        RECT 141.830 142.270 141.970 142.750 ;
        RECT 143.135 142.550 143.425 142.595 ;
        RECT 143.580 142.550 143.900 142.610 ;
        RECT 144.130 142.595 144.270 142.750 ;
        RECT 143.135 142.410 143.900 142.550 ;
        RECT 143.135 142.365 143.425 142.410 ;
        RECT 135.850 142.070 137.830 142.210 ;
        RECT 138.060 142.210 138.380 142.270 ;
        RECT 139.900 142.210 140.220 142.270 ;
        RECT 138.060 142.070 140.220 142.210 ;
        RECT 138.060 142.010 138.380 142.070 ;
        RECT 139.900 142.010 140.220 142.070 ;
        RECT 141.740 142.010 142.060 142.270 ;
        RECT 143.210 142.210 143.350 142.365 ;
        RECT 143.580 142.350 143.900 142.410 ;
        RECT 144.055 142.550 144.345 142.595 ;
        RECT 146.800 142.550 147.120 142.610 ;
        RECT 144.055 142.410 147.120 142.550 ;
        RECT 144.055 142.365 144.345 142.410 ;
        RECT 146.800 142.350 147.120 142.410 ;
        RECT 143.210 142.070 148.410 142.210 ;
        RECT 148.270 141.930 148.410 142.070 ;
        RECT 127.940 141.730 130.930 141.870 ;
        RECT 131.160 141.870 131.480 141.930 ;
        RECT 131.635 141.870 131.925 141.915 ;
        RECT 133.000 141.870 133.320 141.930 ;
        RECT 131.160 141.730 133.320 141.870 ;
        RECT 127.940 141.670 128.260 141.730 ;
        RECT 131.160 141.670 131.480 141.730 ;
        RECT 131.635 141.685 131.925 141.730 ;
        RECT 133.000 141.670 133.320 141.730 ;
        RECT 134.840 141.870 135.160 141.930 ;
        RECT 143.595 141.870 143.885 141.915 ;
        RECT 134.840 141.730 143.885 141.870 ;
        RECT 134.840 141.670 135.160 141.730 ;
        RECT 143.595 141.685 143.885 141.730 ;
        RECT 144.960 141.870 145.280 141.930 ;
        RECT 145.435 141.870 145.725 141.915 ;
        RECT 144.960 141.730 145.725 141.870 ;
        RECT 144.960 141.670 145.280 141.730 ;
        RECT 145.435 141.685 145.725 141.730 ;
        RECT 148.180 141.670 148.500 141.930 ;
        RECT 2.750 141.050 159.030 141.530 ;
        RECT 7.420 140.650 7.740 140.910 ;
        RECT 9.720 140.850 10.040 140.910 ;
        RECT 14.320 140.850 14.640 140.910 ;
        RECT 8.890 140.710 10.040 140.850 ;
        RECT 3.740 140.510 4.060 140.570 ;
        RECT 5.595 140.510 5.885 140.555 ;
        RECT 8.890 140.510 9.030 140.710 ;
        RECT 9.720 140.650 10.040 140.710 ;
        RECT 10.730 140.710 14.640 140.850 ;
        RECT 3.740 140.370 5.350 140.510 ;
        RECT 3.740 140.310 4.060 140.370 ;
        RECT 4.675 139.985 4.965 140.215 ;
        RECT 4.750 139.150 4.890 139.985 ;
        RECT 5.210 139.830 5.350 140.370 ;
        RECT 5.595 140.370 9.030 140.510 ;
        RECT 5.595 140.325 5.885 140.370 ;
        RECT 9.260 140.310 9.580 140.570 ;
        RECT 6.055 139.985 6.345 140.215 ;
        RECT 6.515 140.170 6.805 140.215 ;
        RECT 8.800 140.170 9.120 140.230 ;
        RECT 9.810 140.215 9.950 140.650 ;
        RECT 10.730 140.215 10.870 140.710 ;
        RECT 14.320 140.650 14.640 140.710 ;
        RECT 18.920 140.850 19.240 140.910 ;
        RECT 20.085 140.850 20.375 140.895 ;
        RECT 18.920 140.710 20.375 140.850 ;
        RECT 18.920 140.650 19.240 140.710 ;
        RECT 20.085 140.665 20.375 140.710 ;
        RECT 23.980 140.650 24.300 140.910 ;
        RECT 25.820 140.850 26.140 140.910 ;
        RECT 26.755 140.850 27.045 140.895 ;
        RECT 25.820 140.710 27.045 140.850 ;
        RECT 25.820 140.650 26.140 140.710 ;
        RECT 26.755 140.665 27.045 140.710 ;
        RECT 29.960 140.850 30.280 140.910 ;
        RECT 30.895 140.850 31.185 140.895 ;
        RECT 29.960 140.710 31.185 140.850 ;
        RECT 29.960 140.650 30.280 140.710 ;
        RECT 30.895 140.665 31.185 140.710 ;
        RECT 31.340 140.650 31.660 140.910 ;
        RECT 33.195 140.665 33.485 140.895 ;
        RECT 12.040 140.510 12.330 140.555 ;
        RECT 13.900 140.510 14.190 140.555 ;
        RECT 12.040 140.370 14.190 140.510 ;
        RECT 12.040 140.325 12.330 140.370 ;
        RECT 13.900 140.325 14.190 140.370 ;
        RECT 14.820 140.510 15.110 140.555 ;
        RECT 18.080 140.510 18.370 140.555 ;
        RECT 14.820 140.370 18.370 140.510 ;
        RECT 24.070 140.510 24.210 140.650 ;
        RECT 33.270 140.510 33.410 140.665 ;
        RECT 34.560 140.650 34.880 140.910 ;
        RECT 35.495 140.850 35.785 140.895 ;
        RECT 36.860 140.850 37.180 140.910 ;
        RECT 35.495 140.710 37.180 140.850 ;
        RECT 35.495 140.665 35.785 140.710 ;
        RECT 36.860 140.650 37.180 140.710 ;
        RECT 38.240 140.850 38.560 140.910 ;
        RECT 38.715 140.850 39.005 140.895 ;
        RECT 38.240 140.710 39.005 140.850 ;
        RECT 38.240 140.650 38.560 140.710 ;
        RECT 38.715 140.665 39.005 140.710 ;
        RECT 42.840 140.650 43.160 140.910 ;
        RECT 43.760 140.850 44.080 140.910 ;
        RECT 46.060 140.850 46.380 140.910 ;
        RECT 43.760 140.710 46.380 140.850 ;
        RECT 43.760 140.650 44.080 140.710 ;
        RECT 46.060 140.650 46.380 140.710 ;
        RECT 46.535 140.850 46.825 140.895 ;
        RECT 64.015 140.850 64.305 140.895 ;
        RECT 46.535 140.710 64.305 140.850 ;
        RECT 46.535 140.665 46.825 140.710 ;
        RECT 64.015 140.665 64.305 140.710 ;
        RECT 68.140 140.650 68.460 140.910 ;
        RECT 69.995 140.850 70.285 140.895 ;
        RECT 69.995 140.710 74.350 140.850 ;
        RECT 69.995 140.665 70.285 140.710 ;
        RECT 24.070 140.370 33.410 140.510 ;
        RECT 14.820 140.325 15.110 140.370 ;
        RECT 18.080 140.325 18.370 140.370 ;
        RECT 6.515 140.030 9.120 140.170 ;
        RECT 6.515 139.985 6.805 140.030 ;
        RECT 6.130 139.830 6.270 139.985 ;
        RECT 8.800 139.970 9.120 140.030 ;
        RECT 9.735 139.985 10.025 140.215 ;
        RECT 10.655 139.985 10.945 140.215 ;
        RECT 11.115 140.170 11.405 140.215 ;
        RECT 13.400 140.170 13.720 140.230 ;
        RECT 11.115 140.030 13.720 140.170 ;
        RECT 13.975 140.170 14.190 140.325 ;
        RECT 16.220 140.170 16.510 140.215 ;
        RECT 13.975 140.030 16.510 140.170 ;
        RECT 18.090 140.170 18.230 140.325 ;
        RECT 20.300 140.170 20.620 140.230 ;
        RECT 18.090 140.030 20.620 140.170 ;
        RECT 11.115 139.985 11.405 140.030 ;
        RECT 5.210 139.690 6.270 139.830 ;
        RECT 10.180 139.830 10.500 139.890 ;
        RECT 11.190 139.830 11.330 139.985 ;
        RECT 13.400 139.970 13.720 140.030 ;
        RECT 16.220 139.985 16.510 140.030 ;
        RECT 20.300 139.970 20.620 140.030 ;
        RECT 21.220 140.170 21.540 140.230 ;
        RECT 23.060 140.170 23.380 140.230 ;
        RECT 23.535 140.170 23.825 140.215 ;
        RECT 21.220 140.030 23.825 140.170 ;
        RECT 21.220 139.970 21.540 140.030 ;
        RECT 23.060 139.970 23.380 140.030 ;
        RECT 23.535 139.985 23.825 140.030 ;
        RECT 26.280 140.170 26.600 140.230 ;
        RECT 29.960 140.170 30.280 140.230 ;
        RECT 30.880 140.170 31.200 140.230 ;
        RECT 34.650 140.170 34.790 140.650 ;
        RECT 42.930 140.510 43.070 140.650 ;
        RECT 36.515 140.370 43.070 140.510 ;
        RECT 43.315 140.510 43.605 140.555 ;
        RECT 46.980 140.510 47.300 140.570 ;
        RECT 53.420 140.510 53.740 140.570 ;
        RECT 56.195 140.510 56.485 140.555 ;
        RECT 43.315 140.370 47.300 140.510 ;
        RECT 35.020 140.170 35.340 140.230 ;
        RECT 26.280 140.030 30.280 140.170 ;
        RECT 26.280 139.970 26.600 140.030 ;
        RECT 29.960 139.970 30.280 140.030 ;
        RECT 30.510 140.030 32.490 140.170 ;
        RECT 34.650 140.030 35.340 140.170 ;
        RECT 10.180 139.690 11.330 139.830 ;
        RECT 12.955 139.830 13.245 139.875 ;
        RECT 13.860 139.830 14.180 139.890 ;
        RECT 12.955 139.690 14.180 139.830 ;
        RECT 10.180 139.630 10.500 139.690 ;
        RECT 12.955 139.645 13.245 139.690 ;
        RECT 13.860 139.630 14.180 139.690 ;
        RECT 19.380 139.830 19.700 139.890 ;
        RECT 27.675 139.830 27.965 139.875 ;
        RECT 30.510 139.830 30.650 140.030 ;
        RECT 30.880 139.970 31.200 140.030 ;
        RECT 19.380 139.690 30.650 139.830 ;
        RECT 19.380 139.630 19.700 139.690 ;
        RECT 27.675 139.645 27.965 139.690 ;
        RECT 31.815 139.645 32.105 139.875 ;
        RECT 32.350 139.830 32.490 140.030 ;
        RECT 35.020 139.970 35.340 140.030 ;
        RECT 36.515 139.875 36.655 140.370 ;
        RECT 43.315 140.325 43.605 140.370 ;
        RECT 46.980 140.310 47.300 140.370 ;
        RECT 48.910 140.370 52.730 140.510 ;
        RECT 39.175 140.170 39.465 140.215 ;
        RECT 43.760 140.170 44.080 140.230 ;
        RECT 48.910 140.215 49.050 140.370 ;
        RECT 39.175 140.030 44.080 140.170 ;
        RECT 39.175 139.985 39.465 140.030 ;
        RECT 43.760 139.970 44.080 140.030 ;
        RECT 48.835 139.985 49.125 140.215 ;
        RECT 51.120 139.970 51.440 140.230 ;
        RECT 51.580 139.970 51.900 140.230 ;
        RECT 52.040 139.970 52.360 140.230 ;
        RECT 52.590 140.170 52.730 140.370 ;
        RECT 53.420 140.370 56.485 140.510 ;
        RECT 53.420 140.310 53.740 140.370 ;
        RECT 56.195 140.325 56.485 140.370 ;
        RECT 58.475 140.510 59.125 140.555 ;
        RECT 62.075 140.510 62.365 140.555 ;
        RECT 64.460 140.510 64.780 140.570 ;
        RECT 58.475 140.370 64.780 140.510 ;
        RECT 68.230 140.510 68.370 140.650 ;
        RECT 71.375 140.510 71.665 140.555 ;
        RECT 68.230 140.370 71.665 140.510 ;
        RECT 58.475 140.325 59.125 140.370 ;
        RECT 61.775 140.325 62.365 140.370 ;
        RECT 54.340 140.170 54.660 140.230 ;
        RECT 52.590 140.030 54.660 140.170 ;
        RECT 54.340 139.970 54.660 140.030 ;
        RECT 54.815 139.985 55.105 140.215 ;
        RECT 55.280 140.170 55.570 140.215 ;
        RECT 57.115 140.170 57.405 140.215 ;
        RECT 60.695 140.170 60.985 140.215 ;
        RECT 55.280 140.030 60.985 140.170 ;
        RECT 55.280 139.985 55.570 140.030 ;
        RECT 57.115 139.985 57.405 140.030 ;
        RECT 60.695 139.985 60.985 140.030 ;
        RECT 61.775 140.010 62.065 140.325 ;
        RECT 64.460 140.310 64.780 140.370 ;
        RECT 71.375 140.325 71.665 140.370 ;
        RECT 64.920 140.170 65.240 140.230 ;
        RECT 70.915 140.170 71.205 140.215 ;
        RECT 71.820 140.170 72.140 140.230 ;
        RECT 64.920 140.030 69.750 140.170 ;
        RECT 36.415 139.830 36.705 139.875 ;
        RECT 32.350 139.690 36.705 139.830 ;
        RECT 36.415 139.645 36.705 139.690 ;
        RECT 37.320 139.830 37.640 139.890 ;
        RECT 37.795 139.830 38.085 139.875 ;
        RECT 46.995 139.830 47.285 139.875 ;
        RECT 37.320 139.690 38.085 139.830 ;
        RECT 5.580 139.490 5.900 139.550 ;
        RECT 7.895 139.490 8.185 139.535 ;
        RECT 5.580 139.350 8.185 139.490 ;
        RECT 5.580 139.290 5.900 139.350 ;
        RECT 7.895 139.305 8.185 139.350 ;
        RECT 11.580 139.490 11.870 139.535 ;
        RECT 13.440 139.490 13.730 139.535 ;
        RECT 16.220 139.490 16.510 139.535 ;
        RECT 11.580 139.350 16.510 139.490 ;
        RECT 11.580 139.305 11.870 139.350 ;
        RECT 13.440 139.305 13.730 139.350 ;
        RECT 16.220 139.305 16.510 139.350 ;
        RECT 24.900 139.490 25.220 139.550 ;
        RECT 29.055 139.490 29.345 139.535 ;
        RECT 24.900 139.350 29.345 139.490 ;
        RECT 24.900 139.290 25.220 139.350 ;
        RECT 29.055 139.305 29.345 139.350 ;
        RECT 30.420 139.490 30.740 139.550 ;
        RECT 31.890 139.490 32.030 139.645 ;
        RECT 37.320 139.630 37.640 139.690 ;
        RECT 37.795 139.645 38.085 139.690 ;
        RECT 42.010 139.690 47.285 139.830 ;
        RECT 42.010 139.535 42.150 139.690 ;
        RECT 46.995 139.645 47.285 139.690 ;
        RECT 50.675 139.830 50.965 139.875 ;
        RECT 51.210 139.830 51.350 139.970 ;
        RECT 50.675 139.690 51.350 139.830 ;
        RECT 50.675 139.645 50.965 139.690 ;
        RECT 54.890 139.550 55.030 139.985 ;
        RECT 64.920 139.970 65.240 140.030 ;
        RECT 56.640 139.830 56.960 139.890 ;
        RECT 66.775 139.830 67.065 139.875 ;
        RECT 56.640 139.690 67.065 139.830 ;
        RECT 56.640 139.630 56.960 139.690 ;
        RECT 66.775 139.645 67.065 139.690 ;
        RECT 67.220 139.630 67.540 139.890 ;
        RECT 69.075 139.645 69.365 139.875 ;
        RECT 69.610 139.830 69.750 140.030 ;
        RECT 70.915 140.030 72.140 140.170 ;
        RECT 70.915 139.985 71.205 140.030 ;
        RECT 71.820 139.970 72.140 140.030 ;
        RECT 72.280 140.170 72.600 140.230 ;
        RECT 72.750 140.170 73.040 140.215 ;
        RECT 72.280 140.030 73.040 140.170 ;
        RECT 72.280 139.970 72.600 140.030 ;
        RECT 72.750 139.985 73.040 140.030 ;
        RECT 73.215 139.985 73.505 140.215 ;
        RECT 73.290 139.830 73.430 139.985 ;
        RECT 73.660 139.970 73.980 140.230 ;
        RECT 74.210 140.170 74.350 140.710 ;
        RECT 74.580 140.650 74.900 140.910 ;
        RECT 90.695 140.850 90.985 140.895 ;
        RECT 91.140 140.850 91.460 140.910 ;
        RECT 98.055 140.850 98.345 140.895 ;
        RECT 90.695 140.710 91.460 140.850 ;
        RECT 90.695 140.665 90.985 140.710 ;
        RECT 91.140 140.650 91.460 140.710 ;
        RECT 92.610 140.710 98.345 140.850 ;
        RECT 74.670 140.510 74.810 140.650 ;
        RECT 79.180 140.510 79.500 140.570 ;
        RECT 89.315 140.510 89.605 140.555 ;
        RECT 91.615 140.510 91.905 140.555 ;
        RECT 74.670 140.370 77.570 140.510 ;
        RECT 77.430 140.215 77.570 140.370 ;
        RECT 79.180 140.370 87.690 140.510 ;
        RECT 79.180 140.310 79.500 140.370 ;
        RECT 74.595 140.170 74.885 140.215 ;
        RECT 75.055 140.170 75.345 140.215 ;
        RECT 74.210 140.030 75.345 140.170 ;
        RECT 74.595 139.985 74.885 140.030 ;
        RECT 75.055 139.985 75.345 140.030 ;
        RECT 77.355 139.985 77.645 140.215 ;
        RECT 84.715 140.170 85.005 140.215 ;
        RECT 85.160 140.170 85.480 140.230 ;
        RECT 84.715 140.030 85.480 140.170 ;
        RECT 84.715 139.985 85.005 140.030 ;
        RECT 85.160 139.970 85.480 140.030 ;
        RECT 80.560 139.830 80.880 139.890 ;
        RECT 69.610 139.690 72.965 139.830 ;
        RECT 73.290 139.690 80.880 139.830 ;
        RECT 41.935 139.490 42.225 139.535 ;
        RECT 30.420 139.350 42.225 139.490 ;
        RECT 30.420 139.290 30.740 139.350 ;
        RECT 38.790 139.210 38.930 139.350 ;
        RECT 41.935 139.305 42.225 139.350 ;
        RECT 49.755 139.490 50.045 139.535 ;
        RECT 49.755 139.350 54.570 139.490 ;
        RECT 49.755 139.305 50.045 139.350 ;
        RECT 18.920 139.150 19.240 139.210 ;
        RECT 4.750 139.010 19.240 139.150 ;
        RECT 18.920 138.950 19.240 139.010 ;
        RECT 20.760 138.950 21.080 139.210 ;
        RECT 24.440 138.950 24.760 139.210 ;
        RECT 38.700 138.950 39.020 139.210 ;
        RECT 39.620 139.150 39.940 139.210 ;
        RECT 41.015 139.150 41.305 139.195 ;
        RECT 39.620 139.010 41.305 139.150 ;
        RECT 39.620 138.950 39.940 139.010 ;
        RECT 41.015 138.965 41.305 139.010 ;
        RECT 42.840 139.150 43.160 139.210 ;
        RECT 44.235 139.150 44.525 139.195 ;
        RECT 42.840 139.010 44.525 139.150 ;
        RECT 42.840 138.950 43.160 139.010 ;
        RECT 44.235 138.965 44.525 139.010 ;
        RECT 53.880 138.950 54.200 139.210 ;
        RECT 54.430 139.150 54.570 139.350 ;
        RECT 54.800 139.290 55.120 139.550 ;
        RECT 55.685 139.490 55.975 139.535 ;
        RECT 57.575 139.490 57.865 139.535 ;
        RECT 60.695 139.490 60.985 139.535 ;
        RECT 64.000 139.490 64.320 139.550 ;
        RECT 55.685 139.350 60.985 139.490 ;
        RECT 55.685 139.305 55.975 139.350 ;
        RECT 57.575 139.305 57.865 139.350 ;
        RECT 60.695 139.305 60.985 139.350 ;
        RECT 62.020 139.350 64.320 139.490 ;
        RECT 62.020 139.150 62.160 139.350 ;
        RECT 64.000 139.290 64.320 139.350 ;
        RECT 54.430 139.010 62.160 139.150 ;
        RECT 63.555 139.150 63.845 139.195 ;
        RECT 67.310 139.150 67.450 139.630 ;
        RECT 69.150 139.490 69.290 139.645 ;
        RECT 72.825 139.490 72.965 139.690 ;
        RECT 80.560 139.630 80.880 139.690 ;
        RECT 81.480 139.830 81.800 139.890 ;
        RECT 83.335 139.830 83.625 139.875 ;
        RECT 81.480 139.690 83.625 139.830 ;
        RECT 81.480 139.630 81.800 139.690 ;
        RECT 83.335 139.645 83.625 139.690 ;
        RECT 87.550 139.490 87.690 140.370 ;
        RECT 89.315 140.370 91.905 140.510 ;
        RECT 89.315 140.325 89.605 140.370 ;
        RECT 91.615 140.325 91.905 140.370 ;
        RECT 87.935 139.985 88.225 140.215 ;
        RECT 88.010 139.830 88.150 139.985 ;
        RECT 88.840 139.970 89.160 140.230 ;
        RECT 89.760 140.170 90.080 140.230 ;
        RECT 91.140 140.170 91.460 140.230 ;
        RECT 92.075 140.170 92.365 140.215 ;
        RECT 89.760 140.030 90.910 140.170 ;
        RECT 89.760 139.970 90.080 140.030 ;
        RECT 90.220 139.830 90.540 139.890 ;
        RECT 88.010 139.690 90.540 139.830 ;
        RECT 90.770 139.830 90.910 140.030 ;
        RECT 91.140 140.030 92.365 140.170 ;
        RECT 91.140 139.970 91.460 140.030 ;
        RECT 92.075 139.985 92.365 140.030 ;
        RECT 92.610 139.830 92.750 140.710 ;
        RECT 98.055 140.665 98.345 140.710 ;
        RECT 98.960 140.850 99.280 140.910 ;
        RECT 100.815 140.850 101.105 140.895 ;
        RECT 105.860 140.850 106.180 140.910 ;
        RECT 98.960 140.710 101.105 140.850 ;
        RECT 94.360 140.310 94.680 140.570 ;
        RECT 98.130 140.510 98.270 140.665 ;
        RECT 98.960 140.650 99.280 140.710 ;
        RECT 100.815 140.665 101.105 140.710 ;
        RECT 102.270 140.710 106.180 140.850 ;
        RECT 99.880 140.510 100.200 140.570 ;
        RECT 102.270 140.555 102.410 140.710 ;
        RECT 105.860 140.650 106.180 140.710 ;
        RECT 111.840 140.650 112.160 140.910 ;
        RECT 114.600 140.850 114.920 140.910 ;
        RECT 115.980 140.850 116.300 140.910 ;
        RECT 122.420 140.850 122.740 140.910 ;
        RECT 114.600 140.710 116.300 140.850 ;
        RECT 114.600 140.650 114.920 140.710 ;
        RECT 115.980 140.650 116.300 140.710 ;
        RECT 121.130 140.710 122.740 140.850 ;
        RECT 98.130 140.370 100.200 140.510 ;
        RECT 99.880 140.310 100.200 140.370 ;
        RECT 102.195 140.325 102.485 140.555 ;
        RECT 102.640 140.310 102.960 140.570 ;
        RECT 111.930 140.510 112.070 140.650 ;
        RECT 119.215 140.510 119.505 140.555 ;
        RECT 120.580 140.510 120.900 140.570 ;
        RECT 106.870 140.370 108.850 140.510 ;
        RECT 90.770 139.690 92.750 139.830 ;
        RECT 94.450 139.830 94.590 140.310 ;
        RECT 97.580 140.215 97.900 140.230 ;
        RECT 97.580 139.985 98.050 140.215 ;
        RECT 97.580 139.970 97.900 139.985 ;
        RECT 100.340 139.970 100.660 140.230 ;
        RECT 101.260 140.215 101.580 140.230 ;
        RECT 101.260 139.985 101.795 140.215 ;
        RECT 103.100 140.170 103.420 140.230 ;
        RECT 103.570 140.170 103.860 140.215 ;
        RECT 103.100 140.030 103.860 140.170 ;
        RECT 101.260 139.970 101.580 139.985 ;
        RECT 103.100 139.970 103.420 140.030 ;
        RECT 103.570 139.985 103.860 140.030 ;
        RECT 104.035 140.170 104.325 140.215 ;
        RECT 104.480 140.170 104.800 140.230 ;
        RECT 106.870 140.215 107.010 140.370 ;
        RECT 108.710 140.230 108.850 140.370 ;
        RECT 111.010 140.370 120.900 140.510 ;
        RECT 104.035 140.030 104.800 140.170 ;
        RECT 104.035 139.985 104.325 140.030 ;
        RECT 104.480 139.970 104.800 140.030 ;
        RECT 106.795 139.985 107.085 140.215 ;
        RECT 107.715 139.985 108.005 140.215 ;
        RECT 98.500 139.830 98.820 139.890 ;
        RECT 94.450 139.690 98.820 139.830 ;
        RECT 90.220 139.630 90.540 139.690 ;
        RECT 98.500 139.630 98.820 139.690 ;
        RECT 105.400 139.830 105.720 139.890 ;
        RECT 107.790 139.830 107.930 139.985 ;
        RECT 108.160 139.970 108.480 140.230 ;
        RECT 108.620 139.970 108.940 140.230 ;
        RECT 109.080 139.970 109.400 140.230 ;
        RECT 111.010 140.215 111.150 140.370 ;
        RECT 119.215 140.325 119.505 140.370 ;
        RECT 120.580 140.310 120.900 140.370 ;
        RECT 110.935 139.985 111.225 140.215 ;
        RECT 111.855 140.170 112.145 140.215 ;
        RECT 112.760 140.170 113.080 140.230 ;
        RECT 114.140 140.170 114.460 140.230 ;
        RECT 116.915 140.170 117.205 140.215 ;
        RECT 111.855 140.030 113.910 140.170 ;
        RECT 111.855 139.985 112.145 140.030 ;
        RECT 112.760 139.970 113.080 140.030 ;
        RECT 109.170 139.830 109.310 139.970 ;
        RECT 113.770 139.830 113.910 140.030 ;
        RECT 114.140 140.030 117.205 140.170 ;
        RECT 114.140 139.970 114.460 140.030 ;
        RECT 116.915 139.985 117.205 140.030 ;
        RECT 117.360 139.970 117.680 140.230 ;
        RECT 117.820 140.170 118.140 140.230 ;
        RECT 121.130 140.215 121.270 140.710 ;
        RECT 122.420 140.650 122.740 140.710 ;
        RECT 125.640 140.650 125.960 140.910 ;
        RECT 126.100 140.850 126.420 140.910 ;
        RECT 129.335 140.850 129.625 140.895 ;
        RECT 131.160 140.850 131.480 140.910 ;
        RECT 126.100 140.710 128.630 140.850 ;
        RECT 126.100 140.650 126.420 140.710 ;
        RECT 125.730 140.510 125.870 140.650 ;
        RECT 126.575 140.510 126.865 140.555 ;
        RECT 125.730 140.370 126.865 140.510 ;
        RECT 126.575 140.325 126.865 140.370 ;
        RECT 120.135 140.170 120.425 140.215 ;
        RECT 117.820 140.030 120.425 140.170 ;
        RECT 117.820 139.970 118.140 140.030 ;
        RECT 120.135 139.985 120.425 140.030 ;
        RECT 121.055 139.985 121.345 140.215 ;
        RECT 121.975 140.170 122.265 140.215 ;
        RECT 121.975 140.030 124.030 140.170 ;
        RECT 121.975 139.985 122.265 140.030 ;
        RECT 115.980 139.830 116.300 139.890 ;
        RECT 105.400 139.690 109.310 139.830 ;
        RECT 110.320 139.690 113.450 139.830 ;
        RECT 113.770 139.690 116.300 139.830 ;
        RECT 105.400 139.630 105.720 139.690 ;
        RECT 94.820 139.490 95.140 139.550 ;
        RECT 99.895 139.490 100.185 139.535 ;
        RECT 109.540 139.490 109.860 139.550 ;
        RECT 69.150 139.350 72.510 139.490 ;
        RECT 72.825 139.350 84.470 139.490 ;
        RECT 87.550 139.350 95.140 139.490 ;
        RECT 63.555 139.010 67.450 139.150 ;
        RECT 69.075 139.150 69.365 139.195 ;
        RECT 71.360 139.150 71.680 139.210 ;
        RECT 69.075 139.010 71.680 139.150 ;
        RECT 72.370 139.150 72.510 139.350 ;
        RECT 72.740 139.150 73.060 139.210 ;
        RECT 72.370 139.010 73.060 139.150 ;
        RECT 63.555 138.965 63.845 139.010 ;
        RECT 69.075 138.965 69.365 139.010 ;
        RECT 71.360 138.950 71.680 139.010 ;
        RECT 72.740 138.950 73.060 139.010 ;
        RECT 75.040 139.150 75.360 139.210 ;
        RECT 78.275 139.150 78.565 139.195 ;
        RECT 75.040 139.010 78.565 139.150 ;
        RECT 75.040 138.950 75.360 139.010 ;
        RECT 78.275 138.965 78.565 139.010 ;
        RECT 82.855 139.150 83.145 139.195 ;
        RECT 83.775 139.150 84.065 139.195 ;
        RECT 82.855 139.010 84.065 139.150 ;
        RECT 84.330 139.150 84.470 139.350 ;
        RECT 94.820 139.290 95.140 139.350 ;
        RECT 96.520 139.350 97.810 139.490 ;
        RECT 96.520 139.150 96.660 139.350 ;
        RECT 84.330 139.010 96.660 139.150 ;
        RECT 82.855 138.965 83.145 139.010 ;
        RECT 83.775 138.965 84.065 139.010 ;
        RECT 97.120 138.950 97.440 139.210 ;
        RECT 97.670 139.150 97.810 139.350 ;
        RECT 99.895 139.350 109.860 139.490 ;
        RECT 99.895 139.305 100.185 139.350 ;
        RECT 109.540 139.290 109.860 139.350 ;
        RECT 101.260 139.150 101.580 139.210 ;
        RECT 97.670 139.010 101.580 139.150 ;
        RECT 101.260 138.950 101.580 139.010 ;
        RECT 102.640 139.150 102.960 139.210 ;
        RECT 110.320 139.150 110.460 139.690 ;
        RECT 111.380 139.490 111.700 139.550 ;
        RECT 112.775 139.490 113.065 139.535 ;
        RECT 111.380 139.350 113.065 139.490 ;
        RECT 113.310 139.490 113.450 139.690 ;
        RECT 115.980 139.630 116.300 139.690 ;
        RECT 116.440 139.630 116.760 139.890 ;
        RECT 117.450 139.830 117.590 139.970 ;
        RECT 121.500 139.830 121.820 139.890 ;
        RECT 117.450 139.690 121.820 139.830 ;
        RECT 121.500 139.630 121.820 139.690 ;
        RECT 122.880 139.630 123.200 139.890 ;
        RECT 123.890 139.830 124.030 140.030 ;
        RECT 124.260 139.970 124.580 140.230 ;
        RECT 125.195 139.985 125.485 140.215 ;
        RECT 125.660 140.170 125.950 140.215 ;
        RECT 126.100 140.170 126.420 140.230 ;
        RECT 127.940 140.215 128.260 140.230 ;
        RECT 125.660 140.030 126.420 140.170 ;
        RECT 125.660 139.985 125.950 140.030 ;
        RECT 124.720 139.830 125.040 139.890 ;
        RECT 123.890 139.690 125.040 139.830 ;
        RECT 124.720 139.630 125.040 139.690 ;
        RECT 125.270 139.490 125.410 139.985 ;
        RECT 126.100 139.970 126.420 140.030 ;
        RECT 127.035 139.985 127.325 140.215 ;
        RECT 127.725 139.985 128.260 140.215 ;
        RECT 127.110 139.830 127.250 139.985 ;
        RECT 127.940 139.970 128.260 139.985 ;
        RECT 128.490 139.830 128.630 140.710 ;
        RECT 129.335 140.710 131.480 140.850 ;
        RECT 129.335 140.665 129.625 140.710 ;
        RECT 131.160 140.650 131.480 140.710 ;
        RECT 132.080 140.650 132.400 140.910 ;
        RECT 142.675 140.850 142.965 140.895 ;
        RECT 144.040 140.850 144.360 140.910 ;
        RECT 144.975 140.850 145.265 140.895 ;
        RECT 142.675 140.710 145.265 140.850 ;
        RECT 142.675 140.665 142.965 140.710 ;
        RECT 132.170 140.510 132.310 140.650 ;
        RECT 140.360 140.510 140.680 140.570 ;
        RECT 142.750 140.510 142.890 140.665 ;
        RECT 144.040 140.650 144.360 140.710 ;
        RECT 144.975 140.665 145.265 140.710 ;
        RECT 146.800 140.650 147.120 140.910 ;
        RECT 132.170 140.370 134.150 140.510 ;
        RECT 128.875 140.120 129.165 140.215 ;
        RECT 129.780 140.120 130.100 140.230 ;
        RECT 128.875 139.985 130.100 140.120 ;
        RECT 130.255 139.985 130.545 140.215 ;
        RECT 130.700 140.170 131.020 140.230 ;
        RECT 134.010 140.215 134.150 140.370 ;
        RECT 139.990 140.370 142.890 140.510 ;
        RECT 133.015 140.170 133.305 140.215 ;
        RECT 130.700 140.030 133.305 140.170 ;
        RECT 128.950 139.980 130.100 139.985 ;
        RECT 129.780 139.970 130.100 139.980 ;
        RECT 130.330 139.830 130.470 139.985 ;
        RECT 130.700 139.970 131.020 140.030 ;
        RECT 133.015 139.985 133.305 140.030 ;
        RECT 133.935 139.985 134.225 140.215 ;
        RECT 134.840 140.170 135.160 140.230 ;
        RECT 139.990 140.215 140.130 140.370 ;
        RECT 140.360 140.310 140.680 140.370 ;
        RECT 135.775 140.170 136.065 140.215 ;
        RECT 134.840 140.030 136.065 140.170 ;
        RECT 134.840 139.970 135.160 140.030 ;
        RECT 135.775 139.985 136.065 140.030 ;
        RECT 139.915 139.985 140.205 140.215 ;
        RECT 142.200 140.170 142.520 140.230 ;
        RECT 146.890 140.170 147.030 140.650 ;
        RECT 147.275 140.170 147.565 140.215 ;
        RECT 142.200 140.030 146.570 140.170 ;
        RECT 146.890 140.030 147.565 140.170 ;
        RECT 142.200 139.970 142.520 140.030 ;
        RECT 127.110 139.690 128.170 139.830 ;
        RECT 128.490 139.690 130.470 139.830 ;
        RECT 132.540 139.830 132.860 139.890 ;
        RECT 134.395 139.830 134.685 139.875 ;
        RECT 132.540 139.690 134.685 139.830 ;
        RECT 113.310 139.350 123.110 139.490 ;
        RECT 111.380 139.290 111.700 139.350 ;
        RECT 112.775 139.305 113.065 139.350 ;
        RECT 102.640 139.010 110.460 139.150 ;
        RECT 110.935 139.150 111.225 139.195 ;
        RECT 114.140 139.150 114.460 139.210 ;
        RECT 114.615 139.150 114.905 139.195 ;
        RECT 110.935 139.010 114.905 139.150 ;
        RECT 102.640 138.950 102.960 139.010 ;
        RECT 110.935 138.965 111.225 139.010 ;
        RECT 114.140 138.950 114.460 139.010 ;
        RECT 114.615 138.965 114.905 139.010 ;
        RECT 115.520 138.950 115.840 139.210 ;
        RECT 117.820 139.150 118.140 139.210 ;
        RECT 118.755 139.150 119.045 139.195 ;
        RECT 117.820 139.010 119.045 139.150 ;
        RECT 117.820 138.950 118.140 139.010 ;
        RECT 118.755 138.965 119.045 139.010 ;
        RECT 122.420 138.950 122.740 139.210 ;
        RECT 122.970 139.150 123.110 139.350 ;
        RECT 125.270 139.350 127.710 139.490 ;
        RECT 125.270 139.210 125.410 139.350 ;
        RECT 127.570 139.210 127.710 139.350 ;
        RECT 123.585 139.150 123.875 139.195 ;
        RECT 122.970 139.010 123.875 139.150 ;
        RECT 123.585 138.965 123.875 139.010 ;
        RECT 125.180 138.950 125.500 139.210 ;
        RECT 127.480 138.950 127.800 139.210 ;
        RECT 128.030 139.150 128.170 139.690 ;
        RECT 132.540 139.630 132.860 139.690 ;
        RECT 134.395 139.645 134.685 139.690 ;
        RECT 135.300 139.830 135.620 139.890 ;
        RECT 137.615 139.830 137.905 139.875 ;
        RECT 144.960 139.830 145.280 139.890 ;
        RECT 135.300 139.690 137.905 139.830 ;
        RECT 135.300 139.630 135.620 139.690 ;
        RECT 137.615 139.645 137.905 139.690 ;
        RECT 140.910 139.690 145.280 139.830 ;
        RECT 128.415 139.490 128.705 139.535 ;
        RECT 133.000 139.490 133.320 139.550 ;
        RECT 128.415 139.350 133.320 139.490 ;
        RECT 128.415 139.305 128.705 139.350 ;
        RECT 133.000 139.290 133.320 139.350 ;
        RECT 133.460 139.490 133.780 139.550 ;
        RECT 140.910 139.535 141.050 139.690 ;
        RECT 144.960 139.630 145.280 139.690 ;
        RECT 140.835 139.490 141.125 139.535 ;
        RECT 133.460 139.350 141.125 139.490 ;
        RECT 133.460 139.290 133.780 139.350 ;
        RECT 140.835 139.305 141.125 139.350 ;
        RECT 143.595 139.490 143.885 139.535 ;
        RECT 145.420 139.490 145.740 139.550 ;
        RECT 143.595 139.350 145.740 139.490 ;
        RECT 146.430 139.490 146.570 140.030 ;
        RECT 147.275 139.985 147.565 140.030 ;
        RECT 146.815 139.490 147.105 139.535 ;
        RECT 146.430 139.350 147.105 139.490 ;
        RECT 143.595 139.305 143.885 139.350 ;
        RECT 145.420 139.290 145.740 139.350 ;
        RECT 146.815 139.305 147.105 139.350 ;
        RECT 129.780 139.150 130.100 139.210 ;
        RECT 128.030 139.010 130.100 139.150 ;
        RECT 129.780 138.950 130.100 139.010 ;
        RECT 130.240 139.150 130.560 139.210 ;
        RECT 131.175 139.150 131.465 139.195 ;
        RECT 130.240 139.010 131.465 139.150 ;
        RECT 130.240 138.950 130.560 139.010 ;
        RECT 131.175 138.965 131.465 139.010 ;
        RECT 132.095 139.150 132.385 139.195 ;
        RECT 132.540 139.150 132.860 139.210 ;
        RECT 132.095 139.010 132.860 139.150 ;
        RECT 132.095 138.965 132.385 139.010 ;
        RECT 132.540 138.950 132.860 139.010 ;
        RECT 142.200 139.150 142.520 139.210 ;
        RECT 142.675 139.150 142.965 139.195 ;
        RECT 142.200 139.010 142.965 139.150 ;
        RECT 142.200 138.950 142.520 139.010 ;
        RECT 142.675 138.965 142.965 139.010 ;
        RECT 143.120 139.150 143.440 139.210 ;
        RECT 144.055 139.150 144.345 139.195 ;
        RECT 143.120 139.010 144.345 139.150 ;
        RECT 143.120 138.950 143.440 139.010 ;
        RECT 144.055 138.965 144.345 139.010 ;
        RECT 144.975 139.150 145.265 139.195 ;
        RECT 147.350 139.150 147.490 139.985 ;
        RECT 148.180 139.970 148.500 140.230 ;
        RECT 144.975 139.010 147.490 139.150 ;
        RECT 144.975 138.965 145.265 139.010 ;
        RECT 147.720 138.950 148.040 139.210 ;
        RECT 2.750 138.330 158.230 138.810 ;
        RECT 23.980 138.130 24.300 138.190 ;
        RECT 13.720 137.990 24.300 138.130 ;
        RECT 5.085 137.790 5.375 137.835 ;
        RECT 6.975 137.790 7.265 137.835 ;
        RECT 10.095 137.790 10.385 137.835 ;
        RECT 5.085 137.650 10.385 137.790 ;
        RECT 5.085 137.605 5.375 137.650 ;
        RECT 6.975 137.605 7.265 137.650 ;
        RECT 10.095 137.605 10.385 137.650 ;
        RECT 4.200 137.250 4.520 137.510 ;
        RECT 11.560 137.450 11.880 137.510 ;
        RECT 11.190 137.310 11.880 137.450 ;
        RECT 4.680 137.110 4.970 137.155 ;
        RECT 6.515 137.110 6.805 137.155 ;
        RECT 10.095 137.110 10.385 137.155 ;
        RECT 11.190 137.130 11.330 137.310 ;
        RECT 11.560 137.250 11.880 137.310 ;
        RECT 4.680 136.970 10.385 137.110 ;
        RECT 4.680 136.925 4.970 136.970 ;
        RECT 6.515 136.925 6.805 136.970 ;
        RECT 10.095 136.925 10.385 136.970 ;
        RECT 5.580 136.570 5.900 136.830 ;
        RECT 11.175 136.815 11.465 137.130 ;
        RECT 12.020 137.110 12.340 137.170 ;
        RECT 13.720 137.110 13.860 137.990 ;
        RECT 23.980 137.930 24.300 137.990 ;
        RECT 30.895 138.130 31.185 138.175 ;
        RECT 34.100 138.130 34.420 138.190 ;
        RECT 37.780 138.130 38.100 138.190 ;
        RECT 30.895 137.990 34.420 138.130 ;
        RECT 30.895 137.945 31.185 137.990 ;
        RECT 34.100 137.930 34.420 137.990 ;
        RECT 34.650 137.990 38.100 138.130 ;
        RECT 14.320 137.790 14.640 137.850 ;
        RECT 23.025 137.790 23.315 137.835 ;
        RECT 24.915 137.790 25.205 137.835 ;
        RECT 28.035 137.790 28.325 137.835 ;
        RECT 14.320 137.650 22.370 137.790 ;
        RECT 14.320 137.590 14.640 137.650 ;
        RECT 19.380 137.250 19.700 137.510 ;
        RECT 20.760 137.250 21.080 137.510 ;
        RECT 22.230 137.495 22.370 137.650 ;
        RECT 23.025 137.650 28.325 137.790 ;
        RECT 23.025 137.605 23.315 137.650 ;
        RECT 24.915 137.605 25.205 137.650 ;
        RECT 28.035 137.605 28.325 137.650 ;
        RECT 32.275 137.790 32.565 137.835 ;
        RECT 34.650 137.790 34.790 137.990 ;
        RECT 37.780 137.930 38.100 137.990 ;
        RECT 39.160 138.130 39.480 138.190 ;
        RECT 47.440 138.130 47.760 138.190 ;
        RECT 39.160 137.990 47.760 138.130 ;
        RECT 39.160 137.930 39.480 137.990 ;
        RECT 47.440 137.930 47.760 137.990 ;
        RECT 51.580 137.930 51.900 138.190 ;
        RECT 53.435 138.130 53.725 138.175 ;
        RECT 59.320 138.130 59.610 138.175 ;
        RECT 53.435 137.990 59.610 138.130 ;
        RECT 53.435 137.945 53.725 137.990 ;
        RECT 59.320 137.945 59.610 137.990 ;
        RECT 69.765 138.130 70.055 138.175 ;
        RECT 81.495 138.130 81.785 138.175 ;
        RECT 69.765 137.990 81.785 138.130 ;
        RECT 69.765 137.945 70.055 137.990 ;
        RECT 81.495 137.945 81.785 137.990 ;
        RECT 83.780 138.130 84.100 138.190 ;
        RECT 88.395 138.130 88.685 138.175 ;
        RECT 83.780 137.990 96.890 138.130 ;
        RECT 83.780 137.930 84.100 137.990 ;
        RECT 88.395 137.945 88.685 137.990 ;
        RECT 32.275 137.650 34.790 137.790 ;
        RECT 35.135 137.790 35.425 137.835 ;
        RECT 38.255 137.790 38.545 137.835 ;
        RECT 40.145 137.790 40.435 137.835 ;
        RECT 35.135 137.650 40.435 137.790 ;
        RECT 32.275 137.605 32.565 137.650 ;
        RECT 35.135 137.605 35.425 137.650 ;
        RECT 38.255 137.605 38.545 137.650 ;
        RECT 40.145 137.605 40.435 137.650 ;
        RECT 43.725 137.790 44.015 137.835 ;
        RECT 45.615 137.790 45.905 137.835 ;
        RECT 48.735 137.790 49.025 137.835 ;
        RECT 43.725 137.650 49.025 137.790 ;
        RECT 43.725 137.605 44.015 137.650 ;
        RECT 45.615 137.605 45.905 137.650 ;
        RECT 48.735 137.605 49.025 137.650 ;
        RECT 54.800 137.790 55.120 137.850 ;
        RECT 58.905 137.790 59.195 137.835 ;
        RECT 60.795 137.790 61.085 137.835 ;
        RECT 63.915 137.790 64.205 137.835 ;
        RECT 54.800 137.650 58.250 137.790 ;
        RECT 54.800 137.590 55.120 137.650 ;
        RECT 22.155 137.450 22.445 137.495 ;
        RECT 23.980 137.450 24.300 137.510 ;
        RECT 22.155 137.310 24.300 137.450 ;
        RECT 22.155 137.265 22.445 137.310 ;
        RECT 23.980 137.250 24.300 137.310 ;
        RECT 46.060 137.450 46.380 137.510 ;
        RECT 57.115 137.450 57.405 137.495 ;
        RECT 57.560 137.450 57.880 137.510 ;
        RECT 58.110 137.495 58.250 137.650 ;
        RECT 58.905 137.650 64.205 137.790 ;
        RECT 58.905 137.605 59.195 137.650 ;
        RECT 60.795 137.605 61.085 137.650 ;
        RECT 63.915 137.605 64.205 137.650 ;
        RECT 66.760 137.590 67.080 137.850 ;
        RECT 70.900 137.590 71.220 137.850 ;
        RECT 73.200 137.790 73.520 137.850 ;
        RECT 79.195 137.790 79.485 137.835 ;
        RECT 80.560 137.790 80.880 137.850 ;
        RECT 72.370 137.650 80.880 137.790 ;
        RECT 46.060 137.310 50.430 137.450 ;
        RECT 46.060 137.250 46.380 137.310 ;
        RECT 12.020 136.970 13.860 137.110 ;
        RECT 15.255 137.110 15.545 137.155 ;
        RECT 18.475 137.110 18.765 137.155 ;
        RECT 20.850 137.110 20.990 137.250 ;
        RECT 15.255 136.970 16.390 137.110 ;
        RECT 12.020 136.910 12.340 136.970 ;
        RECT 15.255 136.925 15.545 136.970 ;
        RECT 7.875 136.770 8.525 136.815 ;
        RECT 11.175 136.770 11.765 136.815 ;
        RECT 7.875 136.630 11.765 136.770 ;
        RECT 7.875 136.585 8.525 136.630 ;
        RECT 11.475 136.585 11.765 136.630 ;
        RECT 12.020 136.430 12.340 136.490 ;
        RECT 12.955 136.430 13.245 136.475 ;
        RECT 12.020 136.290 13.245 136.430 ;
        RECT 12.020 136.230 12.340 136.290 ;
        RECT 12.955 136.245 13.245 136.290 ;
        RECT 14.320 136.230 14.640 136.490 ;
        RECT 16.250 136.475 16.390 136.970 ;
        RECT 18.475 136.970 20.990 137.110 ;
        RECT 22.620 137.110 22.910 137.155 ;
        RECT 24.455 137.110 24.745 137.155 ;
        RECT 28.035 137.110 28.325 137.155 ;
        RECT 22.620 136.970 28.325 137.110 ;
        RECT 18.475 136.925 18.765 136.970 ;
        RECT 22.620 136.925 22.910 136.970 ;
        RECT 24.455 136.925 24.745 136.970 ;
        RECT 28.035 136.925 28.325 136.970 ;
        RECT 23.520 136.570 23.840 136.830 ;
        RECT 29.115 136.815 29.405 137.130 ;
        RECT 29.960 137.110 30.280 137.170 ;
        RECT 29.960 136.970 32.950 137.110 ;
        RECT 29.960 136.910 30.280 136.970 ;
        RECT 25.815 136.770 26.465 136.815 ;
        RECT 29.115 136.770 29.705 136.815 ;
        RECT 30.880 136.770 31.200 136.830 ;
        RECT 25.815 136.630 31.200 136.770 ;
        RECT 25.815 136.585 26.465 136.630 ;
        RECT 29.415 136.585 29.705 136.630 ;
        RECT 16.175 136.245 16.465 136.475 ;
        RECT 16.620 136.430 16.940 136.490 ;
        RECT 18.015 136.430 18.305 136.475 ;
        RECT 16.620 136.290 18.305 136.430 ;
        RECT 16.620 136.230 16.940 136.290 ;
        RECT 18.015 136.245 18.305 136.290 ;
        RECT 20.300 136.430 20.620 136.490 ;
        RECT 30.050 136.430 30.190 136.630 ;
        RECT 30.880 136.570 31.200 136.630 ;
        RECT 20.300 136.290 30.190 136.430 ;
        RECT 32.810 136.430 32.950 136.970 ;
        RECT 34.055 136.815 34.345 137.130 ;
        RECT 35.135 137.110 35.425 137.155 ;
        RECT 38.715 137.110 39.005 137.155 ;
        RECT 40.550 137.110 40.840 137.155 ;
        RECT 35.135 136.970 40.840 137.110 ;
        RECT 35.135 136.925 35.425 136.970 ;
        RECT 38.715 136.925 39.005 136.970 ;
        RECT 40.550 136.925 40.840 136.970 ;
        RECT 41.015 137.110 41.305 137.155 ;
        RECT 42.855 137.110 43.145 137.155 ;
        RECT 41.015 136.970 43.145 137.110 ;
        RECT 41.015 136.925 41.305 136.970 ;
        RECT 42.855 136.925 43.145 136.970 ;
        RECT 43.320 137.110 43.610 137.155 ;
        RECT 45.155 137.110 45.445 137.155 ;
        RECT 48.735 137.110 49.025 137.155 ;
        RECT 43.320 136.970 49.025 137.110 ;
        RECT 43.320 136.925 43.610 136.970 ;
        RECT 45.155 136.925 45.445 136.970 ;
        RECT 48.735 136.925 49.025 136.970 ;
        RECT 33.755 136.770 34.345 136.815 ;
        RECT 35.940 136.770 36.260 136.830 ;
        RECT 36.995 136.770 37.645 136.815 ;
        RECT 33.755 136.630 37.645 136.770 ;
        RECT 33.755 136.585 34.045 136.630 ;
        RECT 35.940 136.570 36.260 136.630 ;
        RECT 36.995 136.585 37.645 136.630 ;
        RECT 39.160 136.770 39.480 136.830 ;
        RECT 39.635 136.770 39.925 136.815 ;
        RECT 39.160 136.630 39.925 136.770 ;
        RECT 39.160 136.570 39.480 136.630 ;
        RECT 39.635 136.585 39.925 136.630 ;
        RECT 40.080 136.770 40.400 136.830 ;
        RECT 41.090 136.770 41.230 136.925 ;
        RECT 40.080 136.630 41.230 136.770 ;
        RECT 40.080 136.570 40.400 136.630 ;
        RECT 44.220 136.570 44.540 136.830 ;
        RECT 49.815 136.815 50.105 137.130 ;
        RECT 50.290 136.815 50.430 137.310 ;
        RECT 52.155 137.310 55.950 137.450 ;
        RECT 46.515 136.770 47.165 136.815 ;
        RECT 49.815 136.770 50.430 136.815 ;
        RECT 51.580 136.770 51.900 136.830 ;
        RECT 46.515 136.630 51.900 136.770 ;
        RECT 46.515 136.585 47.165 136.630 ;
        RECT 50.115 136.585 50.405 136.630 ;
        RECT 51.580 136.570 51.900 136.630 ;
        RECT 52.155 136.430 52.295 137.310 ;
        RECT 55.810 137.155 55.950 137.310 ;
        RECT 57.115 137.310 57.880 137.450 ;
        RECT 57.115 137.265 57.405 137.310 ;
        RECT 57.560 137.250 57.880 137.310 ;
        RECT 58.035 137.450 58.325 137.495 ;
        RECT 62.620 137.450 62.940 137.510 ;
        RECT 58.035 137.310 62.940 137.450 ;
        RECT 58.035 137.265 58.325 137.310 ;
        RECT 62.620 137.250 62.940 137.310 ;
        RECT 52.515 137.110 52.805 137.155 ;
        RECT 52.515 136.970 54.110 137.110 ;
        RECT 52.515 136.925 52.805 136.970 ;
        RECT 53.970 136.475 54.110 136.970 ;
        RECT 55.735 136.925 56.025 137.155 ;
        RECT 58.500 137.110 58.790 137.155 ;
        RECT 60.335 137.110 60.625 137.155 ;
        RECT 63.915 137.110 64.205 137.155 ;
        RECT 58.500 136.970 64.205 137.110 ;
        RECT 58.500 136.925 58.790 136.970 ;
        RECT 60.335 136.925 60.625 136.970 ;
        RECT 63.915 136.925 64.205 136.970 ;
        RECT 64.460 137.110 64.780 137.170 ;
        RECT 64.995 137.110 65.285 137.130 ;
        RECT 64.460 136.970 65.285 137.110 ;
        RECT 55.810 136.770 55.950 136.925 ;
        RECT 64.460 136.910 64.780 136.970 ;
        RECT 58.940 136.770 59.260 136.830 ;
        RECT 64.995 136.815 65.285 136.970 ;
        RECT 55.810 136.630 59.260 136.770 ;
        RECT 58.940 136.570 59.260 136.630 ;
        RECT 61.695 136.770 62.345 136.815 ;
        RECT 64.995 136.770 65.585 136.815 ;
        RECT 61.695 136.630 65.585 136.770 ;
        RECT 61.695 136.585 62.345 136.630 ;
        RECT 65.295 136.585 65.585 136.630 ;
        RECT 32.810 136.290 52.295 136.430 ;
        RECT 20.300 136.230 20.620 136.290 ;
        RECT 53.895 136.245 54.185 136.475 ;
        RECT 55.720 136.430 56.040 136.490 ;
        RECT 56.195 136.430 56.485 136.475 ;
        RECT 66.850 136.430 66.990 137.590 ;
        RECT 72.370 137.495 72.510 137.650 ;
        RECT 73.200 137.590 73.520 137.650 ;
        RECT 79.195 137.605 79.485 137.650 ;
        RECT 80.560 137.590 80.880 137.650 ;
        RECT 84.240 137.790 84.560 137.850 ;
        RECT 96.215 137.790 96.505 137.835 ;
        RECT 84.240 137.650 89.070 137.790 ;
        RECT 84.240 137.590 84.560 137.650 ;
        RECT 68.155 137.450 68.445 137.495 ;
        RECT 68.155 137.310 72.050 137.450 ;
        RECT 68.155 137.265 68.445 137.310 ;
        RECT 69.150 137.155 69.290 137.310 ;
        RECT 68.615 136.925 68.905 137.155 ;
        RECT 69.075 136.925 69.365 137.155 ;
        RECT 68.690 136.770 68.830 136.925 ;
        RECT 70.440 136.910 70.760 137.170 ;
        RECT 71.360 136.910 71.680 137.170 ;
        RECT 71.910 137.110 72.050 137.310 ;
        RECT 72.295 137.265 72.585 137.495 ;
        RECT 76.420 137.450 76.740 137.510 ;
        RECT 84.715 137.450 85.005 137.495 ;
        RECT 85.620 137.450 85.940 137.510 ;
        RECT 86.555 137.450 86.845 137.495 ;
        RECT 72.830 137.310 75.270 137.450 ;
        RECT 72.830 137.110 72.970 137.310 ;
        RECT 71.910 136.970 72.970 137.110 ;
        RECT 73.145 137.110 73.435 137.155 ;
        RECT 74.580 137.110 74.900 137.170 ;
        RECT 73.145 136.970 74.900 137.110 ;
        RECT 75.130 137.110 75.270 137.310 ;
        RECT 76.420 137.310 81.710 137.450 ;
        RECT 76.420 137.250 76.740 137.310 ;
        RECT 78.720 137.110 79.040 137.170 ;
        RECT 80.115 137.110 80.405 137.155 ;
        RECT 75.130 136.970 79.040 137.110 ;
        RECT 73.145 136.925 73.435 136.970 ;
        RECT 74.580 136.910 74.900 136.970 ;
        RECT 78.720 136.910 79.040 136.970 ;
        RECT 79.270 136.970 80.405 137.110 ;
        RECT 74.670 136.770 74.810 136.910 ;
        RECT 77.355 136.770 77.645 136.815 ;
        RECT 68.690 136.630 70.210 136.770 ;
        RECT 74.670 136.630 77.645 136.770 ;
        RECT 70.070 136.490 70.210 136.630 ;
        RECT 77.355 136.585 77.645 136.630 ;
        RECT 55.720 136.290 66.990 136.430 ;
        RECT 55.720 136.230 56.040 136.290 ;
        RECT 56.195 136.245 56.485 136.290 ;
        RECT 69.980 136.230 70.300 136.490 ;
        RECT 74.595 136.430 74.885 136.475 ;
        RECT 76.880 136.430 77.200 136.490 ;
        RECT 79.270 136.430 79.410 136.970 ;
        RECT 80.115 136.925 80.405 136.970 ;
        RECT 80.575 137.110 80.865 137.155 ;
        RECT 81.020 137.110 81.340 137.170 ;
        RECT 80.575 136.970 81.340 137.110 ;
        RECT 80.575 136.925 80.865 136.970 ;
        RECT 81.020 136.910 81.340 136.970 ;
        RECT 81.570 136.815 81.710 137.310 ;
        RECT 84.715 137.310 86.845 137.450 ;
        RECT 84.715 137.265 85.005 137.310 ;
        RECT 85.620 137.250 85.940 137.310 ;
        RECT 86.555 137.265 86.845 137.310 ;
        RECT 84.255 137.110 84.545 137.155 ;
        RECT 85.160 137.110 85.480 137.170 ;
        RECT 88.930 137.155 89.070 137.650 ;
        RECT 91.690 137.650 96.505 137.790 ;
        RECT 90.220 137.250 90.540 137.510 ;
        RECT 91.690 137.495 91.830 137.650 ;
        RECT 96.215 137.605 96.505 137.650 ;
        RECT 91.615 137.265 91.905 137.495 ;
        RECT 92.060 137.250 92.380 137.510 ;
        RECT 84.255 136.970 85.480 137.110 ;
        RECT 84.255 136.925 84.545 136.970 ;
        RECT 85.160 136.910 85.480 136.970 ;
        RECT 88.855 137.110 89.145 137.155 ;
        RECT 88.855 136.970 90.450 137.110 ;
        RECT 88.855 136.925 89.145 136.970 ;
        RECT 81.495 136.770 81.785 136.815 ;
        RECT 90.310 136.770 90.450 136.970 ;
        RECT 90.680 136.910 91.000 137.170 ;
        RECT 91.155 137.110 91.445 137.155 ;
        RECT 92.150 137.110 92.290 137.250 ;
        RECT 91.155 136.970 92.290 137.110 ;
        RECT 96.750 137.110 96.890 137.990 ;
        RECT 98.040 137.930 98.360 138.190 ;
        RECT 104.955 138.130 105.245 138.175 ;
        RECT 108.620 138.130 108.940 138.190 ;
        RECT 104.955 137.990 108.940 138.130 ;
        RECT 104.955 137.945 105.245 137.990 ;
        RECT 108.620 137.930 108.940 137.990 ;
        RECT 111.380 137.930 111.700 138.190 ;
        RECT 113.695 138.130 113.985 138.175 ;
        RECT 117.835 138.130 118.125 138.175 ;
        RECT 121.040 138.130 121.360 138.190 ;
        RECT 113.695 137.990 114.830 138.130 ;
        RECT 113.695 137.945 113.985 137.990 ;
        RECT 98.500 137.790 98.820 137.850 ;
        RECT 98.500 137.650 104.250 137.790 ;
        RECT 98.500 137.590 98.820 137.650 ;
        RECT 97.120 137.450 97.440 137.510 ;
        RECT 104.110 137.495 104.250 137.650 ;
        RECT 105.400 137.590 105.720 137.850 ;
        RECT 108.160 137.590 108.480 137.850 ;
        RECT 104.035 137.450 104.325 137.495 ;
        RECT 105.490 137.450 105.630 137.590 ;
        RECT 97.120 137.310 99.190 137.450 ;
        RECT 97.120 137.250 97.440 137.310 ;
        RECT 97.595 137.110 97.885 137.155 ;
        RECT 98.500 137.110 98.820 137.170 ;
        RECT 99.050 137.155 99.190 137.310 ;
        RECT 104.035 137.310 105.630 137.450 ;
        RECT 104.035 137.265 104.325 137.310 ;
        RECT 96.750 136.970 97.350 137.110 ;
        RECT 91.155 136.925 91.445 136.970 ;
        RECT 96.660 136.770 96.980 136.830 ;
        RECT 79.730 136.630 81.250 136.770 ;
        RECT 79.730 136.475 79.870 136.630 ;
        RECT 74.595 136.290 79.410 136.430 ;
        RECT 74.595 136.245 74.885 136.290 ;
        RECT 76.880 136.230 77.200 136.290 ;
        RECT 79.655 136.245 79.945 136.475 ;
        RECT 81.110 136.430 81.250 136.630 ;
        RECT 81.495 136.630 89.530 136.770 ;
        RECT 90.310 136.630 96.980 136.770 ;
        RECT 81.495 136.585 81.785 136.630 ;
        RECT 82.400 136.430 82.720 136.490 ;
        RECT 81.110 136.290 82.720 136.430 ;
        RECT 82.400 136.230 82.720 136.290 ;
        RECT 86.080 136.230 86.400 136.490 ;
        RECT 89.390 136.475 89.530 136.630 ;
        RECT 96.660 136.570 96.980 136.630 ;
        RECT 89.315 136.245 89.605 136.475 ;
        RECT 96.200 136.430 96.520 136.490 ;
        RECT 97.210 136.430 97.350 136.970 ;
        RECT 97.595 136.970 98.820 137.110 ;
        RECT 97.595 136.925 97.885 136.970 ;
        RECT 98.500 136.910 98.820 136.970 ;
        RECT 98.975 136.925 99.265 137.155 ;
        RECT 105.415 137.110 105.705 137.155 ;
        RECT 108.250 137.110 108.390 137.590 ;
        RECT 109.555 137.450 109.845 137.495 ;
        RECT 110.460 137.450 110.780 137.510 ;
        RECT 109.555 137.310 110.780 137.450 ;
        RECT 111.470 137.450 111.610 137.930 ;
        RECT 114.690 137.450 114.830 137.990 ;
        RECT 117.835 137.990 121.360 138.130 ;
        RECT 117.835 137.945 118.125 137.990 ;
        RECT 121.040 137.930 121.360 137.990 ;
        RECT 124.720 137.930 125.040 138.190 ;
        RECT 126.575 138.130 126.865 138.175 ;
        RECT 128.860 138.130 129.180 138.190 ;
        RECT 126.575 137.990 129.180 138.130 ;
        RECT 126.575 137.945 126.865 137.990 ;
        RECT 128.860 137.930 129.180 137.990 ;
        RECT 129.780 138.130 130.100 138.190 ;
        RECT 132.540 138.130 132.860 138.190 ;
        RECT 129.780 137.990 132.860 138.130 ;
        RECT 129.780 137.930 130.100 137.990 ;
        RECT 132.540 137.930 132.860 137.990 ;
        RECT 133.460 138.130 133.780 138.190 ;
        RECT 136.235 138.130 136.525 138.175 ;
        RECT 143.120 138.130 143.440 138.190 ;
        RECT 133.460 137.990 136.525 138.130 ;
        RECT 133.460 137.930 133.780 137.990 ;
        RECT 136.235 137.945 136.525 137.990 ;
        RECT 136.770 137.990 143.440 138.130 ;
        RECT 115.060 137.790 115.380 137.850 ;
        RECT 119.215 137.790 119.505 137.835 ;
        RECT 121.960 137.790 122.280 137.850 ;
        RECT 115.060 137.650 119.505 137.790 ;
        RECT 115.060 137.590 115.380 137.650 ;
        RECT 119.215 137.605 119.505 137.650 ;
        RECT 119.750 137.650 122.280 137.790 ;
        RECT 116.440 137.450 116.760 137.510 ;
        RECT 119.750 137.450 119.890 137.650 ;
        RECT 121.960 137.590 122.280 137.650 ;
        RECT 123.800 137.590 124.120 137.850 ;
        RECT 124.810 137.790 124.950 137.930 ;
        RECT 127.495 137.790 127.785 137.835 ;
        RECT 124.810 137.650 127.785 137.790 ;
        RECT 127.495 137.605 127.785 137.650 ;
        RECT 124.275 137.450 124.565 137.495 ;
        RECT 127.955 137.450 128.245 137.495 ;
        RECT 111.470 137.310 113.450 137.450 ;
        RECT 114.690 137.310 119.890 137.450 ;
        RECT 120.670 137.310 124.030 137.450 ;
        RECT 109.555 137.265 109.845 137.310 ;
        RECT 110.460 137.250 110.780 137.310 ;
        RECT 109.095 137.110 109.385 137.155 ;
        RECT 110.935 137.110 111.225 137.155 ;
        RECT 105.415 136.970 108.390 137.110 ;
        RECT 108.710 136.970 109.385 137.110 ;
        RECT 105.415 136.925 105.705 136.970 ;
        RECT 101.260 136.770 101.580 136.830 ;
        RECT 105.875 136.770 106.165 136.815 ;
        RECT 101.260 136.630 106.165 136.770 ;
        RECT 101.260 136.570 101.580 136.630 ;
        RECT 105.875 136.585 106.165 136.630 ;
        RECT 108.710 136.490 108.850 136.970 ;
        RECT 109.095 136.925 109.385 136.970 ;
        RECT 110.320 136.970 111.225 137.110 ;
        RECT 110.320 136.770 110.460 136.970 ;
        RECT 110.935 136.925 111.225 136.970 ;
        RECT 111.840 137.110 112.160 137.170 ;
        RECT 113.310 137.155 113.450 137.310 ;
        RECT 116.440 137.250 116.760 137.310 ;
        RECT 111.840 136.970 112.990 137.110 ;
        RECT 111.840 136.910 112.160 136.970 ;
        RECT 109.170 136.630 110.460 136.770 ;
        RECT 109.170 136.490 109.310 136.630 ;
        RECT 102.180 136.430 102.500 136.490 ;
        RECT 96.200 136.290 102.500 136.430 ;
        RECT 96.200 136.230 96.520 136.290 ;
        RECT 102.180 136.230 102.500 136.290 ;
        RECT 102.640 136.230 102.960 136.490 ;
        RECT 108.620 136.230 108.940 136.490 ;
        RECT 109.080 136.230 109.400 136.490 ;
        RECT 112.300 136.230 112.620 136.490 ;
        RECT 112.850 136.430 112.990 136.970 ;
        RECT 113.235 136.925 113.525 137.155 ;
        RECT 114.140 136.910 114.460 137.170 ;
        RECT 114.600 137.110 114.920 137.170 ;
        RECT 119.290 137.155 120.350 137.160 ;
        RECT 120.670 137.155 120.810 137.310 ;
        RECT 115.075 137.110 115.365 137.155 ;
        RECT 114.600 136.970 115.365 137.110 ;
        RECT 114.600 136.910 114.920 136.970 ;
        RECT 115.075 136.925 115.365 136.970 ;
        RECT 115.535 137.110 115.825 137.155 ;
        RECT 119.290 137.110 120.425 137.155 ;
        RECT 115.535 137.020 120.425 137.110 ;
        RECT 115.535 136.970 119.430 137.020 ;
        RECT 115.535 136.925 115.825 136.970 ;
        RECT 120.135 136.925 120.425 137.020 ;
        RECT 120.595 136.925 120.885 137.155 ;
        RECT 114.230 136.770 114.370 136.910 ;
        RECT 115.610 136.770 115.750 136.925 ;
        RECT 114.230 136.630 115.750 136.770 ;
        RECT 115.980 136.770 116.300 136.830 ;
        RECT 116.455 136.770 116.745 136.815 ;
        RECT 115.980 136.630 116.745 136.770 ;
        RECT 115.980 136.570 116.300 136.630 ;
        RECT 116.455 136.585 116.745 136.630 ;
        RECT 116.900 136.770 117.220 136.830 ;
        RECT 117.375 136.770 117.665 136.815 ;
        RECT 116.900 136.630 117.665 136.770 ;
        RECT 116.900 136.570 117.220 136.630 ;
        RECT 117.375 136.585 117.665 136.630 ;
        RECT 119.200 136.570 119.520 136.830 ;
        RECT 121.960 136.570 122.280 136.830 ;
        RECT 123.890 136.770 124.030 137.310 ;
        RECT 124.275 137.310 128.245 137.450 ;
        RECT 128.950 137.450 129.090 137.930 ;
        RECT 136.770 137.450 136.910 137.990 ;
        RECT 143.120 137.930 143.440 137.990 ;
        RECT 128.950 137.310 134.150 137.450 ;
        RECT 124.275 137.265 124.565 137.310 ;
        RECT 127.955 137.265 128.245 137.310 ;
        RECT 127.020 136.910 127.340 137.170 ;
        RECT 128.415 137.110 128.705 137.155 ;
        RECT 132.095 137.110 132.385 137.155 ;
        RECT 128.415 136.970 132.385 137.110 ;
        RECT 128.415 136.925 128.705 136.970 ;
        RECT 132.095 136.925 132.385 136.970 ;
        RECT 133.000 136.910 133.320 137.170 ;
        RECT 134.010 137.155 134.150 137.310 ;
        RECT 134.470 137.310 136.910 137.450 ;
        RECT 139.915 137.450 140.205 137.495 ;
        RECT 140.360 137.450 140.680 137.510 ;
        RECT 139.915 137.310 140.680 137.450 ;
        RECT 134.470 137.155 134.610 137.310 ;
        RECT 139.915 137.265 140.205 137.310 ;
        RECT 133.935 136.925 134.225 137.155 ;
        RECT 134.395 136.925 134.685 137.155 ;
        RECT 138.995 137.110 139.285 137.155 ;
        RECT 134.930 136.970 139.285 137.110 ;
        RECT 127.110 136.770 127.250 136.910 ;
        RECT 129.335 136.770 129.625 136.815 ;
        RECT 123.890 136.630 126.790 136.770 ;
        RECT 127.110 136.630 129.625 136.770 ;
        RECT 119.660 136.430 119.980 136.490 ;
        RECT 112.850 136.290 119.980 136.430 ;
        RECT 122.050 136.430 122.190 136.570 ;
        RECT 124.735 136.430 125.025 136.475 ;
        RECT 122.050 136.290 125.025 136.430 ;
        RECT 126.650 136.430 126.790 136.630 ;
        RECT 129.335 136.585 129.625 136.630 ;
        RECT 129.780 136.770 130.100 136.830 ;
        RECT 133.460 136.770 133.780 136.830 ;
        RECT 129.780 136.630 133.780 136.770 ;
        RECT 129.780 136.570 130.100 136.630 ;
        RECT 133.460 136.570 133.780 136.630 ;
        RECT 134.930 136.490 135.070 136.970 ;
        RECT 138.995 136.925 139.285 136.970 ;
        RECT 136.235 136.770 136.525 136.815 ;
        RECT 136.680 136.770 137.000 136.830 ;
        RECT 136.235 136.630 137.000 136.770 ;
        RECT 136.235 136.585 136.525 136.630 ;
        RECT 136.680 136.570 137.000 136.630 ;
        RECT 137.155 136.770 137.445 136.815 ;
        RECT 139.990 136.770 140.130 137.265 ;
        RECT 140.360 137.250 140.680 137.310 ;
        RECT 141.370 137.310 147.950 137.450 ;
        RECT 141.370 137.155 141.510 137.310 ;
        RECT 147.810 137.170 147.950 137.310 ;
        RECT 141.295 136.925 141.585 137.155 ;
        RECT 141.740 137.110 142.060 137.170 ;
        RECT 142.215 137.110 142.505 137.155 ;
        RECT 145.420 137.110 145.740 137.170 ;
        RECT 147.275 137.110 147.565 137.155 ;
        RECT 141.740 136.970 144.960 137.110 ;
        RECT 141.740 136.910 142.060 136.970 ;
        RECT 142.215 136.925 142.505 136.970 ;
        RECT 137.155 136.630 140.130 136.770 ;
        RECT 137.155 136.585 137.445 136.630 ;
        RECT 140.360 136.570 140.680 136.830 ;
        RECT 144.820 136.770 144.960 136.970 ;
        RECT 145.420 136.970 147.565 137.110 ;
        RECT 145.420 136.910 145.740 136.970 ;
        RECT 147.275 136.925 147.565 136.970 ;
        RECT 147.720 136.910 148.040 137.170 ;
        RECT 145.895 136.770 146.185 136.815 ;
        RECT 144.820 136.630 146.185 136.770 ;
        RECT 145.895 136.585 146.185 136.630 ;
        RECT 146.815 136.770 147.105 136.815 ;
        RECT 147.810 136.770 147.950 136.910 ;
        RECT 146.815 136.630 147.950 136.770 ;
        RECT 146.815 136.585 147.105 136.630 ;
        RECT 134.840 136.430 135.160 136.490 ;
        RECT 126.650 136.290 135.160 136.430 ;
        RECT 119.660 136.230 119.980 136.290 ;
        RECT 124.735 136.245 125.025 136.290 ;
        RECT 134.840 136.230 135.160 136.290 ;
        RECT 135.315 136.430 135.605 136.475 ;
        RECT 135.760 136.430 136.080 136.490 ;
        RECT 135.315 136.290 136.080 136.430 ;
        RECT 135.315 136.245 135.605 136.290 ;
        RECT 135.760 136.230 136.080 136.290 ;
        RECT 138.060 136.230 138.380 136.490 ;
        RECT 141.280 136.430 141.600 136.490 ;
        RECT 144.975 136.430 145.265 136.475 ;
        RECT 141.280 136.290 145.265 136.430 ;
        RECT 141.280 136.230 141.600 136.290 ;
        RECT 144.975 136.245 145.265 136.290 ;
        RECT 148.180 136.230 148.500 136.490 ;
        RECT 2.750 135.610 159.030 136.090 ;
        RECT 5.120 135.210 5.440 135.470 ;
        RECT 5.595 135.410 5.885 135.455 ;
        RECT 6.040 135.410 6.360 135.470 ;
        RECT 5.595 135.270 6.360 135.410 ;
        RECT 5.595 135.225 5.885 135.270 ;
        RECT 6.040 135.210 6.360 135.270 ;
        RECT 8.340 135.210 8.660 135.470 ;
        RECT 10.195 135.410 10.485 135.455 ;
        RECT 12.940 135.410 13.260 135.470 ;
        RECT 10.195 135.270 13.260 135.410 ;
        RECT 10.195 135.225 10.485 135.270 ;
        RECT 12.940 135.210 13.260 135.270 ;
        RECT 14.320 135.210 14.640 135.470 ;
        RECT 21.235 135.410 21.525 135.455 ;
        RECT 23.060 135.410 23.380 135.470 ;
        RECT 21.235 135.270 23.380 135.410 ;
        RECT 21.235 135.225 21.525 135.270 ;
        RECT 23.060 135.210 23.380 135.270 ;
        RECT 24.455 135.225 24.745 135.455 ;
        RECT 4.675 134.730 4.965 134.775 ;
        RECT 5.210 134.730 5.350 135.210 ;
        RECT 4.675 134.590 5.350 134.730 ;
        RECT 6.975 134.730 7.265 134.775 ;
        RECT 8.430 134.730 8.570 135.210 ;
        RECT 10.640 135.070 10.960 135.130 ;
        RECT 13.400 135.070 13.720 135.130 ;
        RECT 10.640 134.930 13.720 135.070 ;
        RECT 10.640 134.870 10.960 134.930 ;
        RECT 12.020 134.730 12.340 134.790 ;
        RECT 12.570 134.775 12.710 134.930 ;
        RECT 13.400 134.870 13.720 134.930 ;
        RECT 13.875 135.070 14.165 135.115 ;
        RECT 14.410 135.070 14.550 135.210 ;
        RECT 13.875 134.930 14.550 135.070 ;
        RECT 16.155 135.070 16.805 135.115 ;
        RECT 19.755 135.070 20.045 135.115 ;
        RECT 20.300 135.070 20.620 135.130 ;
        RECT 16.155 134.930 20.620 135.070 ;
        RECT 13.875 134.885 14.165 134.930 ;
        RECT 16.155 134.885 16.805 134.930 ;
        RECT 19.455 134.885 20.045 134.930 ;
        RECT 6.975 134.590 8.570 134.730 ;
        RECT 10.730 134.590 12.340 134.730 ;
        RECT 4.675 134.545 4.965 134.590 ;
        RECT 6.975 134.545 7.265 134.590 ;
        RECT 10.730 134.435 10.870 134.590 ;
        RECT 12.020 134.530 12.340 134.590 ;
        RECT 12.495 134.545 12.785 134.775 ;
        RECT 12.960 134.730 13.250 134.775 ;
        RECT 14.795 134.730 15.085 134.775 ;
        RECT 18.375 134.730 18.665 134.775 ;
        RECT 12.960 134.590 18.665 134.730 ;
        RECT 12.960 134.545 13.250 134.590 ;
        RECT 14.795 134.545 15.085 134.590 ;
        RECT 18.375 134.545 18.665 134.590 ;
        RECT 19.455 134.570 19.745 134.885 ;
        RECT 20.300 134.870 20.620 134.930 ;
        RECT 23.075 134.730 23.365 134.775 ;
        RECT 24.530 134.730 24.670 135.225 ;
        RECT 26.280 135.210 26.600 135.470 ;
        RECT 37.320 135.410 37.640 135.470 ;
        RECT 30.510 135.270 37.640 135.410 ;
        RECT 29.960 135.070 30.280 135.130 ;
        RECT 23.075 134.590 24.670 134.730 ;
        RECT 26.370 134.930 30.280 135.070 ;
        RECT 23.075 134.545 23.365 134.590 ;
        RECT 10.655 134.205 10.945 134.435 ;
        RECT 11.575 134.390 11.865 134.435 ;
        RECT 16.620 134.390 16.940 134.450 ;
        RECT 26.370 134.390 26.510 134.930 ;
        RECT 29.960 134.870 30.280 134.930 ;
        RECT 26.755 134.730 27.045 134.775 ;
        RECT 29.040 134.730 29.360 134.790 ;
        RECT 26.755 134.590 29.360 134.730 ;
        RECT 26.755 134.545 27.045 134.590 ;
        RECT 29.040 134.530 29.360 134.590 ;
        RECT 11.575 134.250 13.170 134.390 ;
        RECT 11.575 134.205 11.865 134.250 ;
        RECT 4.660 133.850 4.980 134.110 ;
        RECT 5.120 134.050 5.440 134.110 ;
        RECT 8.355 134.050 8.645 134.095 ;
        RECT 5.120 133.910 8.645 134.050 ;
        RECT 5.120 133.850 5.440 133.910 ;
        RECT 8.355 133.865 8.645 133.910 ;
        RECT 4.750 133.710 4.890 133.850 ;
        RECT 13.030 133.770 13.170 134.250 ;
        RECT 16.620 134.250 26.510 134.390 ;
        RECT 27.675 134.390 27.965 134.435 ;
        RECT 30.510 134.390 30.650 135.270 ;
        RECT 37.320 135.210 37.640 135.270 ;
        RECT 37.780 135.410 38.100 135.470 ;
        RECT 40.555 135.410 40.845 135.455 ;
        RECT 44.680 135.410 45.000 135.470 ;
        RECT 37.780 135.270 45.000 135.410 ;
        RECT 37.780 135.210 38.100 135.270 ;
        RECT 40.555 135.225 40.845 135.270 ;
        RECT 44.680 135.210 45.000 135.270 ;
        RECT 53.420 135.210 53.740 135.470 ;
        RECT 54.800 135.210 55.120 135.470 ;
        RECT 59.400 135.410 59.720 135.470 ;
        RECT 70.440 135.410 70.760 135.470 ;
        RECT 72.755 135.410 73.045 135.455 ;
        RECT 59.400 135.270 66.530 135.410 ;
        RECT 59.400 135.210 59.720 135.270 ;
        RECT 30.895 135.070 31.185 135.115 ;
        RECT 32.720 135.070 33.040 135.130 ;
        RECT 35.940 135.115 36.260 135.130 ;
        RECT 30.895 134.930 33.040 135.070 ;
        RECT 30.895 134.885 31.185 134.930 ;
        RECT 32.720 134.870 33.040 134.930 ;
        RECT 35.475 135.070 36.260 135.115 ;
        RECT 39.075 135.070 39.365 135.115 ;
        RECT 35.475 134.930 39.365 135.070 ;
        RECT 35.475 134.885 36.260 134.930 ;
        RECT 35.940 134.870 36.260 134.885 ;
        RECT 38.775 134.885 39.365 134.930 ;
        RECT 43.415 135.070 43.705 135.115 ;
        RECT 46.060 135.070 46.380 135.130 ;
        RECT 46.655 135.070 47.305 135.115 ;
        RECT 54.890 135.070 55.030 135.210 ;
        RECT 59.855 135.070 60.505 135.115 ;
        RECT 63.455 135.070 63.745 135.115 ;
        RECT 43.415 134.930 47.305 135.070 ;
        RECT 43.415 134.885 44.005 134.930 ;
        RECT 32.280 134.730 32.570 134.775 ;
        RECT 34.115 134.730 34.405 134.775 ;
        RECT 37.695 134.730 37.985 134.775 ;
        RECT 32.280 134.590 37.985 134.730 ;
        RECT 32.280 134.545 32.570 134.590 ;
        RECT 34.115 134.545 34.405 134.590 ;
        RECT 37.695 134.545 37.985 134.590 ;
        RECT 38.775 134.570 39.065 134.885 ;
        RECT 43.715 134.570 44.005 134.885 ;
        RECT 46.060 134.870 46.380 134.930 ;
        RECT 46.655 134.885 47.305 134.930 ;
        RECT 50.750 134.930 56.410 135.070 ;
        RECT 50.750 134.775 50.890 134.930 ;
        RECT 56.270 134.790 56.410 134.930 ;
        RECT 59.855 134.930 63.745 135.070 ;
        RECT 59.855 134.885 60.505 134.930 ;
        RECT 63.155 134.885 63.745 134.930 ;
        RECT 63.155 134.790 63.445 134.885 ;
        RECT 44.795 134.730 45.085 134.775 ;
        RECT 48.375 134.730 48.665 134.775 ;
        RECT 50.210 134.730 50.500 134.775 ;
        RECT 44.795 134.590 50.500 134.730 ;
        RECT 44.795 134.545 45.085 134.590 ;
        RECT 48.375 134.545 48.665 134.590 ;
        RECT 50.210 134.545 50.500 134.590 ;
        RECT 50.675 134.545 50.965 134.775 ;
        RECT 52.040 134.530 52.360 134.790 ;
        RECT 52.515 134.730 52.805 134.775 ;
        RECT 53.880 134.730 54.200 134.790 ;
        RECT 52.515 134.590 54.200 134.730 ;
        RECT 52.515 134.545 52.805 134.590 ;
        RECT 53.880 134.530 54.200 134.590 ;
        RECT 54.800 134.530 55.120 134.790 ;
        RECT 56.180 134.530 56.500 134.790 ;
        RECT 56.660 134.730 56.950 134.775 ;
        RECT 58.495 134.730 58.785 134.775 ;
        RECT 62.075 134.730 62.365 134.775 ;
        RECT 56.660 134.590 62.365 134.730 ;
        RECT 56.660 134.545 56.950 134.590 ;
        RECT 58.495 134.545 58.785 134.590 ;
        RECT 62.075 134.545 62.365 134.590 ;
        RECT 63.080 134.570 63.445 134.790 ;
        RECT 66.390 134.775 66.530 135.270 ;
        RECT 70.440 135.270 73.045 135.410 ;
        RECT 70.440 135.210 70.760 135.270 ;
        RECT 72.755 135.225 73.045 135.270 ;
        RECT 73.660 135.410 73.980 135.470 ;
        RECT 75.055 135.410 75.345 135.455 ;
        RECT 75.960 135.410 76.280 135.470 ;
        RECT 73.660 135.270 75.345 135.410 ;
        RECT 73.660 135.210 73.980 135.270 ;
        RECT 75.055 135.225 75.345 135.270 ;
        RECT 75.590 135.270 76.280 135.410 ;
        RECT 69.520 134.870 69.840 135.130 ;
        RECT 75.590 135.070 75.730 135.270 ;
        RECT 75.960 135.210 76.280 135.270 ;
        RECT 76.420 135.210 76.740 135.470 ;
        RECT 76.880 135.210 77.200 135.470 ;
        RECT 77.340 135.410 77.660 135.470 ;
        RECT 77.340 135.270 78.030 135.410 ;
        RECT 77.340 135.210 77.660 135.270 ;
        RECT 74.670 134.930 75.730 135.070 ;
        RECT 63.080 134.530 63.400 134.570 ;
        RECT 66.315 134.545 66.605 134.775 ;
        RECT 72.280 134.530 72.600 134.790 ;
        RECT 73.200 134.530 73.520 134.790 ;
        RECT 74.670 134.775 74.810 134.930 ;
        RECT 73.675 134.545 73.965 134.775 ;
        RECT 74.595 134.545 74.885 134.775 ;
        RECT 75.975 134.730 76.265 134.775 ;
        RECT 76.510 134.730 76.650 135.210 ;
        RECT 76.970 135.070 77.110 135.210 ;
        RECT 76.970 134.930 77.570 135.070 ;
        RECT 75.975 134.590 76.650 134.730 ;
        RECT 75.975 134.545 76.265 134.590 ;
        RECT 27.675 134.250 30.650 134.390 ;
        RECT 16.620 134.190 16.940 134.250 ;
        RECT 27.675 134.205 27.965 134.250 ;
        RECT 31.815 134.205 32.105 134.435 ;
        RECT 13.365 134.050 13.655 134.095 ;
        RECT 15.255 134.050 15.545 134.095 ;
        RECT 18.375 134.050 18.665 134.095 ;
        RECT 13.365 133.910 18.665 134.050 ;
        RECT 13.365 133.865 13.655 133.910 ;
        RECT 15.255 133.865 15.545 133.910 ;
        RECT 18.375 133.865 18.665 133.910 ;
        RECT 19.380 134.050 19.700 134.110 ;
        RECT 31.890 134.050 32.030 134.205 ;
        RECT 33.180 134.190 33.500 134.450 ;
        RECT 35.020 134.390 35.340 134.450 ;
        RECT 49.295 134.390 49.585 134.435 ;
        RECT 57.575 134.390 57.865 134.435 ;
        RECT 35.020 134.250 43.990 134.390 ;
        RECT 35.020 134.190 35.340 134.250 ;
        RECT 43.850 134.110 43.990 134.250 ;
        RECT 49.295 134.250 51.350 134.390 ;
        RECT 49.295 134.205 49.585 134.250 ;
        RECT 19.380 133.910 32.030 134.050 ;
        RECT 32.685 134.050 32.975 134.095 ;
        RECT 34.575 134.050 34.865 134.095 ;
        RECT 37.695 134.050 37.985 134.095 ;
        RECT 32.685 133.910 37.985 134.050 ;
        RECT 19.380 133.850 19.700 133.910 ;
        RECT 32.685 133.865 32.975 133.910 ;
        RECT 34.575 133.865 34.865 133.910 ;
        RECT 37.695 133.865 37.985 133.910 ;
        RECT 43.760 133.850 44.080 134.110 ;
        RECT 51.210 134.095 51.350 134.250 ;
        RECT 55.810 134.250 57.865 134.390 ;
        RECT 55.810 134.095 55.950 134.250 ;
        RECT 57.575 134.205 57.865 134.250 ;
        RECT 69.535 134.205 69.825 134.435 ;
        RECT 44.795 134.050 45.085 134.095 ;
        RECT 47.915 134.050 48.205 134.095 ;
        RECT 49.805 134.050 50.095 134.095 ;
        RECT 44.795 133.910 50.095 134.050 ;
        RECT 44.795 133.865 45.085 133.910 ;
        RECT 47.915 133.865 48.205 133.910 ;
        RECT 49.805 133.865 50.095 133.910 ;
        RECT 51.135 133.865 51.425 134.095 ;
        RECT 55.735 133.865 56.025 134.095 ;
        RECT 57.065 134.050 57.355 134.095 ;
        RECT 58.955 134.050 59.245 134.095 ;
        RECT 62.075 134.050 62.365 134.095 ;
        RECT 57.065 133.910 62.365 134.050 ;
        RECT 57.065 133.865 57.355 133.910 ;
        RECT 58.955 133.865 59.245 133.910 ;
        RECT 62.075 133.865 62.365 133.910 ;
        RECT 64.920 133.850 65.240 134.110 ;
        RECT 65.380 133.850 65.700 134.110 ;
        RECT 65.840 134.050 66.160 134.110 ;
        RECT 67.235 134.050 67.525 134.095 ;
        RECT 65.840 133.910 67.525 134.050 ;
        RECT 65.840 133.850 66.160 133.910 ;
        RECT 67.235 133.865 67.525 133.910 ;
        RECT 6.055 133.710 6.345 133.755 ;
        RECT 4.750 133.570 6.345 133.710 ;
        RECT 6.055 133.525 6.345 133.570 ;
        RECT 12.940 133.510 13.260 133.770 ;
        RECT 23.060 133.710 23.380 133.770 ;
        RECT 23.995 133.710 24.285 133.755 ;
        RECT 23.060 133.570 24.285 133.710 ;
        RECT 23.060 133.510 23.380 133.570 ;
        RECT 23.995 133.525 24.285 133.570 ;
        RECT 30.435 133.710 30.725 133.755 ;
        RECT 30.880 133.710 31.200 133.770 ;
        RECT 35.020 133.710 35.340 133.770 ;
        RECT 30.435 133.570 35.340 133.710 ;
        RECT 30.435 133.525 30.725 133.570 ;
        RECT 30.880 133.510 31.200 133.570 ;
        RECT 35.020 133.510 35.340 133.570 ;
        RECT 41.935 133.710 42.225 133.755 ;
        RECT 46.980 133.710 47.300 133.770 ;
        RECT 41.935 133.570 47.300 133.710 ;
        RECT 69.610 133.710 69.750 134.205 ;
        RECT 69.980 134.190 70.300 134.450 ;
        RECT 72.370 134.390 72.510 134.530 ;
        RECT 73.750 134.390 73.890 134.545 ;
        RECT 76.880 134.530 77.200 134.790 ;
        RECT 77.430 134.775 77.570 134.930 ;
        RECT 77.890 134.775 78.030 135.270 ;
        RECT 78.720 135.210 79.040 135.470 ;
        RECT 83.780 135.210 84.100 135.470 ;
        RECT 84.240 135.210 84.560 135.470 ;
        RECT 85.620 135.210 85.940 135.470 ;
        RECT 87.935 135.410 88.225 135.455 ;
        RECT 88.840 135.410 89.160 135.470 ;
        RECT 87.935 135.270 89.160 135.410 ;
        RECT 87.935 135.225 88.225 135.270 ;
        RECT 88.840 135.210 89.160 135.270 ;
        RECT 90.220 135.210 90.540 135.470 ;
        RECT 90.680 135.210 91.000 135.470 ;
        RECT 91.600 135.410 91.920 135.470 ;
        RECT 109.080 135.410 109.400 135.470 ;
        RECT 91.600 135.270 109.400 135.410 ;
        RECT 91.600 135.210 91.920 135.270 ;
        RECT 109.080 135.210 109.400 135.270 ;
        RECT 109.540 135.210 109.860 135.470 ;
        RECT 115.060 135.410 115.380 135.470 ;
        RECT 111.930 135.270 115.380 135.410 ;
        RECT 77.355 134.545 77.645 134.775 ;
        RECT 77.815 134.545 78.105 134.775 ;
        RECT 80.575 134.545 80.865 134.775 ;
        RECT 81.495 134.545 81.785 134.775 ;
        RECT 83.870 134.730 84.010 135.210 ;
        RECT 84.330 135.070 84.470 135.210 ;
        RECT 85.175 135.070 85.465 135.115 ;
        RECT 84.330 134.930 85.465 135.070 ;
        RECT 85.175 134.885 85.465 134.930 ;
        RECT 85.710 134.775 85.850 135.210 ;
        RECT 86.080 135.070 86.400 135.130 ;
        RECT 90.310 135.070 90.450 135.210 ;
        RECT 91.155 135.070 91.445 135.115 ;
        RECT 103.115 135.070 103.405 135.115 ;
        RECT 105.860 135.070 106.180 135.130 ;
        RECT 86.080 134.930 89.070 135.070 ;
        RECT 90.310 134.930 91.445 135.070 ;
        RECT 86.080 134.870 86.400 134.930 ;
        RECT 88.930 134.775 89.070 134.930 ;
        RECT 91.155 134.885 91.445 134.930 ;
        RECT 95.370 134.930 103.405 135.070 ;
        RECT 84.255 134.730 84.545 134.775 ;
        RECT 83.870 134.590 84.545 134.730 ;
        RECT 84.255 134.545 84.545 134.590 ;
        RECT 85.635 134.545 85.925 134.775 ;
        RECT 88.855 134.730 89.145 134.775 ;
        RECT 88.855 134.590 89.990 134.730 ;
        RECT 88.855 134.545 89.145 134.590 ;
        RECT 72.370 134.250 73.890 134.390 ;
        RECT 73.750 134.050 73.890 134.250 ;
        RECT 74.135 134.390 74.425 134.435 ;
        RECT 75.500 134.390 75.820 134.450 ;
        RECT 80.650 134.390 80.790 134.545 ;
        RECT 74.135 134.250 80.790 134.390 ;
        RECT 74.135 134.205 74.425 134.250 ;
        RECT 75.500 134.190 75.820 134.250 ;
        RECT 81.020 134.190 81.340 134.450 ;
        RECT 77.800 134.050 78.120 134.110 ;
        RECT 73.750 133.910 78.120 134.050 ;
        RECT 77.800 133.850 78.120 133.910 ;
        RECT 78.260 134.050 78.580 134.110 ;
        RECT 81.570 134.050 81.710 134.545 ;
        RECT 89.315 134.205 89.605 134.435 ;
        RECT 89.850 134.390 89.990 134.590 ;
        RECT 92.535 134.545 92.825 134.775 ;
        RECT 91.155 134.390 91.445 134.435 ;
        RECT 89.850 134.250 91.445 134.390 ;
        RECT 91.155 134.205 91.445 134.250 ;
        RECT 78.260 133.910 81.710 134.050 ;
        RECT 89.390 134.050 89.530 134.205 ;
        RECT 90.680 134.050 91.000 134.110 ;
        RECT 92.610 134.050 92.750 134.545 ;
        RECT 89.390 133.910 92.750 134.050 ;
        RECT 78.260 133.850 78.580 133.910 ;
        RECT 90.680 133.850 91.000 133.910 ;
        RECT 82.860 133.710 83.180 133.770 ;
        RECT 69.610 133.570 83.180 133.710 ;
        RECT 41.935 133.525 42.225 133.570 ;
        RECT 46.980 133.510 47.300 133.570 ;
        RECT 82.860 133.510 83.180 133.570 ;
        RECT 83.320 133.510 83.640 133.770 ;
        RECT 85.160 133.710 85.480 133.770 ;
        RECT 86.095 133.710 86.385 133.755 ;
        RECT 85.160 133.570 86.385 133.710 ;
        RECT 85.160 133.510 85.480 133.570 ;
        RECT 86.095 133.525 86.385 133.570 ;
        RECT 88.840 133.710 89.160 133.770 ;
        RECT 92.075 133.710 92.365 133.755 ;
        RECT 88.840 133.570 92.365 133.710 ;
        RECT 88.840 133.510 89.160 133.570 ;
        RECT 92.075 133.525 92.365 133.570 ;
        RECT 93.900 133.710 94.220 133.770 ;
        RECT 95.370 133.710 95.510 134.930 ;
        RECT 96.200 134.530 96.520 134.790 ;
        RECT 96.660 134.730 96.980 134.790 ;
        RECT 99.510 134.775 99.650 134.930 ;
        RECT 103.115 134.885 103.405 134.930 ;
        RECT 103.650 134.930 106.180 135.070 ;
        RECT 102.180 134.775 102.500 134.790 ;
        RECT 97.135 134.730 97.425 134.775 ;
        RECT 97.595 134.730 97.885 134.775 ;
        RECT 96.660 134.590 97.885 134.730 ;
        RECT 96.660 134.530 96.980 134.590 ;
        RECT 97.135 134.545 97.425 134.590 ;
        RECT 97.595 134.545 97.885 134.590 ;
        RECT 99.435 134.545 99.725 134.775 ;
        RECT 102.170 134.730 102.500 134.775 ;
        RECT 101.985 134.590 102.500 134.730 ;
        RECT 102.170 134.545 102.500 134.590 ;
        RECT 102.655 134.730 102.945 134.775 ;
        RECT 103.650 134.730 103.790 134.930 ;
        RECT 105.860 134.870 106.180 134.930 ;
        RECT 108.620 134.870 108.940 135.130 ;
        RECT 102.655 134.590 103.790 134.730 ;
        RECT 102.655 134.545 102.945 134.590 ;
        RECT 102.180 134.530 102.500 134.545 ;
        RECT 104.020 134.530 104.340 134.790 ;
        RECT 104.480 134.730 104.800 134.790 ;
        RECT 108.175 134.730 108.465 134.775 ;
        RECT 109.170 134.730 109.310 135.210 ;
        RECT 104.480 134.590 107.930 134.730 ;
        RECT 104.480 134.530 104.800 134.590 ;
        RECT 98.040 134.190 98.360 134.450 ;
        RECT 99.895 134.390 100.185 134.435 ;
        RECT 104.105 134.390 104.245 134.530 ;
        RECT 107.790 134.390 107.930 134.590 ;
        RECT 108.175 134.590 109.310 134.730 ;
        RECT 108.175 134.545 108.465 134.590 ;
        RECT 99.895 134.250 103.790 134.390 ;
        RECT 104.105 134.250 107.010 134.390 ;
        RECT 107.790 134.250 109.310 134.390 ;
        RECT 99.895 134.205 100.185 134.250 ;
        RECT 95.740 134.050 96.060 134.110 ;
        RECT 101.275 134.050 101.565 134.095 ;
        RECT 95.740 133.910 101.565 134.050 ;
        RECT 95.740 133.850 96.060 133.910 ;
        RECT 101.275 133.865 101.565 133.910 ;
        RECT 96.675 133.710 96.965 133.755 ;
        RECT 93.900 133.570 96.965 133.710 ;
        RECT 93.900 133.510 94.220 133.570 ;
        RECT 96.675 133.525 96.965 133.570 ;
        RECT 97.120 133.710 97.440 133.770 ;
        RECT 100.815 133.710 101.105 133.755 ;
        RECT 97.120 133.570 101.105 133.710 ;
        RECT 103.650 133.710 103.790 134.250 ;
        RECT 106.870 134.110 107.010 134.250 ;
        RECT 109.170 134.110 109.310 134.250 ;
        RECT 106.780 133.850 107.100 134.110 ;
        RECT 109.080 133.850 109.400 134.110 ;
        RECT 109.630 134.050 109.770 135.210 ;
        RECT 110.475 134.730 110.765 134.775 ;
        RECT 111.380 134.730 111.700 134.790 ;
        RECT 110.475 134.590 111.700 134.730 ;
        RECT 110.475 134.545 110.765 134.590 ;
        RECT 111.380 134.530 111.700 134.590 ;
        RECT 110.015 134.390 110.305 134.435 ;
        RECT 111.930 134.390 112.070 135.270 ;
        RECT 115.060 135.210 115.380 135.270 ;
        RECT 115.520 135.210 115.840 135.470 ;
        RECT 117.820 135.210 118.140 135.470 ;
        RECT 121.040 135.210 121.360 135.470 ;
        RECT 121.960 135.410 122.280 135.470 ;
        RECT 125.640 135.410 125.960 135.470 ;
        RECT 128.860 135.410 129.180 135.470 ;
        RECT 121.960 135.270 125.960 135.410 ;
        RECT 121.960 135.210 122.280 135.270 ;
        RECT 125.640 135.210 125.960 135.270 ;
        RECT 128.030 135.270 129.180 135.410 ;
        RECT 112.760 135.070 113.080 135.130 ;
        RECT 115.610 135.070 115.750 135.210 ;
        RECT 112.760 134.930 114.830 135.070 ;
        RECT 115.610 134.930 116.670 135.070 ;
        RECT 112.760 134.870 113.080 134.930 ;
        RECT 114.690 134.790 114.830 134.930 ;
        RECT 112.315 134.730 112.605 134.775 ;
        RECT 113.235 134.730 113.525 134.775 ;
        RECT 114.140 134.730 114.460 134.790 ;
        RECT 112.315 134.590 112.990 134.730 ;
        RECT 112.315 134.545 112.605 134.590 ;
        RECT 110.015 134.250 112.070 134.390 ;
        RECT 110.015 134.205 110.305 134.250 ;
        RECT 112.850 134.050 112.990 134.590 ;
        RECT 113.235 134.590 114.460 134.730 ;
        RECT 113.235 134.545 113.525 134.590 ;
        RECT 114.140 134.530 114.460 134.590 ;
        RECT 114.600 134.530 114.920 134.790 ;
        RECT 116.530 134.775 116.670 134.930 ;
        RECT 115.535 134.545 115.825 134.775 ;
        RECT 115.995 134.545 116.285 134.775 ;
        RECT 116.455 134.545 116.745 134.775 ;
        RECT 117.910 134.730 118.050 135.210 ;
        RECT 126.100 135.070 126.420 135.130 ;
        RECT 128.030 135.070 128.170 135.270 ;
        RECT 128.860 135.210 129.180 135.270 ;
        RECT 131.620 135.410 131.940 135.470 ;
        RECT 131.620 135.270 138.750 135.410 ;
        RECT 131.620 135.210 131.940 135.270 ;
        RECT 132.095 135.070 132.385 135.115 ;
        RECT 132.540 135.070 132.860 135.130 ;
        RECT 126.100 134.930 128.170 135.070 ;
        RECT 126.100 134.870 126.420 134.930 ;
        RECT 118.295 134.730 118.585 134.775 ;
        RECT 116.990 134.590 118.585 134.730 ;
        RECT 109.630 133.910 112.990 134.050 ;
        RECT 115.610 134.050 115.750 134.545 ;
        RECT 116.070 134.390 116.210 134.545 ;
        RECT 116.990 134.390 117.130 134.590 ;
        RECT 118.295 134.545 118.585 134.590 ;
        RECT 119.675 134.545 119.965 134.775 ;
        RECT 120.135 134.730 120.425 134.775 ;
        RECT 122.420 134.730 122.740 134.790 ;
        RECT 120.135 134.590 122.740 134.730 ;
        RECT 120.135 134.545 120.425 134.590 ;
        RECT 116.070 134.250 117.130 134.390 ;
        RECT 117.835 134.390 118.125 134.435 ;
        RECT 119.750 134.390 119.890 134.545 ;
        RECT 122.420 134.530 122.740 134.590 ;
        RECT 124.735 134.730 125.025 134.775 ;
        RECT 125.640 134.730 125.960 134.790 ;
        RECT 128.030 134.775 128.170 134.930 ;
        RECT 128.490 134.930 132.860 135.070 ;
        RECT 128.490 134.790 128.630 134.930 ;
        RECT 132.095 134.885 132.385 134.930 ;
        RECT 132.540 134.870 132.860 134.930 ;
        RECT 133.175 135.070 133.465 135.115 ;
        RECT 134.380 135.070 134.700 135.130 ;
        RECT 138.610 135.115 138.750 135.270 ;
        RECT 133.175 134.930 134.700 135.070 ;
        RECT 133.175 134.885 133.465 134.930 ;
        RECT 134.380 134.870 134.700 134.930 ;
        RECT 135.850 134.930 138.290 135.070 ;
        RECT 124.735 134.590 127.250 134.730 ;
        RECT 124.735 134.545 125.025 134.590 ;
        RECT 125.640 134.530 125.960 134.590 ;
        RECT 117.835 134.250 119.890 134.390 ;
        RECT 125.195 134.390 125.485 134.435 ;
        RECT 126.560 134.390 126.880 134.450 ;
        RECT 125.195 134.250 126.880 134.390 ;
        RECT 127.110 134.390 127.250 134.590 ;
        RECT 127.955 134.545 128.245 134.775 ;
        RECT 128.400 134.530 128.720 134.790 ;
        RECT 129.335 134.545 129.625 134.775 ;
        RECT 129.795 134.730 130.085 134.775 ;
        RECT 131.620 134.730 131.940 134.790 ;
        RECT 129.795 134.590 131.940 134.730 ;
        RECT 129.795 134.545 130.085 134.590 ;
        RECT 129.410 134.390 129.550 134.545 ;
        RECT 131.620 134.530 131.940 134.590 ;
        RECT 133.920 134.730 134.240 134.790 ;
        RECT 135.315 134.730 135.605 134.775 ;
        RECT 133.920 134.590 135.605 134.730 ;
        RECT 133.920 134.530 134.240 134.590 ;
        RECT 135.315 134.545 135.605 134.590 ;
        RECT 134.010 134.390 134.150 134.530 ;
        RECT 135.850 134.435 135.990 134.930 ;
        RECT 137.615 134.730 137.905 134.775 ;
        RECT 136.310 134.590 137.905 134.730 ;
        RECT 138.150 134.730 138.290 134.930 ;
        RECT 138.535 134.885 138.825 135.115 ;
        RECT 139.455 134.885 139.745 135.115 ;
        RECT 139.530 134.730 139.670 134.885 ;
        RECT 138.150 134.590 139.670 134.730 ;
        RECT 127.110 134.250 134.150 134.390 ;
        RECT 117.835 134.205 118.125 134.250 ;
        RECT 125.195 134.205 125.485 134.250 ;
        RECT 126.560 134.190 126.880 134.250 ;
        RECT 135.775 134.205 136.065 134.435 ;
        RECT 115.980 134.050 116.300 134.110 ;
        RECT 127.940 134.050 128.260 134.110 ;
        RECT 131.620 134.050 131.940 134.110 ;
        RECT 115.610 133.910 116.300 134.050 ;
        RECT 109.630 133.710 109.770 133.910 ;
        RECT 103.650 133.570 109.770 133.710 ;
        RECT 112.850 133.710 112.990 133.910 ;
        RECT 115.980 133.850 116.300 133.910 ;
        RECT 116.530 133.910 127.710 134.050 ;
        RECT 116.530 133.710 116.670 133.910 ;
        RECT 127.570 133.770 127.710 133.910 ;
        RECT 127.940 133.910 131.940 134.050 ;
        RECT 127.940 133.850 128.260 133.910 ;
        RECT 131.620 133.850 131.940 133.910 ;
        RECT 132.540 134.050 132.860 134.110 ;
        RECT 133.935 134.050 134.225 134.095 ;
        RECT 136.310 134.050 136.450 134.590 ;
        RECT 137.615 134.545 137.905 134.590 ;
        RECT 132.540 133.910 136.450 134.050 ;
        RECT 137.155 134.050 137.445 134.095 ;
        RECT 137.600 134.050 137.920 134.110 ;
        RECT 137.155 133.910 137.920 134.050 ;
        RECT 132.540 133.850 132.860 133.910 ;
        RECT 133.935 133.865 134.225 133.910 ;
        RECT 137.155 133.865 137.445 133.910 ;
        RECT 137.600 133.850 137.920 133.910 ;
        RECT 112.850 133.570 116.670 133.710 ;
        RECT 116.900 133.710 117.220 133.770 ;
        RECT 118.755 133.710 119.045 133.755 ;
        RECT 116.900 133.570 119.045 133.710 ;
        RECT 97.120 133.510 97.440 133.570 ;
        RECT 100.815 133.525 101.105 133.570 ;
        RECT 116.900 133.510 117.220 133.570 ;
        RECT 118.755 133.525 119.045 133.570 ;
        RECT 119.200 133.710 119.520 133.770 ;
        RECT 123.355 133.710 123.645 133.755 ;
        RECT 119.200 133.570 123.645 133.710 ;
        RECT 119.200 133.510 119.520 133.570 ;
        RECT 123.355 133.525 123.645 133.570 ;
        RECT 127.020 133.510 127.340 133.770 ;
        RECT 127.480 133.510 127.800 133.770 ;
        RECT 131.160 133.710 131.480 133.770 ;
        RECT 133.015 133.710 133.305 133.755 ;
        RECT 131.160 133.570 133.305 133.710 ;
        RECT 131.160 133.510 131.480 133.570 ;
        RECT 133.015 133.525 133.305 133.570 ;
        RECT 133.460 133.710 133.780 133.770 ;
        RECT 134.840 133.710 135.160 133.770 ;
        RECT 148.180 133.710 148.500 133.770 ;
        RECT 133.460 133.570 148.500 133.710 ;
        RECT 133.460 133.510 133.780 133.570 ;
        RECT 134.840 133.510 135.160 133.570 ;
        RECT 148.180 133.510 148.500 133.570 ;
        RECT 2.750 132.890 158.230 133.370 ;
        RECT 5.135 132.690 5.425 132.735 ;
        RECT 5.580 132.690 5.900 132.750 ;
        RECT 5.135 132.550 5.900 132.690 ;
        RECT 5.135 132.505 5.425 132.550 ;
        RECT 5.580 132.490 5.900 132.550 ;
        RECT 23.060 132.690 23.380 132.750 ;
        RECT 23.900 132.690 24.190 132.735 ;
        RECT 23.060 132.550 24.190 132.690 ;
        RECT 23.060 132.490 23.380 132.550 ;
        RECT 23.900 132.505 24.190 132.550 ;
        RECT 31.355 132.690 31.645 132.735 ;
        RECT 33.640 132.690 33.960 132.750 ;
        RECT 31.355 132.550 33.960 132.690 ;
        RECT 31.355 132.505 31.645 132.550 ;
        RECT 33.640 132.490 33.960 132.550 ;
        RECT 35.940 132.490 36.260 132.750 ;
        RECT 37.320 132.490 37.640 132.750 ;
        RECT 41.015 132.690 41.305 132.735 ;
        RECT 44.220 132.690 44.540 132.750 ;
        RECT 41.015 132.550 44.540 132.690 ;
        RECT 41.015 132.505 41.305 132.550 ;
        RECT 44.220 132.490 44.540 132.550 ;
        RECT 47.900 132.690 48.220 132.750 ;
        RECT 48.835 132.690 49.125 132.735 ;
        RECT 47.900 132.550 49.125 132.690 ;
        RECT 47.900 132.490 48.220 132.550 ;
        RECT 48.835 132.505 49.125 132.550 ;
        RECT 52.040 132.490 52.360 132.750 ;
        RECT 54.355 132.690 54.645 132.735 ;
        RECT 54.800 132.690 55.120 132.750 ;
        RECT 54.355 132.550 55.120 132.690 ;
        RECT 54.355 132.505 54.645 132.550 ;
        RECT 54.800 132.490 55.120 132.550 ;
        RECT 71.360 132.690 71.680 132.750 ;
        RECT 73.675 132.690 73.965 132.735 ;
        RECT 71.360 132.550 73.965 132.690 ;
        RECT 71.360 132.490 71.680 132.550 ;
        RECT 73.675 132.505 73.965 132.550 ;
        RECT 75.515 132.690 75.805 132.735 ;
        RECT 78.260 132.690 78.580 132.750 ;
        RECT 75.515 132.550 78.580 132.690 ;
        RECT 75.515 132.505 75.805 132.550 ;
        RECT 78.260 132.490 78.580 132.550 ;
        RECT 80.100 132.690 80.420 132.750 ;
        RECT 94.835 132.690 95.125 132.735 ;
        RECT 80.100 132.550 95.125 132.690 ;
        RECT 80.100 132.490 80.420 132.550 ;
        RECT 94.835 132.505 95.125 132.550 ;
        RECT 98.500 132.690 98.820 132.750 ;
        RECT 114.600 132.690 114.920 132.750 ;
        RECT 98.500 132.550 110.690 132.690 ;
        RECT 98.500 132.490 98.820 132.550 ;
        RECT 6.465 132.350 6.755 132.395 ;
        RECT 8.355 132.350 8.645 132.395 ;
        RECT 11.475 132.350 11.765 132.395 ;
        RECT 6.465 132.210 11.765 132.350 ;
        RECT 6.465 132.165 6.755 132.210 ;
        RECT 8.355 132.165 8.645 132.210 ;
        RECT 11.475 132.165 11.765 132.210 ;
        RECT 13.860 132.350 14.180 132.410 ;
        RECT 19.380 132.350 19.700 132.410 ;
        RECT 13.860 132.210 19.700 132.350 ;
        RECT 13.860 132.150 14.180 132.210 ;
        RECT 19.380 132.150 19.700 132.210 ;
        RECT 23.485 132.350 23.775 132.395 ;
        RECT 25.375 132.350 25.665 132.395 ;
        RECT 28.495 132.350 28.785 132.395 ;
        RECT 36.030 132.350 36.170 132.490 ;
        RECT 23.485 132.210 28.785 132.350 ;
        RECT 23.485 132.165 23.775 132.210 ;
        RECT 25.375 132.165 25.665 132.210 ;
        RECT 28.495 132.165 28.785 132.210 ;
        RECT 30.970 132.210 36.170 132.350 ;
        RECT 37.410 132.350 37.550 132.490 ;
        RECT 46.520 132.350 46.840 132.410 ;
        RECT 37.410 132.210 43.990 132.350 ;
        RECT 5.120 131.810 5.440 132.070 ;
        RECT 5.595 132.010 5.885 132.055 ;
        RECT 10.180 132.010 10.500 132.070 ;
        RECT 5.595 131.870 10.500 132.010 ;
        RECT 5.595 131.825 5.885 131.870 ;
        RECT 10.180 131.810 10.500 131.870 ;
        RECT 14.320 132.010 14.640 132.070 ;
        RECT 16.160 132.010 16.480 132.070 ;
        RECT 14.320 131.870 16.480 132.010 ;
        RECT 14.320 131.810 14.640 131.870 ;
        RECT 16.160 131.810 16.480 131.870 ;
        RECT 18.935 132.010 19.225 132.055 ;
        RECT 30.420 132.010 30.740 132.070 ;
        RECT 18.935 131.870 30.740 132.010 ;
        RECT 18.935 131.825 19.225 131.870 ;
        RECT 4.215 131.670 4.505 131.715 ;
        RECT 5.210 131.670 5.350 131.810 ;
        RECT 4.215 131.530 5.350 131.670 ;
        RECT 6.060 131.670 6.350 131.715 ;
        RECT 7.895 131.670 8.185 131.715 ;
        RECT 11.475 131.670 11.765 131.715 ;
        RECT 6.060 131.530 11.765 131.670 ;
        RECT 4.215 131.485 4.505 131.530 ;
        RECT 6.060 131.485 6.350 131.530 ;
        RECT 7.895 131.485 8.185 131.530 ;
        RECT 11.475 131.485 11.765 131.530 ;
        RECT 12.020 131.670 12.340 131.730 ;
        RECT 12.555 131.670 12.845 131.690 ;
        RECT 13.860 131.670 14.180 131.730 ;
        RECT 15.240 131.670 15.560 131.730 ;
        RECT 19.010 131.670 19.150 131.825 ;
        RECT 30.420 131.810 30.740 131.870 ;
        RECT 12.020 131.530 13.630 131.670 ;
        RECT 12.020 131.470 12.340 131.530 ;
        RECT 6.960 131.130 7.280 131.390 ;
        RECT 12.555 131.375 12.845 131.530 ;
        RECT 9.255 131.330 9.905 131.375 ;
        RECT 12.555 131.330 13.145 131.375 ;
        RECT 9.255 131.190 13.145 131.330 ;
        RECT 13.490 131.330 13.630 131.530 ;
        RECT 13.860 131.530 19.150 131.670 ;
        RECT 13.860 131.470 14.180 131.530 ;
        RECT 15.240 131.470 15.560 131.530 ;
        RECT 20.300 131.470 20.620 131.730 ;
        RECT 22.155 131.485 22.445 131.715 ;
        RECT 20.390 131.330 20.530 131.470 ;
        RECT 13.490 131.190 20.530 131.330 ;
        RECT 22.230 131.330 22.370 131.485 ;
        RECT 22.600 131.470 22.920 131.730 ;
        RECT 23.080 131.670 23.370 131.715 ;
        RECT 24.915 131.670 25.205 131.715 ;
        RECT 28.495 131.670 28.785 131.715 ;
        RECT 23.080 131.530 28.785 131.670 ;
        RECT 23.080 131.485 23.370 131.530 ;
        RECT 24.915 131.485 25.205 131.530 ;
        RECT 28.495 131.485 28.785 131.530 ;
        RECT 29.500 131.690 29.820 131.730 ;
        RECT 29.500 131.670 29.865 131.690 ;
        RECT 30.970 131.670 31.110 132.210 ;
        RECT 37.780 132.010 38.100 132.070 ;
        RECT 38.330 132.055 38.470 132.210 ;
        RECT 35.110 131.870 38.100 132.010 ;
        RECT 29.500 131.530 31.110 131.670 ;
        RECT 32.275 131.670 32.565 131.715 ;
        RECT 35.110 131.670 35.250 131.870 ;
        RECT 37.780 131.810 38.100 131.870 ;
        RECT 38.255 131.825 38.545 132.055 ;
        RECT 42.840 132.010 43.160 132.070 ;
        RECT 43.850 132.055 43.990 132.210 ;
        RECT 44.770 132.210 46.840 132.350 ;
        RECT 44.770 132.055 44.910 132.210 ;
        RECT 46.520 132.150 46.840 132.210 ;
        RECT 46.995 132.350 47.285 132.395 ;
        RECT 52.130 132.350 52.270 132.490 ;
        RECT 46.995 132.210 52.270 132.350 ;
        RECT 69.980 132.350 70.300 132.410 ;
        RECT 75.040 132.350 75.360 132.410 ;
        RECT 69.980 132.210 75.360 132.350 ;
        RECT 46.995 132.165 47.285 132.210 ;
        RECT 69.980 132.150 70.300 132.210 ;
        RECT 40.170 131.870 43.160 132.010 ;
        RECT 32.275 131.530 35.250 131.670 ;
        RECT 35.480 131.670 35.800 131.730 ;
        RECT 40.170 131.715 40.310 131.870 ;
        RECT 42.840 131.810 43.160 131.870 ;
        RECT 43.775 131.825 44.065 132.055 ;
        RECT 44.695 131.825 44.985 132.055 ;
        RECT 46.060 132.010 46.380 132.070 ;
        RECT 52.515 132.010 52.805 132.055 ;
        RECT 52.960 132.010 53.280 132.070 ;
        RECT 46.060 131.870 49.970 132.010 ;
        RECT 46.060 131.810 46.380 131.870 ;
        RECT 37.335 131.670 37.625 131.715 ;
        RECT 35.480 131.530 37.625 131.670 ;
        RECT 29.500 131.470 29.865 131.530 ;
        RECT 32.275 131.485 32.565 131.530 ;
        RECT 35.480 131.470 35.800 131.530 ;
        RECT 37.335 131.485 37.625 131.530 ;
        RECT 40.095 131.485 40.385 131.715 ;
        RECT 41.935 131.670 42.225 131.715 ;
        RECT 49.830 131.670 49.970 131.870 ;
        RECT 52.515 131.870 53.280 132.010 ;
        RECT 52.515 131.825 52.805 131.870 ;
        RECT 52.960 131.810 53.280 131.870 ;
        RECT 53.435 132.010 53.725 132.055 ;
        RECT 57.560 132.010 57.880 132.070 ;
        RECT 53.435 131.870 57.880 132.010 ;
        RECT 53.435 131.825 53.725 131.870 ;
        RECT 57.560 131.810 57.880 131.870 ;
        RECT 64.920 131.810 65.240 132.070 ;
        RECT 67.680 132.010 68.000 132.070 ;
        RECT 68.155 132.010 68.445 132.055 ;
        RECT 67.680 131.870 68.445 132.010 ;
        RECT 67.680 131.810 68.000 131.870 ;
        RECT 68.155 131.825 68.445 131.870 ;
        RECT 56.195 131.670 56.485 131.715 ;
        RECT 41.935 131.530 49.510 131.670 ;
        RECT 49.830 131.530 56.485 131.670 ;
        RECT 41.935 131.485 42.225 131.530 ;
        RECT 24.440 131.330 24.760 131.390 ;
        RECT 29.575 131.375 29.865 131.470 ;
        RECT 22.230 131.190 24.760 131.330 ;
        RECT 9.255 131.145 9.905 131.190 ;
        RECT 12.855 131.145 13.145 131.190 ;
        RECT 24.440 131.130 24.760 131.190 ;
        RECT 26.275 131.330 26.925 131.375 ;
        RECT 29.575 131.330 30.165 131.375 ;
        RECT 26.275 131.190 30.165 131.330 ;
        RECT 26.275 131.145 26.925 131.190 ;
        RECT 29.875 131.145 30.165 131.190 ;
        RECT 30.880 131.330 31.200 131.390 ;
        RECT 35.035 131.330 35.325 131.375 ;
        RECT 37.795 131.330 38.085 131.375 ;
        RECT 30.880 131.190 32.030 131.330 ;
        RECT 30.880 131.130 31.200 131.190 ;
        RECT 16.160 130.790 16.480 131.050 ;
        RECT 16.620 130.990 16.940 131.050 ;
        RECT 18.015 130.990 18.305 131.035 ;
        RECT 16.620 130.850 18.305 130.990 ;
        RECT 16.620 130.790 16.940 130.850 ;
        RECT 18.015 130.805 18.305 130.850 ;
        RECT 18.460 130.790 18.780 131.050 ;
        RECT 21.220 130.790 21.540 131.050 ;
        RECT 31.890 130.990 32.030 131.190 ;
        RECT 35.035 131.190 38.085 131.330 ;
        RECT 35.035 131.145 35.325 131.190 ;
        RECT 37.795 131.145 38.085 131.190 ;
        RECT 43.760 131.330 44.080 131.390 ;
        RECT 45.140 131.330 45.460 131.390 ;
        RECT 43.760 131.190 45.460 131.330 ;
        RECT 43.760 131.130 44.080 131.190 ;
        RECT 45.140 131.130 45.460 131.190 ;
        RECT 48.820 131.130 49.140 131.390 ;
        RECT 35.495 130.990 35.785 131.035 ;
        RECT 31.890 130.850 35.785 130.990 ;
        RECT 35.495 130.805 35.785 130.850 ;
        RECT 42.840 130.790 43.160 131.050 ;
        RECT 47.440 130.990 47.760 131.050 ;
        RECT 47.915 130.990 48.205 131.035 ;
        RECT 47.440 130.850 48.205 130.990 ;
        RECT 49.370 130.990 49.510 131.530 ;
        RECT 56.195 131.485 56.485 131.530 ;
        RECT 56.655 131.670 56.945 131.715 ;
        RECT 65.010 131.670 65.150 131.810 ;
        RECT 56.655 131.530 65.150 131.670 ;
        RECT 70.455 131.670 70.745 131.715 ;
        RECT 70.990 131.670 71.130 132.210 ;
        RECT 75.040 132.150 75.360 132.210 ;
        RECT 77.355 132.350 77.645 132.395 ;
        RECT 88.855 132.350 89.145 132.395 ;
        RECT 77.355 132.210 89.145 132.350 ;
        RECT 77.355 132.165 77.645 132.210 ;
        RECT 88.855 132.165 89.145 132.210 ;
        RECT 89.315 132.350 89.605 132.395 ;
        RECT 91.140 132.350 91.460 132.410 ;
        RECT 102.640 132.350 102.960 132.410 ;
        RECT 89.315 132.210 91.460 132.350 ;
        RECT 89.315 132.165 89.605 132.210 ;
        RECT 91.140 132.150 91.460 132.210 ;
        RECT 96.750 132.210 102.960 132.350 ;
        RECT 81.035 132.010 81.325 132.055 ;
        RECT 81.480 132.010 81.800 132.070 ;
        RECT 71.450 131.870 77.570 132.010 ;
        RECT 71.450 131.715 71.590 131.870 ;
        RECT 70.455 131.530 71.130 131.670 ;
        RECT 56.655 131.485 56.945 131.530 ;
        RECT 70.455 131.485 70.745 131.530 ;
        RECT 71.375 131.485 71.665 131.715 ;
        RECT 71.835 131.670 72.125 131.715 ;
        RECT 71.835 131.530 72.510 131.670 ;
        RECT 71.835 131.485 72.125 131.530 ;
        RECT 49.755 131.330 50.045 131.375 ;
        RECT 52.500 131.330 52.820 131.390 ;
        RECT 49.755 131.190 52.820 131.330 ;
        RECT 56.270 131.330 56.410 131.485 ;
        RECT 58.020 131.330 58.340 131.390 ;
        RECT 69.060 131.330 69.380 131.390 ;
        RECT 56.270 131.190 57.330 131.330 ;
        RECT 49.755 131.145 50.045 131.190 ;
        RECT 52.500 131.130 52.820 131.190 ;
        RECT 50.215 130.990 50.505 131.035 ;
        RECT 49.370 130.850 50.505 130.990 ;
        RECT 47.440 130.790 47.760 130.850 ;
        RECT 47.915 130.805 48.205 130.850 ;
        RECT 50.215 130.805 50.505 130.850 ;
        RECT 52.040 130.790 52.360 131.050 ;
        RECT 57.190 130.990 57.330 131.190 ;
        RECT 58.020 131.190 69.380 131.330 ;
        RECT 58.020 131.130 58.340 131.190 ;
        RECT 69.060 131.130 69.380 131.190 ;
        RECT 72.370 131.050 72.510 131.530 ;
        RECT 75.040 131.470 75.360 131.730 ;
        RECT 75.500 131.470 75.820 131.730 ;
        RECT 76.880 131.470 77.200 131.730 ;
        RECT 75.960 131.130 76.280 131.390 ;
        RECT 67.680 130.990 68.000 131.050 ;
        RECT 57.190 130.850 68.000 130.990 ;
        RECT 67.680 130.790 68.000 130.850 ;
        RECT 72.280 130.790 72.600 131.050 ;
        RECT 75.500 130.990 75.820 131.050 ;
        RECT 76.970 130.990 77.110 131.470 ;
        RECT 77.430 131.330 77.570 131.870 ;
        RECT 81.035 131.870 81.800 132.010 ;
        RECT 81.035 131.825 81.325 131.870 ;
        RECT 81.480 131.810 81.800 131.870 ;
        RECT 82.415 132.010 82.705 132.055 ;
        RECT 83.320 132.010 83.640 132.070 ;
        RECT 82.415 131.870 96.430 132.010 ;
        RECT 82.415 131.825 82.705 131.870 ;
        RECT 83.320 131.810 83.640 131.870 ;
        RECT 77.815 131.670 78.105 131.715 ;
        RECT 80.100 131.670 80.420 131.730 ;
        RECT 84.790 131.715 84.930 131.870 ;
        RECT 77.815 131.530 80.420 131.670 ;
        RECT 77.815 131.485 78.105 131.530 ;
        RECT 80.100 131.470 80.420 131.530 ;
        RECT 81.955 131.485 82.245 131.715 ;
        RECT 84.715 131.485 85.005 131.715 ;
        RECT 85.635 131.485 85.925 131.715 ;
        RECT 86.540 131.670 86.860 131.730 ;
        RECT 88.840 131.670 89.160 131.730 ;
        RECT 93.900 131.670 94.220 131.730 ;
        RECT 86.540 131.530 89.160 131.670 ;
        RECT 81.020 131.330 81.340 131.390 ;
        RECT 77.430 131.190 81.340 131.330 ;
        RECT 82.030 131.330 82.170 131.485 ;
        RECT 84.255 131.330 84.545 131.375 ;
        RECT 85.710 131.330 85.850 131.485 ;
        RECT 86.540 131.470 86.860 131.530 ;
        RECT 88.840 131.470 89.160 131.530 ;
        RECT 89.850 131.530 94.220 131.670 ;
        RECT 89.850 131.330 89.990 131.530 ;
        RECT 93.900 131.470 94.220 131.530 ;
        RECT 95.740 131.470 96.060 131.730 ;
        RECT 96.290 131.715 96.430 131.870 ;
        RECT 96.215 131.485 96.505 131.715 ;
        RECT 82.030 131.190 83.550 131.330 ;
        RECT 81.020 131.130 81.340 131.190 ;
        RECT 83.410 131.050 83.550 131.190 ;
        RECT 84.255 131.190 89.990 131.330 ;
        RECT 90.235 131.330 90.525 131.375 ;
        RECT 96.750 131.330 96.890 132.210 ;
        RECT 102.640 132.150 102.960 132.210 ;
        RECT 98.040 132.010 98.360 132.070 ;
        RECT 98.040 131.870 101.030 132.010 ;
        RECT 98.040 131.810 98.360 131.870 ;
        RECT 97.120 131.470 97.440 131.730 ;
        RECT 97.595 131.670 97.885 131.715 ;
        RECT 98.500 131.670 98.820 131.730 ;
        RECT 97.595 131.530 98.820 131.670 ;
        RECT 97.595 131.485 97.885 131.530 ;
        RECT 97.670 131.330 97.810 131.485 ;
        RECT 98.500 131.470 98.820 131.530 ;
        RECT 100.340 131.470 100.660 131.730 ;
        RECT 100.890 131.715 101.030 131.870 ;
        RECT 100.815 131.670 101.105 131.715 ;
        RECT 101.260 131.670 101.580 131.730 ;
        RECT 100.815 131.530 101.580 131.670 ;
        RECT 100.815 131.485 101.105 131.530 ;
        RECT 101.260 131.470 101.580 131.530 ;
        RECT 101.720 131.470 102.040 131.730 ;
        RECT 102.180 131.470 102.500 131.730 ;
        RECT 103.190 131.670 103.330 132.550 ;
        RECT 109.555 131.825 109.845 132.055 ;
        RECT 104.035 131.670 104.325 131.715 ;
        RECT 103.190 131.530 104.325 131.670 ;
        RECT 104.035 131.485 104.325 131.530 ;
        RECT 104.500 131.485 104.790 131.715 ;
        RECT 90.235 131.190 96.890 131.330 ;
        RECT 97.210 131.190 97.810 131.330 ;
        RECT 101.350 131.330 101.490 131.470 ;
        RECT 104.575 131.330 104.715 131.485 ;
        RECT 105.860 131.470 106.180 131.730 ;
        RECT 106.320 131.715 106.640 131.730 ;
        RECT 106.320 131.670 106.650 131.715 ;
        RECT 108.635 131.670 108.925 131.715 ;
        RECT 109.080 131.670 109.400 131.730 ;
        RECT 106.320 131.530 106.835 131.670 ;
        RECT 108.635 131.530 109.400 131.670 ;
        RECT 109.630 131.670 109.770 131.825 ;
        RECT 110.000 131.810 110.320 132.070 ;
        RECT 110.550 132.010 110.690 132.550 ;
        RECT 114.600 132.550 120.350 132.690 ;
        RECT 114.600 132.490 114.920 132.550 ;
        RECT 112.300 132.350 112.620 132.410 ;
        RECT 115.980 132.350 116.300 132.410 ;
        RECT 111.930 132.210 116.300 132.350 ;
        RECT 111.930 132.055 112.070 132.210 ;
        RECT 112.300 132.150 112.620 132.210 ;
        RECT 115.980 132.150 116.300 132.210 ;
        RECT 117.360 132.150 117.680 132.410 ;
        RECT 120.210 132.350 120.350 132.550 ;
        RECT 120.580 132.490 120.900 132.750 ;
        RECT 129.320 132.490 129.640 132.750 ;
        RECT 131.175 132.690 131.465 132.735 ;
        RECT 131.175 132.550 140.590 132.690 ;
        RECT 131.175 132.505 131.465 132.550 ;
        RECT 123.340 132.350 123.660 132.410 ;
        RECT 131.635 132.350 131.925 132.395 ;
        RECT 120.210 132.210 123.660 132.350 ;
        RECT 110.550 131.870 111.610 132.010 ;
        RECT 109.630 131.530 110.230 131.670 ;
        RECT 106.320 131.485 106.650 131.530 ;
        RECT 108.635 131.485 108.925 131.530 ;
        RECT 106.320 131.470 106.640 131.485 ;
        RECT 109.080 131.470 109.400 131.530 ;
        RECT 101.350 131.190 104.715 131.330 ;
        RECT 105.415 131.330 105.705 131.375 ;
        RECT 105.415 131.190 109.310 131.330 ;
        RECT 84.255 131.145 84.545 131.190 ;
        RECT 90.235 131.145 90.525 131.190 ;
        RECT 97.210 131.050 97.350 131.190 ;
        RECT 105.415 131.145 105.705 131.190 ;
        RECT 75.500 130.850 77.110 130.990 ;
        RECT 75.500 130.790 75.820 130.850 ;
        RECT 83.320 130.790 83.640 131.050 ;
        RECT 85.175 130.990 85.465 131.035 ;
        RECT 85.620 130.990 85.940 131.050 ;
        RECT 85.175 130.850 85.940 130.990 ;
        RECT 85.175 130.805 85.465 130.850 ;
        RECT 85.620 130.790 85.940 130.850 ;
        RECT 97.120 130.790 97.440 131.050 ;
        RECT 98.500 130.990 98.820 131.050 ;
        RECT 99.435 130.990 99.725 131.035 ;
        RECT 98.500 130.850 99.725 130.990 ;
        RECT 98.500 130.790 98.820 130.850 ;
        RECT 99.435 130.805 99.725 130.850 ;
        RECT 101.260 130.990 101.580 131.050 ;
        RECT 105.490 130.990 105.630 131.145 ;
        RECT 109.170 131.050 109.310 131.190 ;
        RECT 101.260 130.850 105.630 130.990 ;
        RECT 101.260 130.790 101.580 130.850 ;
        RECT 107.240 130.790 107.560 131.050 ;
        RECT 107.700 130.790 108.020 131.050 ;
        RECT 109.080 130.990 109.400 131.050 ;
        RECT 110.090 130.990 110.230 131.530 ;
        RECT 111.470 131.050 111.610 131.870 ;
        RECT 111.855 131.825 112.145 132.055 ;
        RECT 113.695 132.010 113.985 132.055 ;
        RECT 120.595 132.010 120.885 132.055 ;
        RECT 113.695 131.870 120.885 132.010 ;
        RECT 113.695 131.825 113.985 131.870 ;
        RECT 120.595 131.825 120.885 131.870 ;
        RECT 112.775 131.670 113.065 131.715 ;
        RECT 115.075 131.670 115.365 131.715 ;
        RECT 115.995 131.670 116.285 131.715 ;
        RECT 116.440 131.670 116.760 131.730 ;
        RECT 122.050 131.715 122.190 132.210 ;
        RECT 123.340 132.150 123.660 132.210 ;
        RECT 130.790 132.210 131.925 132.350 ;
        RECT 124.735 132.010 125.025 132.055 ;
        RECT 126.560 132.010 126.880 132.070 ;
        RECT 124.735 131.870 126.880 132.010 ;
        RECT 124.735 131.825 125.025 131.870 ;
        RECT 126.560 131.810 126.880 131.870 ;
        RECT 112.775 131.530 115.750 131.670 ;
        RECT 112.775 131.485 113.065 131.530 ;
        RECT 115.075 131.485 115.365 131.530 ;
        RECT 109.080 130.850 110.230 130.990 ;
        RECT 111.380 130.990 111.700 131.050 ;
        RECT 115.060 130.990 115.380 131.050 ;
        RECT 111.380 130.850 115.380 130.990 ;
        RECT 115.610 130.990 115.750 131.530 ;
        RECT 115.995 131.530 116.760 131.670 ;
        RECT 115.995 131.485 116.285 131.530 ;
        RECT 116.440 131.470 116.760 131.530 ;
        RECT 117.375 131.485 117.665 131.715 ;
        RECT 118.295 131.670 118.585 131.715 ;
        RECT 118.295 131.530 121.730 131.670 ;
        RECT 118.295 131.485 118.585 131.530 ;
        RECT 117.450 131.330 117.590 131.485 ;
        RECT 121.590 131.330 121.730 131.530 ;
        RECT 121.975 131.485 122.265 131.715 ;
        RECT 124.260 131.470 124.580 131.730 ;
        RECT 125.195 131.670 125.485 131.715 ;
        RECT 125.640 131.670 125.960 131.730 ;
        RECT 125.195 131.530 125.960 131.670 ;
        RECT 125.195 131.485 125.485 131.530 ;
        RECT 125.640 131.470 125.960 131.530 ;
        RECT 127.480 131.470 127.800 131.730 ;
        RECT 128.415 131.485 128.705 131.715 ;
        RECT 128.875 131.485 129.165 131.715 ;
        RECT 130.255 131.670 130.545 131.715 ;
        RECT 130.790 131.670 130.930 132.210 ;
        RECT 131.635 132.165 131.925 132.210 ;
        RECT 138.075 132.350 138.365 132.395 ;
        RECT 139.915 132.350 140.205 132.395 ;
        RECT 138.075 132.210 140.205 132.350 ;
        RECT 138.075 132.165 138.365 132.210 ;
        RECT 139.915 132.165 140.205 132.210 ;
        RECT 132.080 132.010 132.400 132.070 ;
        RECT 140.450 132.055 140.590 132.550 ;
        RECT 132.080 131.870 139.210 132.010 ;
        RECT 132.080 131.810 132.400 131.870 ;
        RECT 132.540 131.715 132.860 131.730 ;
        RECT 133.090 131.715 133.230 131.870 ;
        RECT 132.530 131.670 132.860 131.715 ;
        RECT 130.255 131.530 130.930 131.670 ;
        RECT 132.170 131.530 132.860 131.670 ;
        RECT 130.255 131.485 130.545 131.530 ;
        RECT 124.350 131.330 124.490 131.470 ;
        RECT 117.450 131.190 119.430 131.330 ;
        RECT 121.590 131.190 124.490 131.330 ;
        RECT 117.820 130.990 118.140 131.050 ;
        RECT 118.740 130.990 119.060 131.050 ;
        RECT 119.290 131.035 119.430 131.190 ;
        RECT 127.940 131.130 128.260 131.390 ;
        RECT 115.610 130.850 119.060 130.990 ;
        RECT 109.080 130.790 109.400 130.850 ;
        RECT 111.380 130.790 111.700 130.850 ;
        RECT 115.060 130.790 115.380 130.850 ;
        RECT 117.820 130.790 118.140 130.850 ;
        RECT 118.740 130.790 119.060 130.850 ;
        RECT 119.215 130.805 119.505 131.035 ;
        RECT 123.800 130.790 124.120 131.050 ;
        RECT 127.035 130.990 127.325 131.035 ;
        RECT 128.490 130.990 128.630 131.485 ;
        RECT 128.950 131.330 129.090 131.485 ;
        RECT 132.170 131.330 132.310 131.530 ;
        RECT 132.530 131.485 132.860 131.530 ;
        RECT 133.015 131.485 133.305 131.715 ;
        RECT 134.380 131.670 134.700 131.730 ;
        RECT 134.185 131.530 134.700 131.670 ;
        RECT 132.540 131.470 132.860 131.485 ;
        RECT 134.380 131.470 134.700 131.530 ;
        RECT 134.840 131.470 135.160 131.730 ;
        RECT 135.300 131.470 135.620 131.730 ;
        RECT 135.760 131.470 136.080 131.730 ;
        RECT 136.220 131.670 136.540 131.730 ;
        RECT 136.695 131.670 136.985 131.715 ;
        RECT 136.220 131.530 136.985 131.670 ;
        RECT 136.220 131.470 136.540 131.530 ;
        RECT 136.695 131.485 136.985 131.530 ;
        RECT 137.155 131.485 137.445 131.715 ;
        RECT 128.950 131.190 132.310 131.330 ;
        RECT 133.460 131.130 133.780 131.390 ;
        RECT 137.230 131.330 137.370 131.485 ;
        RECT 134.470 131.190 137.370 131.330 ;
        RECT 137.600 131.330 137.920 131.390 ;
        RECT 138.535 131.330 138.825 131.375 ;
        RECT 137.600 131.190 138.825 131.330 ;
        RECT 139.070 131.330 139.210 131.870 ;
        RECT 140.375 131.825 140.665 132.055 ;
        RECT 139.455 131.670 139.745 131.715 ;
        RECT 139.900 131.670 140.220 131.730 ;
        RECT 139.455 131.530 140.220 131.670 ;
        RECT 139.455 131.485 139.745 131.530 ;
        RECT 139.900 131.470 140.220 131.530 ;
        RECT 140.360 131.330 140.680 131.390 ;
        RECT 139.070 131.190 140.680 131.330 ;
        RECT 133.550 130.990 133.690 131.130 ;
        RECT 134.470 131.050 134.610 131.190 ;
        RECT 137.600 131.130 137.920 131.190 ;
        RECT 138.535 131.145 138.825 131.190 ;
        RECT 140.360 131.130 140.680 131.190 ;
        RECT 140.820 131.130 141.140 131.390 ;
        RECT 127.035 130.850 133.690 130.990 ;
        RECT 127.035 130.805 127.325 130.850 ;
        RECT 134.380 130.790 134.700 131.050 ;
        RECT 2.750 130.170 159.030 130.650 ;
        RECT 10.180 129.970 10.500 130.030 ;
        RECT 22.600 129.970 22.920 130.030 ;
        RECT 23.980 129.970 24.300 130.030 ;
        RECT 34.100 129.970 34.420 130.030 ;
        RECT 46.060 129.970 46.380 130.030 ;
        RECT 10.180 129.830 31.570 129.970 ;
        RECT 10.180 129.770 10.500 129.830 ;
        RECT 22.600 129.770 22.920 129.830 ;
        RECT 23.980 129.770 24.300 129.830 ;
        RECT 8.340 129.090 8.660 129.350 ;
        RECT 10.270 129.335 10.410 129.770 ;
        RECT 13.855 129.630 14.505 129.675 ;
        RECT 17.455 129.630 17.745 129.675 ;
        RECT 20.300 129.630 20.620 129.690 ;
        RECT 13.855 129.490 20.620 129.630 ;
        RECT 13.855 129.445 14.505 129.490 ;
        RECT 17.155 129.445 17.745 129.490 ;
        RECT 10.195 129.105 10.485 129.335 ;
        RECT 10.660 129.290 10.950 129.335 ;
        RECT 12.495 129.290 12.785 129.335 ;
        RECT 16.075 129.290 16.365 129.335 ;
        RECT 10.660 129.150 16.365 129.290 ;
        RECT 10.660 129.105 10.950 129.150 ;
        RECT 12.495 129.105 12.785 129.150 ;
        RECT 16.075 129.105 16.365 129.150 ;
        RECT 17.155 129.130 17.445 129.445 ;
        RECT 20.300 129.430 20.620 129.490 ;
        RECT 20.775 129.630 21.065 129.675 ;
        RECT 21.220 129.630 21.540 129.690 ;
        RECT 20.775 129.490 21.540 129.630 ;
        RECT 20.775 129.445 21.065 129.490 ;
        RECT 21.220 129.430 21.540 129.490 ;
        RECT 23.055 129.630 23.705 129.675 ;
        RECT 26.655 129.630 26.945 129.675 ;
        RECT 29.500 129.630 29.820 129.690 ;
        RECT 23.055 129.490 29.820 129.630 ;
        RECT 23.055 129.445 23.705 129.490 ;
        RECT 26.355 129.445 26.945 129.490 ;
        RECT 19.380 129.090 19.700 129.350 ;
        RECT 19.860 129.290 20.150 129.335 ;
        RECT 21.695 129.290 21.985 129.335 ;
        RECT 25.275 129.290 25.565 129.335 ;
        RECT 19.860 129.150 25.565 129.290 ;
        RECT 19.860 129.105 20.150 129.150 ;
        RECT 21.695 129.105 21.985 129.150 ;
        RECT 25.275 129.105 25.565 129.150 ;
        RECT 26.355 129.130 26.645 129.445 ;
        RECT 29.500 129.430 29.820 129.490 ;
        RECT 30.880 129.430 31.200 129.690 ;
        RECT 29.975 129.290 30.265 129.335 ;
        RECT 30.970 129.290 31.110 129.430 ;
        RECT 29.975 129.150 31.110 129.290 ;
        RECT 29.975 129.105 30.265 129.150 ;
        RECT 11.560 128.750 11.880 129.010 ;
        RECT 18.920 128.750 19.240 129.010 ;
        RECT 28.120 128.750 28.440 129.010 ;
        RECT 31.430 128.995 31.570 129.830 ;
        RECT 32.810 129.830 34.420 129.970 ;
        RECT 32.810 129.675 32.950 129.830 ;
        RECT 34.100 129.770 34.420 129.830 ;
        RECT 42.470 129.830 46.380 129.970 ;
        RECT 42.470 129.690 42.610 129.830 ;
        RECT 46.060 129.770 46.380 129.830 ;
        RECT 46.520 129.970 46.840 130.030 ;
        RECT 49.755 129.970 50.045 130.015 ;
        RECT 46.520 129.830 50.045 129.970 ;
        RECT 46.520 129.770 46.840 129.830 ;
        RECT 49.755 129.785 50.045 129.830 ;
        RECT 56.195 129.785 56.485 130.015 ;
        RECT 57.100 129.970 57.420 130.030 ;
        RECT 59.860 129.970 60.180 130.030 ;
        RECT 65.395 129.970 65.685 130.015 ;
        RECT 74.120 129.970 74.440 130.030 ;
        RECT 57.100 129.830 74.440 129.970 ;
        RECT 35.020 129.675 35.340 129.690 ;
        RECT 32.735 129.445 33.025 129.675 ;
        RECT 35.015 129.630 35.665 129.675 ;
        RECT 38.615 129.630 38.905 129.675 ;
        RECT 35.015 129.490 38.905 129.630 ;
        RECT 35.015 129.445 35.665 129.490 ;
        RECT 38.315 129.445 38.905 129.490 ;
        RECT 35.020 129.430 35.340 129.445 ;
        RECT 31.820 129.290 32.110 129.335 ;
        RECT 33.655 129.290 33.945 129.335 ;
        RECT 37.235 129.290 37.525 129.335 ;
        RECT 31.820 129.150 37.525 129.290 ;
        RECT 31.820 129.105 32.110 129.150 ;
        RECT 33.655 129.105 33.945 129.150 ;
        RECT 37.235 129.105 37.525 129.150 ;
        RECT 38.315 129.130 38.605 129.445 ;
        RECT 41.920 129.430 42.240 129.690 ;
        RECT 42.380 129.430 42.700 129.690 ;
        RECT 44.215 129.630 44.865 129.675 ;
        RECT 45.600 129.630 45.920 129.690 ;
        RECT 47.815 129.630 48.105 129.675 ;
        RECT 44.215 129.490 48.105 129.630 ;
        RECT 56.270 129.630 56.410 129.785 ;
        RECT 57.100 129.770 57.420 129.830 ;
        RECT 59.860 129.770 60.180 129.830 ;
        RECT 65.395 129.785 65.685 129.830 ;
        RECT 74.120 129.770 74.440 129.830 ;
        RECT 74.595 129.970 74.885 130.015 ;
        RECT 75.960 129.970 76.280 130.030 ;
        RECT 74.595 129.830 76.280 129.970 ;
        RECT 74.595 129.785 74.885 129.830 ;
        RECT 75.960 129.770 76.280 129.830 ;
        RECT 76.420 129.970 76.740 130.030 ;
        RECT 81.035 129.970 81.325 130.015 ;
        RECT 76.420 129.830 81.325 129.970 ;
        RECT 76.420 129.770 76.740 129.830 ;
        RECT 81.035 129.785 81.325 129.830 ;
        RECT 89.760 129.770 90.080 130.030 ;
        RECT 90.680 129.770 91.000 130.030 ;
        RECT 95.280 129.970 95.600 130.030 ;
        RECT 101.260 129.970 101.580 130.030 ;
        RECT 95.280 129.830 101.580 129.970 ;
        RECT 95.280 129.770 95.600 129.830 ;
        RECT 101.260 129.770 101.580 129.830 ;
        RECT 101.720 129.970 102.040 130.030 ;
        RECT 104.495 129.970 104.785 130.015 ;
        RECT 101.720 129.830 104.785 129.970 ;
        RECT 101.720 129.770 102.040 129.830 ;
        RECT 104.495 129.785 104.785 129.830 ;
        RECT 104.940 129.770 105.260 130.030 ;
        RECT 107.240 129.770 107.560 130.030 ;
        RECT 108.620 129.970 108.940 130.030 ;
        RECT 108.250 129.830 108.940 129.970 ;
        RECT 58.035 129.630 58.325 129.675 ;
        RECT 56.270 129.490 58.325 129.630 ;
        RECT 44.215 129.445 44.865 129.490 ;
        RECT 45.600 129.430 45.920 129.490 ;
        RECT 47.515 129.445 48.105 129.490 ;
        RECT 58.035 129.445 58.325 129.490 ;
        RECT 60.315 129.630 60.965 129.675 ;
        RECT 63.080 129.630 63.400 129.690 ;
        RECT 63.915 129.630 64.205 129.675 ;
        RECT 60.315 129.490 64.205 129.630 ;
        RECT 60.315 129.445 60.965 129.490 ;
        RECT 41.020 129.290 41.310 129.335 ;
        RECT 42.855 129.290 43.145 129.335 ;
        RECT 46.435 129.290 46.725 129.335 ;
        RECT 41.020 129.150 46.725 129.290 ;
        RECT 41.020 129.105 41.310 129.150 ;
        RECT 42.855 129.105 43.145 129.150 ;
        RECT 46.435 129.105 46.725 129.150 ;
        RECT 47.515 129.130 47.805 129.445 ;
        RECT 63.080 129.430 63.400 129.490 ;
        RECT 63.615 129.445 64.205 129.490 ;
        RECT 52.515 129.290 52.805 129.335 ;
        RECT 48.220 129.150 52.805 129.290 ;
        RECT 31.355 128.950 31.645 128.995 ;
        RECT 40.080 128.950 40.400 129.010 ;
        RECT 40.555 128.950 40.845 128.995 ;
        RECT 44.220 128.950 44.540 129.010 ;
        RECT 31.355 128.810 44.540 128.950 ;
        RECT 31.355 128.765 31.645 128.810 ;
        RECT 40.080 128.750 40.400 128.810 ;
        RECT 40.555 128.765 40.845 128.810 ;
        RECT 44.220 128.750 44.540 128.810 ;
        RECT 46.980 128.950 47.300 129.010 ;
        RECT 48.220 128.950 48.360 129.150 ;
        RECT 52.515 129.105 52.805 129.150 ;
        RECT 55.275 129.290 55.565 129.335 ;
        RECT 55.720 129.290 56.040 129.350 ;
        RECT 55.275 129.150 56.040 129.290 ;
        RECT 55.275 129.105 55.565 129.150 ;
        RECT 55.720 129.090 56.040 129.150 ;
        RECT 56.180 129.290 56.500 129.350 ;
        RECT 56.655 129.290 56.945 129.335 ;
        RECT 56.180 129.150 56.945 129.290 ;
        RECT 56.180 129.090 56.500 129.150 ;
        RECT 56.655 129.105 56.945 129.150 ;
        RECT 57.120 129.290 57.410 129.335 ;
        RECT 58.955 129.290 59.245 129.335 ;
        RECT 62.535 129.290 62.825 129.335 ;
        RECT 57.120 129.150 62.825 129.290 ;
        RECT 57.120 129.105 57.410 129.150 ;
        RECT 58.955 129.105 59.245 129.150 ;
        RECT 62.535 129.105 62.825 129.150 ;
        RECT 63.615 129.130 63.905 129.445 ;
        RECT 69.060 129.430 69.380 129.690 ;
        RECT 69.980 129.630 70.300 129.690 ;
        RECT 76.510 129.630 76.650 129.770 ;
        RECT 105.030 129.630 105.170 129.770 ;
        RECT 107.330 129.630 107.470 129.770 ;
        RECT 108.250 129.675 108.390 129.830 ;
        RECT 108.620 129.770 108.940 129.830 ;
        RECT 109.080 129.770 109.400 130.030 ;
        RECT 110.000 129.970 110.320 130.030 ;
        RECT 115.980 129.970 116.300 130.030 ;
        RECT 119.200 129.970 119.520 130.030 ;
        RECT 110.000 129.830 111.610 129.970 ;
        RECT 110.000 129.770 110.320 129.830 ;
        RECT 69.980 129.490 71.590 129.630 ;
        RECT 69.980 129.430 70.300 129.490 ;
        RECT 71.450 129.335 71.590 129.490 ;
        RECT 76.050 129.490 76.650 129.630 ;
        RECT 87.090 129.490 91.370 129.630 ;
        RECT 71.375 129.105 71.665 129.335 ;
        RECT 72.280 129.090 72.600 129.350 ;
        RECT 46.980 128.810 48.360 128.950 ;
        RECT 49.295 128.950 49.585 128.995 ;
        RECT 49.740 128.950 50.060 129.010 ;
        RECT 49.295 128.810 50.060 128.950 ;
        RECT 46.980 128.750 47.300 128.810 ;
        RECT 49.295 128.765 49.585 128.810 ;
        RECT 49.740 128.750 50.060 128.810 ;
        RECT 52.040 128.750 52.360 129.010 ;
        RECT 58.020 128.950 58.340 129.010 ;
        RECT 57.190 128.810 58.340 128.950 ;
        RECT 6.960 128.610 7.280 128.670 ;
        RECT 7.435 128.610 7.725 128.655 ;
        RECT 6.960 128.470 7.725 128.610 ;
        RECT 6.960 128.410 7.280 128.470 ;
        RECT 7.435 128.425 7.725 128.470 ;
        RECT 11.065 128.610 11.355 128.655 ;
        RECT 12.955 128.610 13.245 128.655 ;
        RECT 16.075 128.610 16.365 128.655 ;
        RECT 11.065 128.470 16.365 128.610 ;
        RECT 11.065 128.425 11.355 128.470 ;
        RECT 12.955 128.425 13.245 128.470 ;
        RECT 16.075 128.425 16.365 128.470 ;
        RECT 20.265 128.610 20.555 128.655 ;
        RECT 22.155 128.610 22.445 128.655 ;
        RECT 25.275 128.610 25.565 128.655 ;
        RECT 20.265 128.470 25.565 128.610 ;
        RECT 20.265 128.425 20.555 128.470 ;
        RECT 22.155 128.425 22.445 128.470 ;
        RECT 25.275 128.425 25.565 128.470 ;
        RECT 32.225 128.610 32.515 128.655 ;
        RECT 34.115 128.610 34.405 128.655 ;
        RECT 37.235 128.610 37.525 128.655 ;
        RECT 32.225 128.470 37.525 128.610 ;
        RECT 32.225 128.425 32.515 128.470 ;
        RECT 34.115 128.425 34.405 128.470 ;
        RECT 37.235 128.425 37.525 128.470 ;
        RECT 41.425 128.610 41.715 128.655 ;
        RECT 43.315 128.610 43.605 128.655 ;
        RECT 46.435 128.610 46.725 128.655 ;
        RECT 41.425 128.470 46.725 128.610 ;
        RECT 52.130 128.610 52.270 128.750 ;
        RECT 57.190 128.610 57.330 128.810 ;
        RECT 58.020 128.750 58.340 128.810 ;
        RECT 52.130 128.470 57.330 128.610 ;
        RECT 57.525 128.610 57.815 128.655 ;
        RECT 59.415 128.610 59.705 128.655 ;
        RECT 62.535 128.610 62.825 128.655 ;
        RECT 57.525 128.470 62.825 128.610 ;
        RECT 72.370 128.610 72.510 129.090 ;
        RECT 72.740 128.750 73.060 129.010 ;
        RECT 76.050 128.995 76.190 129.490 ;
        RECT 87.090 129.350 87.230 129.490 ;
        RECT 76.435 129.290 76.725 129.335 ;
        RECT 76.880 129.290 77.200 129.350 ;
        RECT 76.435 129.150 77.200 129.290 ;
        RECT 76.435 129.105 76.725 129.150 ;
        RECT 76.880 129.090 77.200 129.150 ;
        RECT 82.875 129.290 83.165 129.335 ;
        RECT 86.555 129.290 86.845 129.335 ;
        RECT 87.000 129.290 87.320 129.350 ;
        RECT 82.875 129.150 85.850 129.290 ;
        RECT 82.875 129.105 83.165 129.150 ;
        RECT 85.710 129.010 85.850 129.150 ;
        RECT 86.555 129.150 87.320 129.290 ;
        RECT 86.555 129.105 86.845 129.150 ;
        RECT 87.000 129.090 87.320 129.150 ;
        RECT 87.475 129.290 87.765 129.335 ;
        RECT 87.935 129.290 88.225 129.335 ;
        RECT 87.475 129.150 88.225 129.290 ;
        RECT 87.475 129.105 87.765 129.150 ;
        RECT 87.935 129.105 88.225 129.150 ;
        RECT 88.855 129.290 89.145 129.335 ;
        RECT 89.300 129.290 89.620 129.350 ;
        RECT 91.230 129.335 91.370 129.490 ;
        RECT 93.530 129.490 99.190 129.630 ;
        RECT 93.530 129.335 93.670 129.490 ;
        RECT 88.855 129.150 89.620 129.290 ;
        RECT 88.855 129.105 89.145 129.150 ;
        RECT 89.300 129.090 89.620 129.150 ;
        RECT 90.235 129.105 90.525 129.335 ;
        RECT 91.155 129.105 91.445 129.335 ;
        RECT 92.535 129.105 92.825 129.335 ;
        RECT 93.455 129.105 93.745 129.335 ;
        RECT 95.280 129.290 95.600 129.350 ;
        RECT 99.050 129.335 99.190 129.490 ;
        RECT 104.110 129.490 105.170 129.630 ;
        RECT 106.410 129.490 107.470 129.630 ;
        RECT 93.990 129.150 95.600 129.290 ;
        RECT 75.975 128.765 76.265 128.995 ;
        RECT 83.335 128.765 83.625 128.995 ;
        RECT 85.620 128.950 85.940 129.010 ;
        RECT 90.310 128.950 90.450 129.105 ;
        RECT 85.620 128.810 90.450 128.950 ;
        RECT 92.610 128.950 92.750 129.105 ;
        RECT 93.990 128.950 94.130 129.150 ;
        RECT 95.280 129.090 95.600 129.150 ;
        RECT 98.975 129.290 99.265 129.335 ;
        RECT 100.800 129.290 101.120 129.350 ;
        RECT 98.975 129.150 101.120 129.290 ;
        RECT 98.975 129.105 99.265 129.150 ;
        RECT 100.800 129.090 101.120 129.150 ;
        RECT 101.260 129.290 101.580 129.350 ;
        RECT 104.110 129.335 104.250 129.490 ;
        RECT 104.035 129.290 104.325 129.335 ;
        RECT 101.260 129.150 104.325 129.290 ;
        RECT 101.260 129.090 101.580 129.150 ;
        RECT 104.035 129.105 104.325 129.150 ;
        RECT 104.940 129.090 105.260 129.350 ;
        RECT 106.410 129.335 106.550 129.490 ;
        RECT 108.175 129.445 108.465 129.675 ;
        RECT 109.170 129.630 109.310 129.770 ;
        RECT 109.170 129.490 111.150 129.630 ;
        RECT 107.240 129.335 107.560 129.350 ;
        RECT 106.335 129.105 106.625 129.335 ;
        RECT 107.075 129.105 107.560 129.335 ;
        RECT 107.715 129.105 108.005 129.335 ;
        RECT 108.660 129.290 108.950 129.335 ;
        RECT 109.540 129.290 109.860 129.350 ;
        RECT 111.010 129.335 111.150 129.490 ;
        RECT 111.470 129.335 111.610 129.830 ;
        RECT 115.980 129.830 119.520 129.970 ;
        RECT 115.980 129.770 116.300 129.830 ;
        RECT 119.200 129.770 119.520 129.830 ;
        RECT 120.135 129.970 120.425 130.015 ;
        RECT 130.240 129.970 130.560 130.030 ;
        RECT 120.135 129.830 130.560 129.970 ;
        RECT 120.135 129.785 120.425 129.830 ;
        RECT 130.240 129.770 130.560 129.830 ;
        RECT 131.175 129.970 131.465 130.015 ;
        RECT 133.460 129.970 133.780 130.030 ;
        RECT 131.175 129.830 133.780 129.970 ;
        RECT 131.175 129.785 131.465 129.830 ;
        RECT 133.460 129.770 133.780 129.830 ;
        RECT 140.820 129.770 141.140 130.030 ;
        RECT 121.960 129.430 122.280 129.690 ;
        RECT 124.260 129.630 124.580 129.690 ;
        RECT 140.910 129.630 141.050 129.770 ;
        RECT 124.260 129.490 141.050 129.630 ;
        RECT 124.260 129.430 124.580 129.490 ;
        RECT 108.250 129.150 109.860 129.290 ;
        RECT 107.240 129.090 107.560 129.105 ;
        RECT 92.610 128.810 94.130 128.950 ;
        RECT 94.835 128.950 95.125 128.995 ;
        RECT 99.895 128.950 100.185 128.995 ;
        RECT 94.835 128.810 100.185 128.950 ;
        RECT 72.370 128.470 77.570 128.610 ;
        RECT 41.425 128.425 41.715 128.470 ;
        RECT 43.315 128.425 43.605 128.470 ;
        RECT 46.435 128.425 46.725 128.470 ;
        RECT 57.525 128.425 57.815 128.470 ;
        RECT 59.415 128.425 59.705 128.470 ;
        RECT 62.535 128.425 62.825 128.470 ;
        RECT 77.430 128.330 77.570 128.470 ;
        RECT 83.410 128.330 83.550 128.765 ;
        RECT 85.620 128.750 85.940 128.810 ;
        RECT 94.835 128.765 95.125 128.810 ;
        RECT 99.895 128.765 100.185 128.810 ;
        RECT 103.575 128.950 103.865 128.995 ;
        RECT 104.480 128.950 104.800 129.010 ;
        RECT 107.790 128.950 107.930 129.105 ;
        RECT 103.575 128.810 107.930 128.950 ;
        RECT 103.575 128.765 103.865 128.810 ;
        RECT 104.480 128.750 104.800 128.810 ;
        RECT 87.460 128.610 87.780 128.670 ;
        RECT 91.615 128.610 91.905 128.655 ;
        RECT 87.460 128.470 91.905 128.610 ;
        RECT 87.460 128.410 87.780 128.470 ;
        RECT 91.615 128.425 91.905 128.470 ;
        RECT 98.040 128.610 98.360 128.670 ;
        RECT 100.340 128.610 100.660 128.670 ;
        RECT 108.250 128.610 108.390 129.150 ;
        RECT 108.660 129.105 108.950 129.150 ;
        RECT 109.540 129.090 109.860 129.150 ;
        RECT 110.935 129.105 111.225 129.335 ;
        RECT 111.395 129.105 111.685 129.335 ;
        RECT 114.600 129.290 114.920 129.350 ;
        RECT 117.375 129.290 117.665 129.335 ;
        RECT 114.600 129.150 117.665 129.290 ;
        RECT 114.600 129.090 114.920 129.150 ;
        RECT 117.375 129.105 117.665 129.150 ;
        RECT 119.675 129.290 119.965 129.335 ;
        RECT 120.120 129.290 120.440 129.350 ;
        RECT 119.675 129.150 120.440 129.290 ;
        RECT 119.675 129.105 119.965 129.150 ;
        RECT 120.120 129.090 120.440 129.150 ;
        RECT 121.055 129.290 121.345 129.335 ;
        RECT 121.055 129.150 123.110 129.290 ;
        RECT 121.055 129.105 121.345 129.150 ;
        RECT 109.080 128.950 109.400 129.010 ;
        RECT 109.080 128.810 109.770 128.950 ;
        RECT 109.080 128.750 109.400 128.810 ;
        RECT 109.630 128.655 109.770 128.810 ;
        RECT 116.440 128.750 116.760 129.010 ;
        RECT 116.915 128.765 117.205 128.995 ;
        RECT 117.835 128.765 118.125 128.995 ;
        RECT 118.280 128.950 118.600 129.010 ;
        RECT 121.515 128.950 121.805 128.995 ;
        RECT 118.280 128.810 121.805 128.950 ;
        RECT 122.970 128.950 123.110 129.150 ;
        RECT 123.340 129.090 123.660 129.350 ;
        RECT 123.815 129.290 124.105 129.335 ;
        RECT 125.640 129.290 125.960 129.350 ;
        RECT 123.815 129.150 125.960 129.290 ;
        RECT 123.815 129.105 124.105 129.150 ;
        RECT 125.640 129.090 125.960 129.150 ;
        RECT 128.400 129.090 128.720 129.350 ;
        RECT 129.320 129.290 129.640 129.350 ;
        RECT 130.255 129.290 130.545 129.335 ;
        RECT 129.320 129.150 130.545 129.290 ;
        RECT 129.320 129.090 129.640 129.150 ;
        RECT 130.255 129.105 130.545 129.150 ;
        RECT 131.175 129.290 131.465 129.335 ;
        RECT 132.540 129.290 132.860 129.350 ;
        RECT 137.140 129.290 137.460 129.350 ;
        RECT 131.175 129.150 137.460 129.290 ;
        RECT 131.175 129.105 131.465 129.150 ;
        RECT 128.490 128.950 128.630 129.090 ;
        RECT 122.970 128.810 128.630 128.950 ;
        RECT 98.040 128.470 100.660 128.610 ;
        RECT 98.040 128.410 98.360 128.470 ;
        RECT 100.340 128.410 100.660 128.470 ;
        RECT 104.110 128.470 108.390 128.610 ;
        RECT 104.110 128.330 104.250 128.470 ;
        RECT 109.555 128.425 109.845 128.655 ;
        RECT 110.000 128.410 110.320 128.670 ;
        RECT 30.895 128.270 31.185 128.315 ;
        RECT 33.180 128.270 33.500 128.330 ;
        RECT 30.895 128.130 33.500 128.270 ;
        RECT 30.895 128.085 31.185 128.130 ;
        RECT 33.180 128.070 33.500 128.130 ;
        RECT 40.095 128.270 40.385 128.315 ;
        RECT 43.760 128.270 44.080 128.330 ;
        RECT 40.095 128.130 44.080 128.270 ;
        RECT 40.095 128.085 40.385 128.130 ;
        RECT 43.760 128.070 44.080 128.130 ;
        RECT 45.140 128.270 45.460 128.330 ;
        RECT 57.100 128.270 57.420 128.330 ;
        RECT 45.140 128.130 57.420 128.270 ;
        RECT 45.140 128.070 45.460 128.130 ;
        RECT 57.100 128.070 57.420 128.130 ;
        RECT 77.340 128.070 77.660 128.330 ;
        RECT 83.320 128.070 83.640 128.330 ;
        RECT 84.240 128.270 84.560 128.330 ;
        RECT 102.640 128.270 102.960 128.330 ;
        RECT 84.240 128.130 102.960 128.270 ;
        RECT 84.240 128.070 84.560 128.130 ;
        RECT 102.640 128.070 102.960 128.130 ;
        RECT 104.020 128.070 104.340 128.330 ;
        RECT 115.520 128.070 115.840 128.330 ;
        RECT 116.990 128.270 117.130 128.765 ;
        RECT 117.910 128.610 118.050 128.765 ;
        RECT 118.280 128.750 118.600 128.810 ;
        RECT 121.515 128.765 121.805 128.810 ;
        RECT 128.400 128.610 128.720 128.670 ;
        RECT 117.910 128.470 128.720 128.610 ;
        RECT 130.330 128.610 130.470 129.105 ;
        RECT 132.540 129.090 132.860 129.150 ;
        RECT 137.140 129.090 137.460 129.150 ;
        RECT 138.995 129.290 139.285 129.335 ;
        RECT 138.995 129.150 140.130 129.290 ;
        RECT 138.995 129.105 139.285 129.150 ;
        RECT 133.475 128.950 133.765 128.995 ;
        RECT 133.920 128.950 134.240 129.010 ;
        RECT 133.475 128.810 134.240 128.950 ;
        RECT 133.475 128.765 133.765 128.810 ;
        RECT 133.920 128.750 134.240 128.810 ;
        RECT 135.760 128.950 136.080 129.010 ;
        RECT 137.615 128.950 137.905 128.995 ;
        RECT 139.455 128.950 139.745 128.995 ;
        RECT 135.760 128.810 139.745 128.950 ;
        RECT 135.760 128.750 136.080 128.810 ;
        RECT 137.615 128.765 137.905 128.810 ;
        RECT 139.455 128.765 139.745 128.810 ;
        RECT 134.380 128.610 134.700 128.670 ;
        RECT 139.990 128.610 140.130 129.150 ;
        RECT 130.330 128.470 140.130 128.610 ;
        RECT 128.400 128.410 128.720 128.470 ;
        RECT 134.380 128.410 134.700 128.470 ;
        RECT 117.820 128.270 118.140 128.330 ;
        RECT 116.990 128.130 118.140 128.270 ;
        RECT 117.820 128.070 118.140 128.130 ;
        RECT 121.055 128.270 121.345 128.315 ;
        RECT 122.420 128.270 122.740 128.330 ;
        RECT 121.055 128.130 122.740 128.270 ;
        RECT 121.055 128.085 121.345 128.130 ;
        RECT 122.420 128.070 122.740 128.130 ;
        RECT 124.720 128.070 125.040 128.330 ;
        RECT 135.295 128.270 135.585 128.315 ;
        RECT 136.215 128.270 136.505 128.315 ;
        RECT 135.295 128.130 136.505 128.270 ;
        RECT 135.295 128.085 135.585 128.130 ;
        RECT 136.215 128.085 136.505 128.130 ;
        RECT 2.750 127.450 158.230 127.930 ;
        RECT 8.340 127.250 8.660 127.310 ;
        RECT 9.275 127.250 9.565 127.295 ;
        RECT 8.340 127.110 9.565 127.250 ;
        RECT 8.340 127.050 8.660 127.110 ;
        RECT 9.275 127.065 9.565 127.110 ;
        RECT 11.560 127.250 11.880 127.310 ;
        RECT 13.875 127.250 14.165 127.295 ;
        RECT 11.560 127.110 14.165 127.250 ;
        RECT 11.560 127.050 11.880 127.110 ;
        RECT 13.875 127.065 14.165 127.110 ;
        RECT 16.160 127.050 16.480 127.310 ;
        RECT 18.460 127.250 18.780 127.310 ;
        RECT 18.935 127.250 19.225 127.295 ;
        RECT 18.460 127.110 19.225 127.250 ;
        RECT 18.460 127.050 18.780 127.110 ;
        RECT 18.935 127.065 19.225 127.110 ;
        RECT 29.040 127.050 29.360 127.310 ;
        RECT 33.655 127.250 33.945 127.295 ;
        RECT 34.100 127.250 34.420 127.310 ;
        RECT 33.655 127.110 34.420 127.250 ;
        RECT 33.655 127.065 33.945 127.110 ;
        RECT 34.100 127.050 34.420 127.110 ;
        RECT 39.160 127.250 39.480 127.310 ;
        RECT 40.095 127.250 40.385 127.295 ;
        RECT 39.160 127.110 40.385 127.250 ;
        RECT 39.160 127.050 39.480 127.110 ;
        RECT 40.095 127.065 40.385 127.110 ;
        RECT 41.920 127.250 42.240 127.310 ;
        RECT 42.395 127.250 42.685 127.295 ;
        RECT 41.920 127.110 42.685 127.250 ;
        RECT 41.920 127.050 42.240 127.110 ;
        RECT 42.395 127.065 42.685 127.110 ;
        RECT 42.840 127.250 43.160 127.310 ;
        RECT 55.720 127.250 56.040 127.310 ;
        RECT 58.495 127.250 58.785 127.295 ;
        RECT 42.840 127.110 49.970 127.250 ;
        RECT 42.840 127.050 43.160 127.110 ;
        RECT 12.495 126.570 12.785 126.615 ;
        RECT 13.860 126.570 14.180 126.630 ;
        RECT 12.495 126.430 14.180 126.570 ;
        RECT 12.495 126.385 12.785 126.430 ;
        RECT 13.860 126.370 14.180 126.430 ;
        RECT 14.320 126.370 14.640 126.630 ;
        RECT 11.575 126.230 11.865 126.275 ;
        RECT 14.410 126.230 14.550 126.370 ;
        RECT 11.575 126.090 14.550 126.230 ;
        RECT 14.795 126.230 15.085 126.275 ;
        RECT 16.250 126.230 16.390 127.050 ;
        RECT 34.190 126.770 40.310 126.910 ;
        RECT 18.920 126.570 19.240 126.630 ;
        RECT 21.695 126.570 21.985 126.615 ;
        RECT 18.920 126.430 21.985 126.570 ;
        RECT 18.920 126.370 19.240 126.430 ;
        RECT 21.695 126.385 21.985 126.430 ;
        RECT 32.275 126.570 32.565 126.615 ;
        RECT 33.640 126.570 33.960 126.630 ;
        RECT 32.275 126.430 33.960 126.570 ;
        RECT 32.275 126.385 32.565 126.430 ;
        RECT 33.640 126.370 33.960 126.430 ;
        RECT 14.795 126.090 16.390 126.230 ;
        RECT 11.575 126.045 11.865 126.090 ;
        RECT 14.795 126.045 15.085 126.090 ;
        RECT 11.115 125.890 11.405 125.935 ;
        RECT 12.480 125.890 12.800 125.950 ;
        RECT 34.190 125.890 34.330 126.770 ;
        RECT 38.255 126.570 38.545 126.615 ;
        RECT 38.700 126.570 39.020 126.630 ;
        RECT 38.255 126.430 39.020 126.570 ;
        RECT 40.170 126.570 40.310 126.770 ;
        RECT 43.775 126.725 44.065 126.955 ;
        RECT 44.220 126.910 44.540 126.970 ;
        RECT 44.220 126.770 49.510 126.910 ;
        RECT 42.380 126.570 42.700 126.630 ;
        RECT 40.170 126.430 42.700 126.570 ;
        RECT 38.255 126.385 38.545 126.430 ;
        RECT 34.575 126.230 34.865 126.275 ;
        RECT 35.480 126.230 35.800 126.290 ;
        RECT 36.875 126.230 37.165 126.275 ;
        RECT 34.575 126.090 35.250 126.230 ;
        RECT 34.575 126.045 34.865 126.090 ;
        RECT 11.115 125.750 34.330 125.890 ;
        RECT 11.115 125.705 11.405 125.750 ;
        RECT 12.480 125.690 12.800 125.750 ;
        RECT 35.110 125.595 35.250 126.090 ;
        RECT 35.480 126.090 37.165 126.230 ;
        RECT 35.480 126.030 35.800 126.090 ;
        RECT 36.875 126.045 37.165 126.090 ;
        RECT 36.950 125.890 37.090 126.045 ;
        RECT 38.335 125.890 38.475 126.385 ;
        RECT 38.700 126.370 39.020 126.430 ;
        RECT 42.380 126.370 42.700 126.430 ;
        RECT 39.620 126.230 39.940 126.290 ;
        RECT 41.015 126.230 41.305 126.275 ;
        RECT 39.620 126.090 41.305 126.230 ;
        RECT 39.620 126.030 39.940 126.090 ;
        RECT 41.015 126.045 41.305 126.090 ;
        RECT 43.315 126.230 43.605 126.275 ;
        RECT 43.850 126.230 43.990 126.725 ;
        RECT 44.220 126.710 44.540 126.770 ;
        RECT 49.370 126.615 49.510 126.770 ;
        RECT 46.535 126.570 46.825 126.615 ;
        RECT 43.315 126.090 43.990 126.230 ;
        RECT 44.310 126.430 46.825 126.570 ;
        RECT 43.315 126.045 43.605 126.090 ;
        RECT 44.310 125.890 44.450 126.430 ;
        RECT 46.535 126.385 46.825 126.430 ;
        RECT 49.295 126.385 49.585 126.615 ;
        RECT 49.830 126.570 49.970 127.110 ;
        RECT 55.720 127.110 58.785 127.250 ;
        RECT 55.720 127.050 56.040 127.110 ;
        RECT 58.495 127.065 58.785 127.110 ;
        RECT 74.580 127.050 74.900 127.310 ;
        RECT 76.435 127.250 76.725 127.295 ;
        RECT 76.880 127.250 77.200 127.310 ;
        RECT 76.435 127.110 77.200 127.250 ;
        RECT 76.435 127.065 76.725 127.110 ;
        RECT 76.880 127.050 77.200 127.110 ;
        RECT 77.340 127.050 77.660 127.310 ;
        RECT 83.320 127.050 83.640 127.310 ;
        RECT 84.240 127.250 84.560 127.310 ;
        RECT 83.870 127.110 84.560 127.250 ;
        RECT 50.165 126.910 50.455 126.955 ;
        RECT 52.055 126.910 52.345 126.955 ;
        RECT 55.175 126.910 55.465 126.955 ;
        RECT 50.165 126.770 55.465 126.910 ;
        RECT 50.165 126.725 50.455 126.770 ;
        RECT 52.055 126.725 52.345 126.770 ;
        RECT 55.175 126.725 55.465 126.770 ;
        RECT 57.100 126.710 57.420 126.970 ;
        RECT 58.940 126.910 59.260 126.970 ;
        RECT 58.940 126.770 67.910 126.910 ;
        RECT 58.940 126.710 59.260 126.770 ;
        RECT 50.675 126.570 50.965 126.615 ;
        RECT 49.830 126.430 50.965 126.570 ;
        RECT 50.675 126.385 50.965 126.430 ;
        RECT 45.140 126.230 45.460 126.290 ;
        RECT 45.615 126.230 45.905 126.275 ;
        RECT 45.140 126.090 45.905 126.230 ;
        RECT 45.140 126.030 45.460 126.090 ;
        RECT 45.615 126.045 45.905 126.090 ;
        RECT 49.760 126.230 50.050 126.275 ;
        RECT 51.595 126.230 51.885 126.275 ;
        RECT 55.175 126.230 55.465 126.275 ;
        RECT 49.760 126.090 55.465 126.230 ;
        RECT 49.760 126.045 50.050 126.090 ;
        RECT 51.595 126.045 51.885 126.090 ;
        RECT 55.175 126.045 55.465 126.090 ;
        RECT 52.040 125.890 52.360 125.950 ;
        RECT 56.255 125.935 56.545 126.250 ;
        RECT 52.955 125.890 53.605 125.935 ;
        RECT 56.255 125.890 56.845 125.935 ;
        RECT 36.950 125.750 38.010 125.890 ;
        RECT 38.335 125.750 44.450 125.890 ;
        RECT 45.690 125.750 52.360 125.890 ;
        RECT 35.035 125.365 35.325 125.595 ;
        RECT 37.320 125.350 37.640 125.610 ;
        RECT 37.870 125.550 38.010 125.750 ;
        RECT 45.690 125.550 45.830 125.750 ;
        RECT 52.040 125.690 52.360 125.750 ;
        RECT 52.590 125.750 56.845 125.890 ;
        RECT 57.190 125.890 57.330 126.710 ;
        RECT 57.560 126.570 57.880 126.630 ;
        RECT 67.770 126.615 67.910 126.770 ;
        RECT 61.255 126.570 61.545 126.615 ;
        RECT 57.560 126.430 61.545 126.570 ;
        RECT 57.560 126.370 57.880 126.430 ;
        RECT 61.255 126.385 61.545 126.430 ;
        RECT 67.695 126.385 67.985 126.615 ;
        RECT 69.520 126.570 69.840 126.630 ;
        RECT 71.375 126.570 71.665 126.615 ;
        RECT 69.520 126.430 71.665 126.570 ;
        RECT 69.520 126.370 69.840 126.430 ;
        RECT 71.375 126.385 71.665 126.430 ;
        RECT 76.420 126.370 76.740 126.630 ;
        RECT 77.800 126.570 78.120 126.630 ;
        RECT 79.655 126.570 79.945 126.615 ;
        RECT 83.870 126.570 84.010 127.110 ;
        RECT 84.240 127.050 84.560 127.110 ;
        RECT 87.460 127.050 87.780 127.310 ;
        RECT 92.980 127.250 93.300 127.310 ;
        RECT 94.375 127.250 94.665 127.295 ;
        RECT 92.980 127.110 94.665 127.250 ;
        RECT 92.980 127.050 93.300 127.110 ;
        RECT 94.375 127.065 94.665 127.110 ;
        RECT 98.975 127.250 99.265 127.295 ;
        RECT 98.975 127.110 101.950 127.250 ;
        RECT 98.975 127.065 99.265 127.110 ;
        RECT 99.895 126.910 100.185 126.955 ;
        RECT 77.800 126.430 84.010 126.570 ;
        RECT 84.330 126.770 100.185 126.910 ;
        RECT 101.810 126.910 101.950 127.110 ;
        RECT 102.180 127.050 102.500 127.310 ;
        RECT 102.640 127.250 102.960 127.310 ;
        RECT 110.460 127.250 110.780 127.310 ;
        RECT 115.060 127.250 115.380 127.310 ;
        RECT 102.640 127.110 115.380 127.250 ;
        RECT 102.640 127.050 102.960 127.110 ;
        RECT 110.460 127.050 110.780 127.110 ;
        RECT 115.060 127.050 115.380 127.110 ;
        RECT 115.520 127.050 115.840 127.310 ;
        RECT 116.440 127.050 116.760 127.310 ;
        RECT 120.135 127.250 120.425 127.295 ;
        RECT 120.580 127.250 120.900 127.310 ;
        RECT 117.450 127.110 120.900 127.250 ;
        RECT 103.560 126.910 103.880 126.970 ;
        RECT 101.810 126.770 103.880 126.910 ;
        RECT 77.800 126.370 78.120 126.430 ;
        RECT 79.655 126.385 79.945 126.430 ;
        RECT 59.860 126.230 60.180 126.290 ;
        RECT 60.795 126.230 61.085 126.275 ;
        RECT 59.860 126.090 61.085 126.230 ;
        RECT 59.860 126.030 60.180 126.090 ;
        RECT 60.795 126.045 61.085 126.090 ;
        RECT 69.980 126.030 70.300 126.290 ;
        RECT 70.900 126.030 71.220 126.290 ;
        RECT 76.510 126.230 76.650 126.370 ;
        RECT 76.895 126.230 77.185 126.275 ;
        RECT 76.510 126.090 77.185 126.230 ;
        RECT 76.895 126.045 77.185 126.090 ;
        RECT 78.260 126.030 78.580 126.290 ;
        RECT 79.180 126.030 79.500 126.290 ;
        RECT 83.780 126.030 84.100 126.290 ;
        RECT 84.330 126.275 84.470 126.770 ;
        RECT 99.895 126.725 100.185 126.770 ;
        RECT 98.040 126.570 98.360 126.630 ;
        RECT 84.790 126.430 98.360 126.570 ;
        RECT 84.255 126.045 84.545 126.275 ;
        RECT 60.335 125.890 60.625 125.935 ;
        RECT 67.680 125.890 68.000 125.950 ;
        RECT 81.940 125.890 82.260 125.950 ;
        RECT 57.190 125.750 82.260 125.890 ;
        RECT 83.870 125.890 84.010 126.030 ;
        RECT 84.790 125.890 84.930 126.430 ;
        RECT 85.620 126.030 85.940 126.290 ;
        RECT 86.095 126.045 86.385 126.275 ;
        RECT 87.000 126.230 87.320 126.290 ;
        RECT 89.850 126.275 89.990 126.430 ;
        RECT 98.040 126.370 98.360 126.430 ;
        RECT 98.500 126.570 98.820 126.630 ;
        RECT 99.435 126.570 99.725 126.615 ;
        RECT 98.500 126.430 99.725 126.570 ;
        RECT 99.970 126.570 100.110 126.725 ;
        RECT 103.560 126.710 103.880 126.770 ;
        RECT 109.080 126.710 109.400 126.970 ;
        RECT 115.610 126.910 115.750 127.050 ;
        RECT 114.690 126.770 115.750 126.910 ;
        RECT 104.955 126.570 105.245 126.615 ;
        RECT 108.620 126.570 108.940 126.630 ;
        RECT 99.970 126.430 105.245 126.570 ;
        RECT 98.500 126.370 98.820 126.430 ;
        RECT 99.435 126.385 99.725 126.430 ;
        RECT 104.955 126.385 105.245 126.430 ;
        RECT 107.330 126.430 108.940 126.570 ;
        RECT 88.855 126.230 89.145 126.275 ;
        RECT 87.000 126.090 89.145 126.230 ;
        RECT 86.170 125.890 86.310 126.045 ;
        RECT 87.000 126.030 87.320 126.090 ;
        RECT 88.855 126.045 89.145 126.090 ;
        RECT 89.775 126.045 90.065 126.275 ;
        RECT 90.695 126.230 90.985 126.275 ;
        RECT 97.120 126.230 97.410 126.275 ;
        RECT 98.960 126.230 99.280 126.290 ;
        RECT 90.695 126.090 99.280 126.230 ;
        RECT 90.695 126.045 90.985 126.090 ;
        RECT 97.120 126.045 97.410 126.090 ;
        RECT 83.870 125.750 84.930 125.890 ;
        RECT 85.250 125.750 86.310 125.890 ;
        RECT 87.920 125.890 88.240 125.950 ;
        RECT 90.770 125.890 90.910 126.045 ;
        RECT 98.960 126.030 99.280 126.090 ;
        RECT 99.880 126.030 100.200 126.290 ;
        RECT 100.815 126.230 101.105 126.275 ;
        RECT 101.260 126.230 101.580 126.290 ;
        RECT 100.815 126.090 101.580 126.230 ;
        RECT 100.815 126.045 101.105 126.090 ;
        RECT 101.260 126.030 101.580 126.090 ;
        RECT 104.495 126.230 104.785 126.275 ;
        RECT 107.330 126.230 107.470 126.430 ;
        RECT 108.620 126.370 108.940 126.430 ;
        RECT 104.495 126.090 107.470 126.230 ;
        RECT 107.700 126.230 108.020 126.290 ;
        RECT 109.170 126.275 109.310 126.710 ;
        RECT 114.690 126.275 114.830 126.770 ;
        RECT 115.535 126.385 115.825 126.615 ;
        RECT 108.175 126.230 108.465 126.275 ;
        RECT 107.700 126.090 108.465 126.230 ;
        RECT 104.495 126.045 104.785 126.090 ;
        RECT 107.700 126.030 108.020 126.090 ;
        RECT 108.175 126.045 108.465 126.090 ;
        RECT 109.095 126.045 109.385 126.275 ;
        RECT 113.235 126.230 113.525 126.275 ;
        RECT 109.630 126.090 113.525 126.230 ;
        RECT 87.920 125.750 90.910 125.890 ;
        RECT 92.060 125.890 92.380 125.950 ;
        RECT 93.440 125.890 93.760 125.950 ;
        RECT 92.060 125.750 93.760 125.890 ;
        RECT 37.870 125.410 45.830 125.550 ;
        RECT 46.060 125.350 46.380 125.610 ;
        RECT 51.580 125.550 51.900 125.610 ;
        RECT 52.590 125.550 52.730 125.750 ;
        RECT 52.955 125.705 53.605 125.750 ;
        RECT 56.555 125.705 56.845 125.750 ;
        RECT 60.335 125.705 60.625 125.750 ;
        RECT 67.680 125.690 68.000 125.750 ;
        RECT 81.940 125.690 82.260 125.750 ;
        RECT 51.580 125.410 52.730 125.550 ;
        RECT 53.880 125.550 54.200 125.610 ;
        RECT 58.035 125.550 58.325 125.595 ;
        RECT 53.880 125.410 58.325 125.550 ;
        RECT 51.580 125.350 51.900 125.410 ;
        RECT 53.880 125.350 54.200 125.410 ;
        RECT 58.035 125.365 58.325 125.410 ;
        RECT 82.860 125.550 83.180 125.610 ;
        RECT 85.250 125.595 85.390 125.750 ;
        RECT 87.920 125.690 88.240 125.750 ;
        RECT 92.060 125.690 92.380 125.750 ;
        RECT 93.440 125.690 93.760 125.750 ;
        RECT 104.035 125.890 104.325 125.935 ;
        RECT 106.320 125.890 106.640 125.950 ;
        RECT 109.630 125.890 109.770 126.090 ;
        RECT 113.235 126.045 113.525 126.090 ;
        RECT 114.155 126.045 114.445 126.275 ;
        RECT 114.615 126.045 114.905 126.275 ;
        RECT 104.035 125.750 106.640 125.890 ;
        RECT 104.035 125.705 104.325 125.750 ;
        RECT 106.320 125.690 106.640 125.750 ;
        RECT 106.870 125.750 109.770 125.890 ;
        RECT 110.460 125.890 110.780 125.950 ;
        RECT 110.935 125.890 111.225 125.935 ;
        RECT 110.460 125.750 111.225 125.890 ;
        RECT 85.175 125.550 85.465 125.595 ;
        RECT 82.860 125.410 85.465 125.550 ;
        RECT 82.860 125.350 83.180 125.410 ;
        RECT 85.175 125.365 85.465 125.410 ;
        RECT 88.380 125.350 88.700 125.610 ;
        RECT 94.360 125.595 94.680 125.610 ;
        RECT 94.360 125.365 94.745 125.595 ;
        RECT 94.360 125.350 94.680 125.365 ;
        RECT 95.280 125.350 95.600 125.610 ;
        RECT 96.215 125.550 96.505 125.595 ;
        RECT 96.660 125.550 96.980 125.610 ;
        RECT 96.215 125.410 96.980 125.550 ;
        RECT 96.215 125.365 96.505 125.410 ;
        RECT 96.660 125.350 96.980 125.410 ;
        RECT 97.135 125.550 97.425 125.595 ;
        RECT 99.880 125.550 100.200 125.610 ;
        RECT 97.135 125.410 100.200 125.550 ;
        RECT 97.135 125.365 97.425 125.410 ;
        RECT 99.880 125.350 100.200 125.410 ;
        RECT 100.340 125.550 100.660 125.610 ;
        RECT 106.870 125.550 107.010 125.750 ;
        RECT 110.460 125.690 110.780 125.750 ;
        RECT 110.935 125.705 111.225 125.750 ;
        RECT 111.840 125.690 112.160 125.950 ;
        RECT 100.340 125.410 107.010 125.550 ;
        RECT 100.340 125.350 100.660 125.410 ;
        RECT 107.240 125.350 107.560 125.610 ;
        RECT 110.000 125.350 110.320 125.610 ;
        RECT 114.230 125.550 114.370 126.045 ;
        RECT 115.610 125.890 115.750 126.385 ;
        RECT 115.980 126.230 116.300 126.290 ;
        RECT 116.900 126.230 117.220 126.290 ;
        RECT 117.450 126.275 117.590 127.110 ;
        RECT 120.135 127.065 120.425 127.110 ;
        RECT 120.580 127.050 120.900 127.110 ;
        RECT 124.260 127.050 124.580 127.310 ;
        RECT 124.720 127.250 125.040 127.310 ;
        RECT 124.720 127.110 126.330 127.250 ;
        RECT 124.720 127.050 125.040 127.110 ;
        RECT 118.740 126.710 119.060 126.970 ;
        RECT 118.830 126.570 118.970 126.710 ;
        RECT 118.830 126.430 120.350 126.570 ;
        RECT 115.980 126.090 117.220 126.230 ;
        RECT 115.980 126.030 116.300 126.090 ;
        RECT 116.900 126.030 117.220 126.090 ;
        RECT 117.375 126.045 117.665 126.275 ;
        RECT 119.200 126.030 119.520 126.290 ;
        RECT 120.210 126.275 120.350 126.430 ;
        RECT 120.670 126.275 120.810 127.050 ;
        RECT 124.350 126.910 124.490 127.050 ;
        RECT 122.970 126.770 124.490 126.910 ;
        RECT 121.040 126.570 121.360 126.630 ;
        RECT 121.040 126.430 121.730 126.570 ;
        RECT 121.040 126.370 121.360 126.430 ;
        RECT 121.590 126.275 121.730 126.430 ;
        RECT 122.970 126.275 123.110 126.770 ;
        RECT 125.195 126.725 125.485 126.955 ;
        RECT 123.340 126.370 123.660 126.630 ;
        RECT 120.135 126.045 120.425 126.275 ;
        RECT 120.595 126.045 120.885 126.275 ;
        RECT 121.515 126.045 121.805 126.275 ;
        RECT 121.975 126.045 122.265 126.275 ;
        RECT 122.715 126.090 123.110 126.275 ;
        RECT 123.430 126.230 123.570 126.370 ;
        RECT 124.720 126.275 125.040 126.290 ;
        RECT 123.815 126.230 124.105 126.275 ;
        RECT 123.430 126.090 124.105 126.230 ;
        RECT 122.715 126.045 123.005 126.090 ;
        RECT 123.815 126.045 124.105 126.090 ;
        RECT 124.505 126.045 125.040 126.275 ;
        RECT 125.270 126.230 125.410 126.725 ;
        RECT 126.190 126.275 126.330 127.110 ;
        RECT 128.400 127.050 128.720 127.310 ;
        RECT 133.935 127.250 134.225 127.295 ;
        RECT 135.760 127.250 136.080 127.310 ;
        RECT 133.935 127.110 136.080 127.250 ;
        RECT 133.935 127.065 134.225 127.110 ;
        RECT 135.760 127.050 136.080 127.110 ;
        RECT 134.840 126.910 135.160 126.970 ;
        RECT 127.110 126.770 135.160 126.910 ;
        RECT 127.110 126.275 127.250 126.770 ;
        RECT 134.840 126.710 135.160 126.770 ;
        RECT 135.315 126.570 135.605 126.615 ;
        RECT 137.140 126.570 137.460 126.630 ;
        RECT 133.090 126.430 135.070 126.570 ;
        RECT 125.655 126.230 125.945 126.275 ;
        RECT 125.270 126.090 125.945 126.230 ;
        RECT 125.655 126.045 125.945 126.090 ;
        RECT 126.115 126.045 126.405 126.275 ;
        RECT 127.035 126.045 127.325 126.275 ;
        RECT 127.495 126.045 127.785 126.275 ;
        RECT 127.940 126.230 128.260 126.290 ;
        RECT 133.090 126.275 133.230 126.430 ;
        RECT 134.930 126.275 135.070 126.430 ;
        RECT 135.315 126.430 137.460 126.570 ;
        RECT 135.315 126.385 135.605 126.430 ;
        RECT 133.015 126.230 133.305 126.275 ;
        RECT 127.940 126.090 133.305 126.230 ;
        RECT 118.295 125.890 118.585 125.935 ;
        RECT 119.660 125.890 119.980 125.950 ;
        RECT 121.040 125.890 121.360 125.950 ;
        RECT 115.610 125.750 119.980 125.890 ;
        RECT 118.295 125.705 118.585 125.750 ;
        RECT 119.660 125.690 119.980 125.750 ;
        RECT 120.210 125.750 121.360 125.890 ;
        RECT 120.210 125.550 120.350 125.750 ;
        RECT 121.040 125.690 121.360 125.750 ;
        RECT 114.230 125.410 120.350 125.550 ;
        RECT 120.580 125.350 120.900 125.610 ;
        RECT 122.050 125.550 122.190 126.045 ;
        RECT 124.720 126.030 125.040 126.045 ;
        RECT 123.340 125.690 123.660 125.950 ;
        RECT 125.180 125.690 125.500 125.950 ;
        RECT 126.560 125.890 126.880 125.950 ;
        RECT 127.570 125.890 127.710 126.045 ;
        RECT 127.940 126.030 128.260 126.090 ;
        RECT 133.015 126.045 133.305 126.090 ;
        RECT 134.395 126.045 134.685 126.275 ;
        RECT 134.855 126.045 135.145 126.275 ;
        RECT 126.560 125.750 127.710 125.890 ;
        RECT 134.470 125.890 134.610 126.045 ;
        RECT 135.390 125.890 135.530 126.385 ;
        RECT 137.140 126.370 137.460 126.430 ;
        RECT 134.470 125.750 135.530 125.890 ;
        RECT 126.560 125.690 126.880 125.750 ;
        RECT 125.270 125.550 125.410 125.690 ;
        RECT 122.050 125.410 125.410 125.550 ;
        RECT 132.080 125.350 132.400 125.610 ;
        RECT 136.680 125.350 137.000 125.610 ;
        RECT 2.750 124.730 159.030 125.210 ;
        RECT 37.320 124.530 37.640 124.590 ;
        RECT 38.715 124.530 39.005 124.575 ;
        RECT 37.320 124.390 39.005 124.530 ;
        RECT 37.320 124.330 37.640 124.390 ;
        RECT 38.715 124.345 39.005 124.390 ;
        RECT 46.060 124.530 46.380 124.590 ;
        RECT 47.915 124.530 48.205 124.575 ;
        RECT 46.060 124.390 48.205 124.530 ;
        RECT 46.060 124.330 46.380 124.390 ;
        RECT 47.915 124.345 48.205 124.390 ;
        RECT 77.815 124.530 78.105 124.575 ;
        RECT 78.260 124.530 78.580 124.590 ;
        RECT 77.815 124.390 78.580 124.530 ;
        RECT 77.815 124.345 78.105 124.390 ;
        RECT 78.260 124.330 78.580 124.390 ;
        RECT 86.540 124.330 86.860 124.590 ;
        RECT 87.920 124.330 88.240 124.590 ;
        RECT 88.380 124.530 88.700 124.590 ;
        RECT 88.380 124.390 89.070 124.530 ;
        RECT 88.380 124.330 88.700 124.390 ;
        RECT 67.680 123.990 68.000 124.250 ;
        RECT 78.735 124.190 79.025 124.235 ;
        RECT 76.970 124.050 79.025 124.190 ;
        RECT 76.970 123.910 77.110 124.050 ;
        RECT 78.735 124.005 79.025 124.050 ;
        RECT 79.180 123.990 79.500 124.250 ;
        RECT 88.010 124.190 88.150 124.330 ;
        RECT 84.790 124.050 88.150 124.190 ;
        RECT 88.930 124.190 89.070 124.390 ;
        RECT 91.140 124.330 91.460 124.590 ;
        RECT 92.520 124.530 92.840 124.590 ;
        RECT 94.360 124.530 94.680 124.590 ;
        RECT 106.780 124.530 107.100 124.590 ;
        RECT 109.540 124.530 109.860 124.590 ;
        RECT 92.520 124.390 94.680 124.530 ;
        RECT 92.520 124.330 92.840 124.390 ;
        RECT 94.360 124.330 94.680 124.390 ;
        RECT 94.910 124.390 107.100 124.530 ;
        RECT 93.915 124.190 94.205 124.235 ;
        RECT 94.910 124.190 95.050 124.390 ;
        RECT 106.780 124.330 107.100 124.390 ;
        RECT 107.330 124.390 109.860 124.530 ;
        RECT 104.480 124.190 104.800 124.250 ;
        RECT 107.330 124.190 107.470 124.390 ;
        RECT 109.540 124.330 109.860 124.390 ;
        RECT 111.840 124.530 112.160 124.590 ;
        RECT 113.235 124.530 113.525 124.575 ;
        RECT 111.840 124.390 113.525 124.530 ;
        RECT 111.840 124.330 112.160 124.390 ;
        RECT 113.235 124.345 113.525 124.390 ;
        RECT 116.455 124.530 116.745 124.575 ;
        RECT 116.900 124.530 117.220 124.590 ;
        RECT 127.020 124.530 127.340 124.590 ;
        RECT 130.715 124.530 131.005 124.575 ;
        RECT 133.000 124.530 133.320 124.590 ;
        RECT 135.315 124.530 135.605 124.575 ;
        RECT 116.455 124.390 117.220 124.530 ;
        RECT 116.455 124.345 116.745 124.390 ;
        RECT 116.900 124.330 117.220 124.390 ;
        RECT 119.750 124.390 124.950 124.530 ;
        RECT 88.930 124.050 94.205 124.190 ;
        RECT 41.935 123.850 42.225 123.895 ;
        RECT 43.300 123.850 43.620 123.910 ;
        RECT 41.935 123.710 43.620 123.850 ;
        RECT 41.935 123.665 42.225 123.710 ;
        RECT 43.300 123.650 43.620 123.710 ;
        RECT 48.360 123.850 48.680 123.910 ;
        RECT 50.675 123.850 50.965 123.895 ;
        RECT 48.360 123.710 50.965 123.850 ;
        RECT 48.360 123.650 48.680 123.710 ;
        RECT 50.675 123.665 50.965 123.710 ;
        RECT 69.980 123.650 70.300 123.910 ;
        RECT 70.900 123.650 71.220 123.910 ;
        RECT 71.360 123.650 71.680 123.910 ;
        RECT 75.960 123.650 76.280 123.910 ;
        RECT 76.880 123.650 77.200 123.910 ;
        RECT 78.275 123.665 78.565 123.895 ;
        RECT 79.270 123.845 79.410 123.990 ;
        RECT 75.515 123.325 75.805 123.555 ;
        RECT 75.590 123.170 75.730 123.325 ;
        RECT 76.420 123.310 76.740 123.570 ;
        RECT 78.350 123.510 78.490 123.665 ;
        RECT 79.195 123.615 79.485 123.845 ;
        RECT 83.320 123.650 83.640 123.910 ;
        RECT 84.790 123.895 84.930 124.050 ;
        RECT 93.915 124.005 94.205 124.050 ;
        RECT 94.530 124.050 95.050 124.190 ;
        RECT 97.670 124.050 104.800 124.190 ;
        RECT 84.715 123.665 85.005 123.895 ;
        RECT 87.935 123.850 88.225 123.895 ;
        RECT 88.380 123.850 88.700 123.910 ;
        RECT 89.760 123.850 90.080 123.910 ;
        RECT 92.075 123.850 92.365 123.895 ;
        RECT 87.935 123.710 88.700 123.850 ;
        RECT 87.935 123.665 88.225 123.710 ;
        RECT 88.380 123.650 88.700 123.710 ;
        RECT 88.930 123.710 92.365 123.850 ;
        RECT 78.720 123.510 79.040 123.570 ;
        RECT 78.350 123.370 79.040 123.510 ;
        RECT 78.720 123.310 79.040 123.370 ;
        RECT 81.035 123.510 81.325 123.555 ;
        RECT 82.860 123.510 83.180 123.570 ;
        RECT 81.035 123.370 83.180 123.510 ;
        RECT 81.035 123.325 81.325 123.370 ;
        RECT 82.860 123.310 83.180 123.370 ;
        RECT 86.555 123.510 86.845 123.555 ;
        RECT 88.930 123.510 89.070 123.710 ;
        RECT 89.760 123.650 90.080 123.710 ;
        RECT 92.075 123.665 92.365 123.710 ;
        RECT 92.520 123.650 92.840 123.910 ;
        RECT 92.980 123.650 93.300 123.910 ;
        RECT 94.530 123.850 94.670 124.050 ;
        RECT 93.990 123.710 94.670 123.850 ;
        RECT 86.555 123.370 89.070 123.510 ;
        RECT 86.555 123.325 86.845 123.370 ;
        RECT 89.315 123.325 89.605 123.555 ;
        RECT 90.235 123.510 90.525 123.555 ;
        RECT 92.610 123.510 92.750 123.650 ;
        RECT 90.235 123.370 92.750 123.510 ;
        RECT 90.235 123.325 90.525 123.370 ;
        RECT 89.390 123.170 89.530 123.325 ;
        RECT 90.680 123.170 91.000 123.230 ;
        RECT 93.070 123.170 93.210 123.650 ;
        RECT 93.990 123.570 94.130 123.710 ;
        RECT 95.280 123.650 95.600 123.910 ;
        RECT 95.755 123.850 96.045 123.895 ;
        RECT 96.200 123.850 96.520 123.910 ;
        RECT 95.755 123.710 96.520 123.850 ;
        RECT 95.755 123.665 96.045 123.710 ;
        RECT 96.200 123.650 96.520 123.710 ;
        RECT 96.660 123.650 96.980 123.910 ;
        RECT 97.120 123.650 97.440 123.910 ;
        RECT 93.900 123.310 94.220 123.570 ;
        RECT 94.820 123.510 95.140 123.570 ;
        RECT 97.670 123.510 97.810 124.050 ;
        RECT 104.480 123.990 104.800 124.050 ;
        RECT 105.490 124.050 107.470 124.190 ;
        RECT 98.040 123.840 98.360 123.910 ;
        RECT 98.975 123.840 99.265 123.895 ;
        RECT 98.040 123.700 99.265 123.840 ;
        RECT 98.040 123.650 98.360 123.700 ;
        RECT 98.975 123.665 99.265 123.700 ;
        RECT 99.880 123.650 100.200 123.910 ;
        RECT 104.020 123.650 104.340 123.910 ;
        RECT 104.940 123.650 105.260 123.910 ;
        RECT 105.490 123.895 105.630 124.050 ;
        RECT 107.700 123.990 108.020 124.250 ;
        RECT 117.375 124.190 117.665 124.235 ;
        RECT 110.550 124.050 117.665 124.190 ;
        RECT 105.415 123.665 105.705 123.895 ;
        RECT 106.320 123.650 106.640 123.910 ;
        RECT 108.635 123.850 108.925 123.895 ;
        RECT 107.790 123.710 108.925 123.850 ;
        RECT 94.820 123.370 97.810 123.510 ;
        RECT 98.515 123.510 98.805 123.555 ;
        RECT 99.970 123.510 100.110 123.650 ;
        RECT 98.515 123.370 100.110 123.510 ;
        RECT 101.720 123.510 102.040 123.570 ;
        RECT 105.030 123.510 105.170 123.650 ;
        RECT 107.240 123.510 107.560 123.570 ;
        RECT 101.720 123.370 107.560 123.510 ;
        RECT 94.820 123.310 95.140 123.370 ;
        RECT 98.515 123.325 98.805 123.370 ;
        RECT 101.720 123.310 102.040 123.370 ;
        RECT 107.240 123.310 107.560 123.370 ;
        RECT 75.590 123.030 85.390 123.170 ;
        RECT 89.390 123.030 93.210 123.170 ;
        RECT 98.960 123.170 99.280 123.230 ;
        RECT 107.790 123.215 107.930 123.710 ;
        RECT 108.635 123.665 108.925 123.710 ;
        RECT 110.000 123.650 110.320 123.910 ;
        RECT 110.550 123.230 110.690 124.050 ;
        RECT 117.375 124.005 117.665 124.050 ;
        RECT 110.920 123.650 111.240 123.910 ;
        RECT 111.855 123.665 112.145 123.895 ;
        RECT 116.915 123.850 117.205 123.895 ;
        RECT 114.230 123.710 117.205 123.850 ;
        RECT 111.930 123.510 112.070 123.665 ;
        RECT 114.230 123.555 114.370 123.710 ;
        RECT 116.915 123.665 117.205 123.710 ;
        RECT 117.820 123.650 118.140 123.910 ;
        RECT 119.750 123.895 119.890 124.390 ;
        RECT 124.810 124.250 124.950 124.390 ;
        RECT 127.020 124.390 131.005 124.530 ;
        RECT 127.020 124.330 127.340 124.390 ;
        RECT 130.715 124.345 131.005 124.390 ;
        RECT 131.250 124.390 135.605 124.530 ;
        RECT 123.800 124.190 124.120 124.250 ;
        RECT 121.130 124.050 124.120 124.190 ;
        RECT 121.130 123.895 121.270 124.050 ;
        RECT 123.800 123.990 124.120 124.050 ;
        RECT 124.720 124.190 125.040 124.250 ;
        RECT 127.955 124.190 128.245 124.235 ;
        RECT 124.720 124.050 128.245 124.190 ;
        RECT 124.720 123.990 125.040 124.050 ;
        RECT 127.955 124.005 128.245 124.050 ;
        RECT 119.675 123.665 119.965 123.895 ;
        RECT 120.595 123.665 120.885 123.895 ;
        RECT 121.055 123.665 121.345 123.895 ;
        RECT 121.500 123.850 121.820 123.910 ;
        RECT 121.975 123.850 122.265 123.895 ;
        RECT 121.500 123.710 122.265 123.850 ;
        RECT 114.155 123.510 114.445 123.555 ;
        RECT 111.930 123.370 114.445 123.510 ;
        RECT 103.115 123.170 103.405 123.215 ;
        RECT 98.960 123.030 103.405 123.170 ;
        RECT 82.855 122.830 83.145 122.875 ;
        RECT 83.775 122.830 84.065 122.875 ;
        RECT 82.855 122.690 84.065 122.830 ;
        RECT 85.250 122.830 85.390 123.030 ;
        RECT 90.680 122.970 91.000 123.030 ;
        RECT 98.960 122.970 99.280 123.030 ;
        RECT 103.115 122.985 103.405 123.030 ;
        RECT 107.715 122.985 108.005 123.215 ;
        RECT 110.460 123.170 110.780 123.230 ;
        RECT 108.250 123.030 110.780 123.170 ;
        RECT 94.375 122.830 94.665 122.875 ;
        RECT 85.250 122.690 94.665 122.830 ;
        RECT 82.855 122.645 83.145 122.690 ;
        RECT 83.775 122.645 84.065 122.690 ;
        RECT 94.375 122.645 94.665 122.690 ;
        RECT 94.820 122.830 95.140 122.890 ;
        RECT 108.250 122.830 108.390 123.030 ;
        RECT 110.460 122.970 110.780 123.030 ;
        RECT 94.820 122.690 108.390 122.830 ;
        RECT 108.635 122.830 108.925 122.875 ;
        RECT 109.080 122.830 109.400 122.890 ;
        RECT 108.635 122.690 109.400 122.830 ;
        RECT 94.820 122.630 95.140 122.690 ;
        RECT 108.635 122.645 108.925 122.690 ;
        RECT 109.080 122.630 109.400 122.690 ;
        RECT 111.380 122.830 111.700 122.890 ;
        RECT 111.930 122.830 112.070 123.370 ;
        RECT 114.155 123.325 114.445 123.370 ;
        RECT 114.615 123.510 114.905 123.555 ;
        RECT 117.910 123.510 118.050 123.650 ;
        RECT 120.120 123.510 120.440 123.570 ;
        RECT 114.615 123.370 120.440 123.510 ;
        RECT 120.670 123.510 120.810 123.665 ;
        RECT 121.500 123.650 121.820 123.710 ;
        RECT 121.975 123.665 122.265 123.710 ;
        RECT 122.880 123.650 123.200 123.910 ;
        RECT 126.100 123.850 126.420 123.910 ;
        RECT 123.430 123.710 126.420 123.850 ;
        RECT 123.430 123.510 123.570 123.710 ;
        RECT 126.100 123.650 126.420 123.710 ;
        RECT 127.480 123.650 127.800 123.910 ;
        RECT 128.400 123.650 128.720 123.910 ;
        RECT 129.780 123.650 130.100 123.910 ;
        RECT 130.790 123.570 130.930 124.345 ;
        RECT 131.250 123.895 131.390 124.390 ;
        RECT 133.000 124.330 133.320 124.390 ;
        RECT 135.315 124.345 135.605 124.390 ;
        RECT 137.615 124.190 137.905 124.235 ;
        RECT 132.170 124.050 137.905 124.190 ;
        RECT 132.170 123.910 132.310 124.050 ;
        RECT 137.615 124.005 137.905 124.050 ;
        RECT 131.175 123.665 131.465 123.895 ;
        RECT 132.080 123.650 132.400 123.910 ;
        RECT 133.935 123.665 134.225 123.895 ;
        RECT 120.670 123.370 123.570 123.510 ;
        RECT 123.800 123.510 124.120 123.570 ;
        RECT 126.575 123.510 126.865 123.555 ;
        RECT 127.940 123.510 128.260 123.570 ;
        RECT 123.800 123.370 128.260 123.510 ;
        RECT 114.615 123.325 114.905 123.370 ;
        RECT 120.120 123.310 120.440 123.370 ;
        RECT 123.800 123.310 124.120 123.370 ;
        RECT 126.575 123.325 126.865 123.370 ;
        RECT 127.940 123.310 128.260 123.370 ;
        RECT 130.700 123.510 131.020 123.570 ;
        RECT 134.010 123.510 134.150 123.665 ;
        RECT 130.700 123.370 134.150 123.510 ;
        RECT 134.855 123.510 135.145 123.555 ;
        RECT 134.855 123.370 136.450 123.510 ;
        RECT 130.700 123.310 131.020 123.370 ;
        RECT 134.855 123.325 135.145 123.370 ;
        RECT 117.360 123.170 117.680 123.230 ;
        RECT 121.040 123.170 121.360 123.230 ;
        RECT 129.795 123.170 130.085 123.215 ;
        RECT 117.360 123.030 120.810 123.170 ;
        RECT 117.360 122.970 117.680 123.030 ;
        RECT 111.380 122.690 112.070 122.830 ;
        RECT 111.380 122.630 111.700 122.690 ;
        RECT 118.740 122.630 119.060 122.890 ;
        RECT 120.670 122.830 120.810 123.030 ;
        RECT 121.040 123.030 130.085 123.170 ;
        RECT 121.040 122.970 121.360 123.030 ;
        RECT 129.795 122.985 130.085 123.030 ;
        RECT 132.540 122.970 132.860 123.230 ;
        RECT 136.310 123.215 136.450 123.370 ;
        RECT 136.235 123.170 136.525 123.215 ;
        RECT 136.680 123.170 137.000 123.230 ;
        RECT 136.235 123.030 137.000 123.170 ;
        RECT 136.235 122.985 136.525 123.030 ;
        RECT 136.680 122.970 137.000 123.030 ;
        RECT 121.500 122.830 121.820 122.890 ;
        RECT 123.340 122.830 123.660 122.890 ;
        RECT 120.670 122.690 123.660 122.830 ;
        RECT 121.500 122.630 121.820 122.690 ;
        RECT 123.340 122.630 123.660 122.690 ;
        RECT 123.835 122.830 124.125 122.875 ;
        RECT 124.755 122.830 125.045 122.875 ;
        RECT 123.835 122.690 125.045 122.830 ;
        RECT 123.835 122.645 124.125 122.690 ;
        RECT 124.755 122.645 125.045 122.690 ;
        RECT 2.750 122.010 158.230 122.490 ;
        RECT 72.755 121.810 73.045 121.855 ;
        RECT 76.420 121.810 76.740 121.870 ;
        RECT 72.755 121.670 76.740 121.810 ;
        RECT 72.755 121.625 73.045 121.670 ;
        RECT 76.420 121.610 76.740 121.670 ;
        RECT 79.180 121.610 79.500 121.870 ;
        RECT 85.620 121.810 85.940 121.870 ;
        RECT 85.250 121.670 88.150 121.810 ;
        RECT 75.515 121.470 75.805 121.515 ;
        RECT 79.270 121.470 79.410 121.610 ;
        RECT 75.515 121.330 79.410 121.470 ;
        RECT 75.515 121.285 75.805 121.330 ;
        RECT 74.595 120.790 74.885 120.835 ;
        RECT 75.590 120.790 75.730 121.285 ;
        RECT 77.815 121.130 78.105 121.175 ;
        RECT 85.250 121.130 85.390 121.670 ;
        RECT 85.620 121.610 85.940 121.670 ;
        RECT 87.460 121.470 87.780 121.530 ;
        RECT 85.710 121.330 87.780 121.470 ;
        RECT 88.010 121.470 88.150 121.670 ;
        RECT 90.680 121.610 91.000 121.870 ;
        RECT 94.360 121.610 94.680 121.870 ;
        RECT 96.660 121.810 96.980 121.870 ;
        RECT 96.660 121.670 104.250 121.810 ;
        RECT 96.660 121.610 96.980 121.670 ;
        RECT 98.040 121.470 98.360 121.530 ;
        RECT 88.010 121.330 98.360 121.470 ;
        RECT 85.710 121.175 85.850 121.330 ;
        RECT 87.460 121.270 87.780 121.330 ;
        RECT 98.040 121.270 98.360 121.330 ;
        RECT 99.895 121.470 100.185 121.515 ;
        RECT 99.895 121.330 103.790 121.470 ;
        RECT 99.895 121.285 100.185 121.330 ;
        RECT 77.815 120.990 85.390 121.130 ;
        RECT 77.815 120.945 78.105 120.990 ;
        RECT 85.635 120.945 85.925 121.175 ;
        RECT 87.015 120.945 87.305 121.175 ;
        RECT 95.280 121.130 95.600 121.190 ;
        RECT 95.755 121.130 96.045 121.175 ;
        RECT 99.970 121.130 100.110 121.285 ;
        RECT 103.650 121.175 103.790 121.330 ;
        RECT 91.230 120.990 96.045 121.130 ;
        RECT 74.595 120.650 75.730 120.790 ;
        RECT 77.355 120.790 77.645 120.835 ;
        RECT 82.860 120.790 83.180 120.850 ;
        RECT 85.175 120.790 85.465 120.835 ;
        RECT 77.355 120.650 85.465 120.790 ;
        RECT 74.595 120.605 74.885 120.650 ;
        RECT 77.355 120.605 77.645 120.650 ;
        RECT 82.860 120.590 83.180 120.650 ;
        RECT 85.175 120.605 85.465 120.650 ;
        RECT 73.675 120.450 73.965 120.495 ;
        RECT 87.090 120.450 87.230 120.945 ;
        RECT 91.230 120.450 91.370 120.990 ;
        RECT 95.280 120.930 95.600 120.990 ;
        RECT 95.755 120.945 96.045 120.990 ;
        RECT 97.210 120.990 100.110 121.130 ;
        RECT 97.210 120.835 97.350 120.990 ;
        RECT 102.195 120.945 102.485 121.175 ;
        RECT 103.575 120.945 103.865 121.175 ;
        RECT 91.615 120.790 91.905 120.835 ;
        RECT 91.615 120.650 95.050 120.790 ;
        RECT 91.615 120.605 91.905 120.650 ;
        RECT 92.535 120.450 92.825 120.495 ;
        RECT 73.675 120.310 78.950 120.450 ;
        RECT 87.090 120.310 92.825 120.450 ;
        RECT 94.910 120.450 95.050 120.650 ;
        RECT 97.135 120.605 97.425 120.835 ;
        RECT 97.625 120.790 97.915 120.835 ;
        RECT 98.500 120.790 98.820 120.850 ;
        RECT 101.720 120.790 102.040 120.850 ;
        RECT 97.625 120.650 98.270 120.790 ;
        RECT 97.625 120.605 97.915 120.650 ;
        RECT 98.130 120.450 98.270 120.650 ;
        RECT 98.500 120.650 102.040 120.790 ;
        RECT 98.500 120.590 98.820 120.650 ;
        RECT 101.720 120.590 102.040 120.650 ;
        RECT 102.270 120.510 102.410 120.945 ;
        RECT 104.110 120.850 104.250 121.670 ;
        RECT 104.480 121.610 104.800 121.870 ;
        RECT 105.415 121.810 105.705 121.855 ;
        RECT 106.320 121.810 106.640 121.870 ;
        RECT 105.415 121.670 106.640 121.810 ;
        RECT 105.415 121.625 105.705 121.670 ;
        RECT 106.320 121.610 106.640 121.670 ;
        RECT 111.380 121.610 111.700 121.870 ;
        RECT 118.740 121.610 119.060 121.870 ;
        RECT 121.960 121.610 122.280 121.870 ;
        RECT 122.880 121.810 123.200 121.870 ;
        RECT 125.655 121.810 125.945 121.855 ;
        RECT 126.560 121.810 126.880 121.870 ;
        RECT 122.510 121.670 124.950 121.810 ;
        RECT 104.570 121.470 104.710 121.610 ;
        RECT 117.360 121.470 117.680 121.530 ;
        RECT 104.570 121.330 117.680 121.470 ;
        RECT 104.020 120.590 104.340 120.850 ;
        RECT 104.570 120.790 104.710 121.330 ;
        RECT 117.360 121.270 117.680 121.330 ;
        RECT 109.540 121.130 109.860 121.190 ;
        RECT 118.830 121.130 118.970 121.610 ;
        RECT 122.510 121.470 122.650 121.670 ;
        RECT 122.880 121.610 123.200 121.670 ;
        RECT 109.345 120.990 118.970 121.130 ;
        RECT 122.050 121.330 122.650 121.470 ;
        RECT 124.810 121.470 124.950 121.670 ;
        RECT 125.655 121.670 126.880 121.810 ;
        RECT 125.655 121.625 125.945 121.670 ;
        RECT 126.560 121.610 126.880 121.670 ;
        RECT 127.035 121.810 127.325 121.855 ;
        RECT 127.480 121.810 127.800 121.870 ;
        RECT 129.780 121.810 130.100 121.870 ;
        RECT 132.555 121.810 132.845 121.855 ;
        RECT 127.035 121.670 129.090 121.810 ;
        RECT 127.035 121.625 127.325 121.670 ;
        RECT 127.480 121.610 127.800 121.670 ;
        RECT 128.400 121.470 128.720 121.530 ;
        RECT 124.810 121.330 128.720 121.470 ;
        RECT 109.540 120.930 109.860 120.990 ;
        RECT 106.335 120.790 106.625 120.835 ;
        RECT 104.570 120.650 106.625 120.790 ;
        RECT 106.335 120.605 106.625 120.650 ;
        RECT 107.255 120.605 107.545 120.835 ;
        RECT 107.700 120.790 108.020 120.850 ;
        RECT 110.015 120.790 110.305 120.835 ;
        RECT 107.700 120.650 110.305 120.790 ;
        RECT 102.180 120.450 102.500 120.510 ;
        RECT 106.795 120.450 107.085 120.495 ;
        RECT 94.910 120.310 95.970 120.450 ;
        RECT 98.130 120.310 107.085 120.450 ;
        RECT 107.330 120.450 107.470 120.605 ;
        RECT 107.700 120.590 108.020 120.650 ;
        RECT 110.015 120.605 110.305 120.650 ;
        RECT 108.620 120.450 108.940 120.510 ;
        RECT 122.050 120.450 122.190 121.330 ;
        RECT 124.260 120.930 124.580 121.190 ;
        RECT 123.815 120.800 124.105 120.835 ;
        RECT 123.800 120.540 124.120 120.800 ;
        RECT 124.810 120.790 124.950 121.330 ;
        RECT 128.400 121.270 128.720 121.330 ;
        RECT 128.950 121.130 129.090 121.670 ;
        RECT 129.780 121.670 132.845 121.810 ;
        RECT 129.780 121.610 130.100 121.670 ;
        RECT 132.555 121.625 132.845 121.670 ;
        RECT 133.000 121.610 133.320 121.870 ;
        RECT 130.700 121.270 131.020 121.530 ;
        RECT 126.190 120.990 129.090 121.130 ;
        RECT 126.190 120.835 126.330 120.990 ;
        RECT 125.195 120.790 125.485 120.835 ;
        RECT 124.810 120.650 125.485 120.790 ;
        RECT 125.195 120.605 125.485 120.650 ;
        RECT 126.115 120.605 126.405 120.835 ;
        RECT 126.575 120.605 126.865 120.835 ;
        RECT 130.790 120.790 130.930 121.270 ;
        RECT 131.160 121.130 131.480 121.190 ;
        RECT 132.095 121.130 132.385 121.175 ;
        RECT 139.900 121.130 140.220 121.190 ;
        RECT 131.160 120.990 140.220 121.130 ;
        RECT 131.160 120.930 131.480 120.990 ;
        RECT 132.095 120.945 132.385 120.990 ;
        RECT 139.900 120.930 140.220 120.990 ;
        RECT 133.475 120.790 133.765 120.835 ;
        RECT 130.790 120.650 133.765 120.790 ;
        RECT 133.475 120.605 133.765 120.650 ;
        RECT 107.330 120.310 122.190 120.450 ;
        RECT 124.260 120.450 124.580 120.510 ;
        RECT 126.650 120.450 126.790 120.605 ;
        RECT 124.260 120.310 126.790 120.450 ;
        RECT 73.675 120.265 73.965 120.310 ;
        RECT 78.810 120.170 78.950 120.310 ;
        RECT 92.535 120.265 92.825 120.310 ;
        RECT 95.830 120.170 95.970 120.310 ;
        RECT 102.180 120.250 102.500 120.310 ;
        RECT 106.795 120.265 107.085 120.310 ;
        RECT 108.620 120.250 108.940 120.310 ;
        RECT 124.260 120.250 124.580 120.310 ;
        RECT 132.540 120.250 132.860 120.510 ;
        RECT 78.720 120.110 79.040 120.170 ;
        RECT 94.820 120.110 95.140 120.170 ;
        RECT 78.720 119.970 95.140 120.110 ;
        RECT 78.720 119.910 79.040 119.970 ;
        RECT 94.820 119.910 95.140 119.970 ;
        RECT 95.740 120.110 96.060 120.170 ;
        RECT 98.055 120.110 98.345 120.155 ;
        RECT 95.740 119.970 98.345 120.110 ;
        RECT 95.740 119.910 96.060 119.970 ;
        RECT 98.055 119.925 98.345 119.970 ;
        RECT 104.020 120.110 104.340 120.170 ;
        RECT 132.630 120.110 132.770 120.250 ;
        RECT 104.020 119.970 132.770 120.110 ;
        RECT 104.020 119.910 104.340 119.970 ;
        RECT 2.750 119.290 159.030 119.770 ;
        RECT 94.835 119.090 95.125 119.135 ;
        RECT 96.200 119.090 96.520 119.150 ;
        RECT 94.835 118.950 96.520 119.090 ;
        RECT 94.835 118.905 95.125 118.950 ;
        RECT 96.200 118.890 96.520 118.950 ;
        RECT 96.660 118.890 96.980 119.150 ;
        RECT 102.180 119.090 102.500 119.150 ;
        RECT 97.670 118.950 102.500 119.090 ;
        RECT 70.900 118.750 71.220 118.810 ;
        RECT 70.900 118.610 96.430 118.750 ;
        RECT 70.900 118.550 71.220 118.610 ;
        RECT 94.835 118.410 95.125 118.455 ;
        RECT 95.740 118.410 96.060 118.470 ;
        RECT 94.835 118.270 96.060 118.410 ;
        RECT 94.835 118.225 95.125 118.270 ;
        RECT 95.740 118.210 96.060 118.270 ;
        RECT 95.280 117.870 95.600 118.130 ;
        RECT 96.290 118.070 96.430 118.610 ;
        RECT 96.750 118.455 96.890 118.890 ;
        RECT 97.670 118.455 97.810 118.950 ;
        RECT 102.180 118.890 102.500 118.950 ;
        RECT 106.780 119.090 107.100 119.150 ;
        RECT 131.160 119.090 131.480 119.150 ;
        RECT 106.780 118.950 131.480 119.090 ;
        RECT 106.780 118.890 107.100 118.950 ;
        RECT 131.160 118.890 131.480 118.950 ;
        RECT 109.080 118.750 109.400 118.810 ;
        RECT 98.130 118.610 109.400 118.750 ;
        RECT 96.675 118.225 96.965 118.455 ;
        RECT 97.595 118.225 97.885 118.455 ;
        RECT 98.130 118.070 98.270 118.610 ;
        RECT 109.080 118.550 109.400 118.610 ;
        RECT 98.500 118.210 98.820 118.470 ;
        RECT 96.290 117.930 98.270 118.070 ;
        RECT 96.215 117.390 96.505 117.435 ;
        RECT 97.595 117.390 97.885 117.435 ;
        RECT 96.215 117.250 97.885 117.390 ;
        RECT 96.215 117.205 96.505 117.250 ;
        RECT 97.595 117.205 97.885 117.250 ;
        RECT 2.750 116.570 158.230 117.050 ;
        RECT 2.750 113.850 159.030 114.330 ;
        RECT 3.520 98.480 4.520 112.820 ;
        RECT 6.320 97.510 7.320 111.220 ;
        RECT 6.290 96.510 7.350 97.510 ;
        RECT 11.030 94.670 12.030 112.920 ;
        RECT 15.820 92.560 16.820 112.730 ;
        RECT 18.220 91.390 19.220 112.930 ;
        RECT 21.130 91.390 22.130 91.420 ;
        RECT 18.220 90.390 22.130 91.390 ;
        RECT 21.130 90.360 22.130 90.390 ;
        RECT 23.330 88.460 24.330 112.330 ;
        RECT 25.640 87.580 26.640 112.430 ;
        RECT 26.840 87.580 27.840 87.610 ;
        RECT 25.640 86.580 27.840 87.580 ;
        RECT 26.840 86.550 27.840 86.580 ;
        RECT 29.440 85.760 30.440 112.430 ;
        RECT 130.870 99.510 131.870 99.610 ;
        RECT 31.420 98.510 131.870 99.510 ;
        RECT 31.320 96.510 129.030 97.510 ;
        RECT 31.420 94.700 125.930 95.700 ;
        RECT 31.450 93.590 32.450 93.620 ;
        RECT 31.450 92.590 123.040 93.590 ;
        RECT 31.450 92.560 32.450 92.590 ;
        RECT 31.350 91.390 32.350 91.420 ;
        RECT 31.350 90.390 119.870 91.390 ;
        RECT 31.350 90.360 32.350 90.390 ;
        RECT 31.420 88.490 116.870 89.490 ;
        RECT 31.720 86.580 113.870 87.580 ;
        RECT 112.870 85.760 113.870 86.580 ;
        RECT 115.870 85.760 116.870 88.490 ;
        RECT 118.870 85.760 119.870 90.390 ;
        RECT 122.040 85.760 123.040 92.590 ;
        RECT 124.930 85.760 125.930 94.700 ;
        RECT 128.030 85.760 129.030 96.510 ;
        RECT 130.870 85.760 131.870 98.510 ;
        RECT 29.440 84.760 111.070 85.760 ;
        RECT 112.870 84.760 114.070 85.760 ;
        RECT 115.870 84.760 117.070 85.760 ;
        RECT 118.870 84.760 120.070 85.760 ;
        RECT 121.870 84.760 123.070 85.760 ;
        RECT 124.870 84.760 126.070 85.760 ;
        RECT 127.870 84.760 129.070 85.760 ;
        RECT 130.870 84.760 132.070 85.760 ;
        RECT 110.670 80.060 111.070 84.760 ;
        RECT 113.670 80.060 114.070 84.760 ;
        RECT 116.670 80.060 117.070 84.760 ;
        RECT 119.670 80.060 120.070 84.760 ;
        RECT 122.670 80.060 123.070 84.760 ;
        RECT 125.670 80.060 126.070 84.760 ;
        RECT 128.670 80.060 129.070 84.760 ;
        RECT 131.670 80.060 132.070 84.760 ;
        RECT 110.750 79.775 111.000 80.060 ;
        RECT 113.750 79.775 114.000 80.060 ;
        RECT 116.750 79.775 117.000 80.060 ;
        RECT 119.750 79.775 120.000 80.060 ;
        RECT 122.750 79.775 123.000 80.060 ;
        RECT 125.750 79.775 126.000 80.060 ;
        RECT 128.750 79.775 129.000 80.060 ;
        RECT 131.750 79.775 132.000 80.060 ;
        RECT 102.970 77.700 104.030 78.700 ;
        RECT 103.000 13.840 104.000 77.700 ;
        RECT 106.670 55.860 108.970 56.260 ;
        RECT 106.670 53.060 107.070 55.860 ;
        RECT 106.750 52.775 107.000 53.060 ;
        RECT 108.570 38.760 108.970 55.860 ;
        RECT 110.750 38.760 111.000 39.725 ;
        RECT 113.750 38.760 114.000 39.725 ;
        RECT 116.750 38.760 117.000 39.725 ;
        RECT 119.750 38.760 120.000 39.725 ;
        RECT 122.750 38.760 123.000 39.725 ;
        RECT 125.750 38.760 126.000 39.725 ;
        RECT 128.750 38.860 129.000 39.725 ;
        RECT 131.750 38.860 132.000 39.725 ;
        RECT 108.570 38.360 111.070 38.760 ;
        RECT 110.670 32.960 111.070 38.360 ;
        RECT 112.170 38.360 114.070 38.760 ;
        RECT 110.750 32.775 111.000 32.960 ;
        RECT 102.940 12.840 106.360 13.840 ;
        RECT 103.000 11.760 104.000 12.840 ;
        RECT 106.750 12.360 107.000 12.725 ;
        RECT 102.870 11.460 104.000 11.760 ;
        RECT 106.670 11.460 107.070 12.360 ;
        RECT 110.750 11.460 111.000 12.725 ;
        RECT 112.170 11.460 112.570 38.360 ;
        RECT 113.750 37.620 114.000 38.360 ;
        RECT 113.750 34.060 114.000 34.880 ;
        RECT 116.670 34.060 117.070 38.760 ;
        RECT 113.670 33.660 117.070 34.060 ;
        RECT 113.750 32.775 114.000 33.660 ;
        RECT 116.670 32.960 117.070 33.660 ;
        RECT 118.170 38.360 120.070 38.760 ;
        RECT 116.750 32.775 117.000 32.960 ;
        RECT 113.750 11.460 114.000 12.725 ;
        RECT 116.750 11.460 117.000 12.725 ;
        RECT 118.170 11.460 118.570 38.360 ;
        RECT 119.750 37.620 120.000 38.360 ;
        RECT 119.750 34.060 120.000 34.880 ;
        RECT 122.670 34.060 123.070 38.760 ;
        RECT 119.670 33.660 123.070 34.060 ;
        RECT 119.750 32.775 120.000 33.660 ;
        RECT 122.670 32.960 123.070 33.660 ;
        RECT 124.170 38.360 126.070 38.760 ;
        RECT 122.750 32.775 123.000 32.960 ;
        RECT 119.750 11.460 120.000 12.725 ;
        RECT 122.750 11.460 123.000 12.725 ;
        RECT 124.170 11.460 124.570 38.360 ;
        RECT 125.750 37.620 126.000 38.360 ;
        RECT 125.750 34.060 126.000 34.880 ;
        RECT 128.670 34.060 129.070 38.860 ;
        RECT 125.670 33.660 129.070 34.060 ;
        RECT 125.750 32.775 126.000 33.660 ;
        RECT 128.670 33.060 129.070 33.660 ;
        RECT 131.670 35.460 132.070 38.860 ;
        RECT 135.870 37.760 138.500 38.760 ;
        RECT 135.870 35.460 136.270 37.760 ;
        RECT 137.900 35.670 138.500 37.760 ;
        RECT 131.670 35.060 136.270 35.460 ;
        RECT 128.750 32.775 129.000 33.060 ;
        RECT 125.750 11.460 126.000 12.725 ;
        RECT 128.750 12.260 129.000 12.725 ;
        RECT 128.670 11.560 129.070 12.260 ;
        RECT 131.670 11.560 132.070 35.060 ;
        RECT 102.870 11.060 107.070 11.460 ;
        RECT 110.670 11.060 114.070 11.460 ;
        RECT 116.670 11.060 120.070 11.460 ;
        RECT 122.670 11.060 126.070 11.460 ;
        RECT 128.670 11.160 132.070 11.560 ;
        RECT 102.870 10.760 104.000 11.060 ;
        RECT 103.000 10.750 104.000 10.760 ;
        RECT 106.750 10.620 107.000 11.060 ;
        RECT 110.750 10.620 111.000 11.060 ;
        RECT 113.750 10.620 114.000 11.060 ;
        RECT 116.750 10.620 117.000 11.060 ;
        RECT 119.750 10.620 120.000 11.060 ;
        RECT 122.750 10.620 123.000 11.060 ;
        RECT 125.750 10.620 126.000 11.060 ;
        RECT 128.750 10.620 129.000 11.160 ;
      LAYER met2 ;
        RECT 68.620 221.940 68.900 222.055 ;
        RECT 68.230 221.800 68.900 221.940 ;
        RECT 22.620 221.260 22.900 221.375 ;
        RECT 20.330 220.860 20.590 221.180 ;
        RECT 22.620 221.120 23.750 221.260 ;
        RECT 25.390 221.200 25.650 221.520 ;
        RECT 22.620 221.005 22.900 221.120 ;
        RECT 17.570 220.520 17.830 220.840 ;
        RECT 6.530 218.820 6.790 219.140 ;
        RECT 6.590 217.975 6.730 218.820 ;
        RECT 17.630 218.800 17.770 220.520 ;
        RECT 13.430 218.480 13.690 218.800 ;
        RECT 17.570 218.480 17.830 218.800 ;
        RECT 11.130 218.140 11.390 218.460 ;
        RECT 6.520 217.605 6.800 217.975 ;
        RECT 10.660 216.925 10.940 217.295 ;
        RECT 10.670 216.780 10.930 216.925 ;
        RECT 6.070 215.760 6.330 216.080 ;
        RECT 4.690 215.080 4.950 215.400 ;
        RECT 4.750 209.960 4.890 215.080 ;
        RECT 5.610 212.360 5.870 212.680 ;
        RECT 5.670 211.660 5.810 212.360 ;
        RECT 5.610 211.340 5.870 211.660 ;
        RECT 4.690 209.640 4.950 209.960 ;
        RECT 4.750 208.940 4.890 209.640 ;
        RECT 4.690 208.620 4.950 208.940 ;
        RECT 4.750 208.040 4.890 208.620 ;
        RECT 4.750 207.900 5.350 208.040 ;
        RECT 5.210 202.820 5.350 207.900 ;
        RECT 5.610 207.260 5.870 207.580 ;
        RECT 5.670 206.220 5.810 207.260 ;
        RECT 5.610 205.900 5.870 206.220 ;
        RECT 6.130 204.520 6.270 215.760 ;
        RECT 7.900 214.885 8.180 215.255 ;
        RECT 7.970 213.360 8.110 214.885 ;
        RECT 7.910 213.040 8.170 213.360 ;
        RECT 10.210 212.360 10.470 212.680 ;
        RECT 10.270 206.220 10.410 212.360 ;
        RECT 10.730 206.220 10.870 216.780 ;
        RECT 11.190 216.420 11.330 218.140 ;
        RECT 11.130 216.100 11.390 216.420 ;
        RECT 11.190 210.980 11.330 216.100 ;
        RECT 13.490 214.380 13.630 218.480 ;
        RECT 18.030 218.140 18.290 218.460 ;
        RECT 19.410 218.140 19.670 218.460 ;
        RECT 14.810 217.860 15.070 218.120 ;
        RECT 14.410 217.800 15.070 217.860 ;
        RECT 14.410 217.720 15.010 217.800 ;
        RECT 13.430 214.060 13.690 214.380 ;
        RECT 12.510 213.380 12.770 213.700 ;
        RECT 11.130 210.660 11.390 210.980 ;
        RECT 10.210 205.900 10.470 206.220 ;
        RECT 10.670 205.900 10.930 206.220 ;
        RECT 12.570 205.735 12.710 213.380 ;
        RECT 14.410 213.360 14.550 217.720 ;
        RECT 16.190 215.080 16.450 215.400 ;
        RECT 14.350 213.040 14.610 213.360 ;
        RECT 13.890 212.700 14.150 213.020 ;
        RECT 12.970 212.360 13.230 212.680 ;
        RECT 13.030 207.240 13.170 212.360 ;
        RECT 13.430 210.660 13.690 210.980 ;
        RECT 13.490 209.960 13.630 210.660 ;
        RECT 13.430 209.640 13.690 209.960 ;
        RECT 13.430 207.600 13.690 207.920 ;
        RECT 12.970 206.920 13.230 207.240 ;
        RECT 13.030 205.880 13.170 206.920 ;
        RECT 12.500 205.365 12.780 205.735 ;
        RECT 12.970 205.560 13.230 205.880 ;
        RECT 12.570 205.200 12.710 205.365 ;
        RECT 12.510 204.880 12.770 205.200 ;
        RECT 12.970 204.880 13.230 205.200 ;
        RECT 6.070 204.200 6.330 204.520 ;
        RECT 13.030 203.500 13.170 204.880 ;
        RECT 12.970 203.180 13.230 203.500 ;
        RECT 5.150 202.500 5.410 202.820 ;
        RECT 13.490 202.140 13.630 207.600 ;
        RECT 13.950 206.220 14.090 212.700 ;
        RECT 13.890 205.900 14.150 206.220 ;
        RECT 14.410 204.860 14.550 213.040 ;
        RECT 16.250 213.020 16.390 215.080 ;
        RECT 16.640 214.885 16.920 215.255 ;
        RECT 16.190 212.700 16.450 213.020 ;
        RECT 16.710 211.320 16.850 214.885 ;
        RECT 18.090 213.700 18.230 218.140 ;
        RECT 18.950 217.800 19.210 218.120 ;
        RECT 19.010 216.080 19.150 217.800 ;
        RECT 19.470 217.100 19.610 218.140 ;
        RECT 19.410 216.780 19.670 217.100 ;
        RECT 19.860 216.925 20.140 217.295 ;
        RECT 20.390 217.100 20.530 220.860 ;
        RECT 21.415 219.985 22.955 220.355 ;
        RECT 23.090 217.800 23.350 218.120 ;
        RECT 19.870 216.780 20.130 216.925 ;
        RECT 20.330 216.780 20.590 217.100 ;
        RECT 18.950 215.760 19.210 216.080 ;
        RECT 19.930 215.140 20.070 216.780 ;
        RECT 19.930 215.000 20.990 215.140 ;
        RECT 20.850 213.700 20.990 215.000 ;
        RECT 21.415 214.545 22.955 214.915 ;
        RECT 23.150 214.380 23.290 217.800 ;
        RECT 23.610 216.760 23.750 221.120 ;
        RECT 24.930 219.335 25.190 219.480 ;
        RECT 24.920 218.965 25.200 219.335 ;
        RECT 24.990 217.100 25.130 218.965 ;
        RECT 25.450 217.100 25.590 221.200 ;
        RECT 50.690 220.860 50.950 221.180 ;
        RECT 51.610 220.860 51.870 221.180 ;
        RECT 62.640 221.005 62.920 221.375 ;
        RECT 35.040 220.325 35.320 220.695 ;
        RECT 44.240 220.325 44.520 220.695 ;
        RECT 35.110 219.820 35.250 220.325 ;
        RECT 44.310 219.820 44.450 220.325 ;
        RECT 31.830 219.500 32.090 219.820 ;
        RECT 35.050 219.500 35.310 219.820 ;
        RECT 44.250 219.500 44.510 219.820 ;
        RECT 27.690 218.820 27.950 219.140 ;
        RECT 31.370 218.820 31.630 219.140 ;
        RECT 24.930 216.780 25.190 217.100 ;
        RECT 25.390 216.780 25.650 217.100 ;
        RECT 23.550 216.440 23.810 216.760 ;
        RECT 27.230 216.100 27.490 216.420 ;
        RECT 23.090 214.060 23.350 214.380 ;
        RECT 22.630 213.720 22.890 214.040 ;
        RECT 18.030 213.380 18.290 213.700 ;
        RECT 20.790 213.380 21.050 213.700 ;
        RECT 16.650 211.000 16.910 211.320 ;
        RECT 18.090 210.980 18.230 213.380 ;
        RECT 22.690 212.680 22.830 213.720 ;
        RECT 24.930 212.700 25.190 213.020 ;
        RECT 20.790 212.360 21.050 212.680 ;
        RECT 22.630 212.360 22.890 212.680 ;
        RECT 19.870 211.340 20.130 211.660 ;
        RECT 18.030 210.660 18.290 210.980 ;
        RECT 15.270 210.320 15.530 210.640 ;
        RECT 15.330 208.940 15.470 210.320 ;
        RECT 18.090 210.300 18.230 210.660 ;
        RECT 18.030 209.980 18.290 210.300 ;
        RECT 19.930 209.960 20.070 211.340 ;
        RECT 19.870 209.640 20.130 209.960 ;
        RECT 15.270 208.620 15.530 208.940 ;
        RECT 16.190 207.260 16.450 207.580 ;
        RECT 16.250 206.220 16.390 207.260 ;
        RECT 16.650 206.920 16.910 207.240 ;
        RECT 18.030 206.920 18.290 207.240 ;
        RECT 16.190 205.900 16.450 206.220 ;
        RECT 14.350 204.540 14.610 204.860 ;
        RECT 15.270 204.200 15.530 204.520 ;
        RECT 15.330 203.500 15.470 204.200 ;
        RECT 13.890 203.180 14.150 203.500 ;
        RECT 15.270 203.180 15.530 203.500 ;
        RECT 13.430 201.820 13.690 202.140 ;
        RECT 13.490 201.655 13.630 201.820 ;
        RECT 13.420 201.540 13.700 201.655 ;
        RECT 13.030 201.400 13.700 201.540 ;
        RECT 13.030 200.440 13.170 201.400 ;
        RECT 13.420 201.285 13.700 201.400 ;
        RECT 13.950 200.780 14.090 203.180 ;
        RECT 16.250 203.160 16.390 205.900 ;
        RECT 16.190 202.840 16.450 203.160 ;
        RECT 16.710 202.140 16.850 206.920 ;
        RECT 17.110 205.220 17.370 205.540 ;
        RECT 17.570 205.220 17.830 205.540 ;
        RECT 16.650 201.820 16.910 202.140 ;
        RECT 13.890 200.460 14.150 200.780 ;
        RECT 12.970 200.120 13.230 200.440 ;
        RECT 13.430 199.780 13.690 200.100 ;
        RECT 5.610 199.440 5.870 199.760 ;
        RECT 5.670 198.060 5.810 199.440 ;
        RECT 5.610 197.740 5.870 198.060 ;
        RECT 10.670 197.060 10.930 197.380 ;
        RECT 5.610 194.000 5.870 194.320 ;
        RECT 5.670 192.620 5.810 194.000 ;
        RECT 5.610 192.300 5.870 192.620 ;
        RECT 5.150 191.960 5.410 192.280 ;
        RECT 5.210 189.900 5.350 191.960 ;
        RECT 10.730 191.940 10.870 197.060 ;
        RECT 12.510 196.040 12.770 196.360 ;
        RECT 10.670 191.620 10.930 191.940 ;
        RECT 5.150 189.580 5.410 189.900 ;
        RECT 4.690 187.880 4.950 188.200 ;
        RECT 3.770 186.180 4.030 186.500 ;
        RECT 3.830 140.600 3.970 186.180 ;
        RECT 4.750 186.160 4.890 187.880 ;
        RECT 4.690 185.840 4.950 186.160 ;
        RECT 6.070 185.840 6.330 186.160 ;
        RECT 4.750 180.720 4.890 185.840 ;
        RECT 6.130 184.460 6.270 185.840 ;
        RECT 10.730 184.460 10.870 191.620 ;
        RECT 11.130 185.500 11.390 185.820 ;
        RECT 6.070 184.140 6.330 184.460 ;
        RECT 10.670 184.140 10.930 184.460 ;
        RECT 8.830 183.460 9.090 183.780 ;
        RECT 4.690 180.400 4.950 180.720 ;
        RECT 6.070 180.400 6.330 180.720 ;
        RECT 4.750 177.660 4.890 180.400 ;
        RECT 6.130 179.020 6.270 180.400 ;
        RECT 6.070 178.700 6.330 179.020 ;
        RECT 4.690 177.340 4.950 177.660 ;
        RECT 4.750 175.620 4.890 177.340 ;
        RECT 4.690 175.300 4.950 175.620 ;
        RECT 6.530 174.620 6.790 174.940 ;
        RECT 6.590 173.580 6.730 174.620 ;
        RECT 6.530 173.260 6.790 173.580 ;
        RECT 8.890 173.540 9.030 183.460 ;
        RECT 10.670 183.120 10.930 183.440 ;
        RECT 10.730 178.340 10.870 183.120 ;
        RECT 11.190 180.380 11.330 185.500 ;
        RECT 11.130 180.290 11.390 180.380 ;
        RECT 11.130 180.150 11.790 180.290 ;
        RECT 11.130 180.060 11.390 180.150 ;
        RECT 10.670 178.020 10.930 178.340 ;
        RECT 11.650 175.280 11.790 180.150 ;
        RECT 11.590 174.960 11.850 175.280 ;
        RECT 8.890 173.400 9.490 173.540 ;
        RECT 4.230 169.520 4.490 169.840 ;
        RECT 4.290 164.740 4.430 169.520 ;
        RECT 5.610 169.180 5.870 169.500 ;
        RECT 8.830 169.180 9.090 169.500 ;
        RECT 5.670 168.140 5.810 169.180 ;
        RECT 5.610 167.820 5.870 168.140 ;
        RECT 4.230 164.420 4.490 164.740 ;
        RECT 8.890 164.060 9.030 169.180 ;
        RECT 8.830 163.740 9.090 164.060 ;
        RECT 8.890 161.000 9.030 163.740 ;
        RECT 8.830 160.680 9.090 161.000 ;
        RECT 8.890 158.620 9.030 160.680 ;
        RECT 8.830 158.300 9.090 158.620 ;
        RECT 4.230 153.200 4.490 153.520 ;
        RECT 4.290 148.080 4.430 153.200 ;
        RECT 6.070 152.860 6.330 153.180 ;
        RECT 5.610 150.820 5.870 151.140 ;
        RECT 5.140 148.245 5.420 148.615 ;
        RECT 4.230 147.760 4.490 148.080 ;
        RECT 4.290 142.980 4.430 147.760 ;
        RECT 4.690 147.080 4.950 147.400 ;
        RECT 4.230 142.660 4.490 142.980 ;
        RECT 3.770 140.280 4.030 140.600 ;
        RECT 4.290 137.540 4.430 142.660 ;
        RECT 4.230 137.220 4.490 137.540 ;
        RECT 4.750 134.140 4.890 147.080 ;
        RECT 5.210 145.700 5.350 148.245 ;
        RECT 5.150 145.380 5.410 145.700 ;
        RECT 5.150 144.360 5.410 144.680 ;
        RECT 5.210 135.500 5.350 144.360 ;
        RECT 5.670 139.580 5.810 150.820 ;
        RECT 6.130 148.420 6.270 152.860 ;
        RECT 7.910 151.500 8.170 151.820 ;
        RECT 7.970 151.140 8.110 151.500 ;
        RECT 8.830 151.160 9.090 151.480 ;
        RECT 7.450 150.820 7.710 151.140 ;
        RECT 7.910 150.820 8.170 151.140 ;
        RECT 6.070 148.100 6.330 148.420 ;
        RECT 7.510 145.700 7.650 150.820 ;
        RECT 8.370 150.140 8.630 150.460 ;
        RECT 8.430 146.380 8.570 150.140 ;
        RECT 8.890 150.120 9.030 151.160 ;
        RECT 8.830 149.800 9.090 150.120 ;
        RECT 8.370 146.060 8.630 146.380 ;
        RECT 6.990 145.380 7.250 145.700 ;
        RECT 7.450 145.380 7.710 145.700 ;
        RECT 7.910 145.380 8.170 145.700 ;
        RECT 8.820 145.525 9.100 145.895 ;
        RECT 7.050 143.660 7.190 145.380 ;
        RECT 6.990 143.340 7.250 143.660 ;
        RECT 6.070 142.320 6.330 142.640 ;
        RECT 5.610 139.260 5.870 139.580 ;
        RECT 5.610 136.540 5.870 136.860 ;
        RECT 5.150 135.180 5.410 135.500 ;
        RECT 4.690 133.820 4.950 134.140 ;
        RECT 5.150 133.820 5.410 134.140 ;
        RECT 5.210 132.100 5.350 133.820 ;
        RECT 5.670 132.780 5.810 136.540 ;
        RECT 6.130 135.500 6.270 142.320 ;
        RECT 7.450 140.850 7.710 140.940 ;
        RECT 7.970 140.850 8.110 145.380 ;
        RECT 8.370 144.700 8.630 145.020 ;
        RECT 7.450 140.710 8.110 140.850 ;
        RECT 7.450 140.620 7.710 140.710 ;
        RECT 8.430 135.500 8.570 144.700 ;
        RECT 8.890 140.260 9.030 145.525 ;
        RECT 9.350 140.600 9.490 173.400 ;
        RECT 12.570 172.560 12.710 196.040 ;
        RECT 12.970 193.320 13.230 193.640 ;
        RECT 13.030 191.600 13.170 193.320 ;
        RECT 12.970 191.280 13.230 191.600 ;
        RECT 13.490 188.880 13.630 199.780 ;
        RECT 14.810 199.440 15.070 199.760 ;
        RECT 14.870 198.060 15.010 199.440 ;
        RECT 15.270 198.760 15.530 199.080 ;
        RECT 14.810 197.740 15.070 198.060 ;
        RECT 14.350 197.400 14.610 197.720 ;
        RECT 14.410 197.040 14.550 197.400 ;
        RECT 14.350 196.720 14.610 197.040 ;
        RECT 15.330 196.780 15.470 198.760 ;
        RECT 17.170 198.060 17.310 205.220 ;
        RECT 17.630 203.500 17.770 205.220 ;
        RECT 17.570 203.180 17.830 203.500 ;
        RECT 18.090 202.820 18.230 206.920 ;
        RECT 18.490 205.560 18.750 205.880 ;
        RECT 18.030 202.500 18.290 202.820 ;
        RECT 18.550 199.080 18.690 205.560 ;
        RECT 18.940 201.965 19.220 202.335 ;
        RECT 18.950 201.820 19.210 201.965 ;
        RECT 19.010 200.780 19.150 201.820 ;
        RECT 19.930 201.655 20.070 209.640 ;
        RECT 20.850 208.340 20.990 212.360 ;
        RECT 24.990 211.320 25.130 212.700 ;
        RECT 24.930 211.000 25.190 211.320 ;
        RECT 26.770 209.640 27.030 209.960 ;
        RECT 21.415 209.105 22.955 209.475 ;
        RECT 21.240 208.340 21.520 208.455 ;
        RECT 20.850 208.200 21.520 208.340 ;
        RECT 21.240 208.085 21.520 208.200 ;
        RECT 21.710 207.940 21.970 208.260 ;
        RECT 23.090 207.940 23.350 208.260 ;
        RECT 20.330 206.920 20.590 207.240 ;
        RECT 20.390 206.220 20.530 206.920 ;
        RECT 20.330 205.900 20.590 206.220 ;
        RECT 21.770 205.735 21.910 207.940 ;
        RECT 21.700 205.365 21.980 205.735 ;
        RECT 20.330 204.880 20.590 205.200 ;
        RECT 20.390 202.140 20.530 204.880 ;
        RECT 21.240 204.685 21.520 205.055 ;
        RECT 21.250 204.540 21.510 204.685 ;
        RECT 21.415 203.665 22.955 204.035 ;
        RECT 20.790 202.840 21.050 203.160 ;
        RECT 20.330 201.820 20.590 202.140 ;
        RECT 19.860 201.285 20.140 201.655 ;
        RECT 19.930 200.780 20.070 201.285 ;
        RECT 18.950 200.460 19.210 200.780 ;
        RECT 19.870 200.460 20.130 200.780 ;
        RECT 19.870 199.440 20.130 199.760 ;
        RECT 18.490 198.760 18.750 199.080 ;
        RECT 17.110 197.740 17.370 198.060 ;
        RECT 14.410 196.100 14.550 196.720 ;
        RECT 14.870 196.700 15.470 196.780 ;
        RECT 14.810 196.640 15.470 196.700 ;
        RECT 14.810 196.380 15.070 196.640 ;
        RECT 14.410 195.960 15.470 196.100 ;
        RECT 17.570 196.040 17.830 196.360 ;
        RECT 18.030 196.040 18.290 196.360 ;
        RECT 19.410 196.040 19.670 196.360 ;
        RECT 13.890 194.340 14.150 194.660 ;
        RECT 13.950 189.560 14.090 194.340 ;
        RECT 14.350 191.280 14.610 191.600 ;
        RECT 13.890 189.240 14.150 189.560 ;
        RECT 13.430 188.560 13.690 188.880 ;
        RECT 13.430 186.180 13.690 186.500 ;
        RECT 12.970 185.160 13.230 185.480 ;
        RECT 13.030 183.780 13.170 185.160 ;
        RECT 12.970 183.460 13.230 183.780 ;
        RECT 13.490 178.000 13.630 186.180 ;
        RECT 13.950 185.820 14.090 189.240 ;
        RECT 14.410 188.200 14.550 191.280 ;
        RECT 14.350 187.880 14.610 188.200 ;
        RECT 13.890 185.500 14.150 185.820 ;
        RECT 13.890 183.120 14.150 183.440 ;
        RECT 13.950 181.740 14.090 183.120 ;
        RECT 13.890 181.420 14.150 181.740 ;
        RECT 14.350 180.400 14.610 180.720 ;
        RECT 13.890 179.720 14.150 180.040 ;
        RECT 13.950 178.680 14.090 179.720 ;
        RECT 14.410 179.020 14.550 180.400 ;
        RECT 14.350 178.700 14.610 179.020 ;
        RECT 13.890 178.360 14.150 178.680 ;
        RECT 14.810 178.020 15.070 178.340 ;
        RECT 13.430 177.680 13.690 178.000 ;
        RECT 13.490 172.560 13.630 177.680 ;
        RECT 13.890 175.640 14.150 175.960 ;
        RECT 13.950 173.580 14.090 175.640 ;
        RECT 13.890 173.260 14.150 173.580 ;
        RECT 12.510 172.240 12.770 172.560 ;
        RECT 13.430 172.240 13.690 172.560 ;
        RECT 10.670 171.620 10.930 171.880 ;
        RECT 10.270 171.560 10.930 171.620 ;
        RECT 10.270 171.480 10.870 171.560 ;
        RECT 10.270 167.460 10.410 171.480 ;
        RECT 10.210 167.140 10.470 167.460 ;
        RECT 10.270 157.260 10.410 167.140 ;
        RECT 11.590 166.800 11.850 167.120 ;
        RECT 10.670 164.760 10.930 165.080 ;
        RECT 10.730 162.020 10.870 164.760 ;
        RECT 11.650 164.740 11.790 166.800 ;
        RECT 11.590 164.420 11.850 164.740 ;
        RECT 11.650 162.360 11.790 164.420 ;
        RECT 11.590 162.040 11.850 162.360 ;
        RECT 10.670 161.700 10.930 162.020 ;
        RECT 10.730 158.960 10.870 161.700 ;
        RECT 10.670 158.640 10.930 158.960 ;
        RECT 10.210 156.940 10.470 157.260 ;
        RECT 10.730 156.580 10.870 158.640 ;
        RECT 10.670 156.260 10.930 156.580 ;
        RECT 10.210 155.240 10.470 155.560 ;
        RECT 10.270 152.015 10.410 155.240 ;
        RECT 10.200 151.645 10.480 152.015 ;
        RECT 9.750 150.710 10.010 150.800 ;
        RECT 9.750 150.570 10.410 150.710 ;
        RECT 9.750 150.480 10.010 150.570 ;
        RECT 9.740 144.845 10.020 145.215 ;
        RECT 9.810 140.940 9.950 144.845 ;
        RECT 10.270 142.640 10.410 150.570 ;
        RECT 10.210 142.320 10.470 142.640 ;
        RECT 9.750 140.620 10.010 140.940 ;
        RECT 9.290 140.280 9.550 140.600 ;
        RECT 8.830 139.940 9.090 140.260 ;
        RECT 10.270 139.920 10.410 142.320 ;
        RECT 10.210 139.600 10.470 139.920 ;
        RECT 6.070 135.180 6.330 135.500 ;
        RECT 8.370 135.180 8.630 135.500 ;
        RECT 10.730 135.160 10.870 156.260 ;
        RECT 11.130 150.480 11.390 150.800 ;
        RECT 11.190 148.080 11.330 150.480 ;
        RECT 11.130 147.760 11.390 148.080 ;
        RECT 11.190 142.300 11.330 147.760 ;
        RECT 11.650 145.360 11.790 162.040 ;
        RECT 12.570 159.640 12.710 172.240 ;
        RECT 14.870 170.860 15.010 178.020 ;
        RECT 14.810 170.540 15.070 170.860 ;
        RECT 14.350 169.520 14.610 169.840 ;
        RECT 12.970 168.840 13.230 169.160 ;
        RECT 13.030 167.460 13.170 168.840 ;
        RECT 14.410 168.140 14.550 169.520 ;
        RECT 14.810 169.180 15.070 169.500 ;
        RECT 14.350 167.820 14.610 168.140 ;
        RECT 12.970 167.140 13.230 167.460 ;
        RECT 12.970 165.100 13.230 165.420 ;
        RECT 13.030 162.700 13.170 165.100 ;
        RECT 13.890 163.400 14.150 163.720 ;
        RECT 13.950 162.700 14.090 163.400 ;
        RECT 12.970 162.380 13.230 162.700 ;
        RECT 13.890 162.380 14.150 162.700 ;
        RECT 13.890 161.360 14.150 161.680 ;
        RECT 12.510 159.320 12.770 159.640 ;
        RECT 12.050 155.920 12.310 156.240 ;
        RECT 12.110 154.540 12.250 155.920 ;
        RECT 12.050 154.220 12.310 154.540 ;
        RECT 12.570 154.200 12.710 159.320 ;
        RECT 12.970 156.940 13.230 157.260 ;
        RECT 12.510 153.880 12.770 154.200 ;
        RECT 12.570 146.040 12.710 153.880 ;
        RECT 13.030 147.400 13.170 156.940 ;
        RECT 13.950 148.760 14.090 161.360 ;
        RECT 14.870 153.180 15.010 169.180 ;
        RECT 15.330 153.180 15.470 195.960 ;
        RECT 17.110 194.000 17.370 194.320 ;
        RECT 15.730 191.620 15.990 191.940 ;
        RECT 15.790 186.840 15.930 191.620 ;
        RECT 16.190 190.600 16.450 190.920 ;
        RECT 16.650 190.600 16.910 190.920 ;
        RECT 15.730 186.520 15.990 186.840 ;
        RECT 15.730 175.300 15.990 175.620 ;
        RECT 15.790 155.560 15.930 175.300 ;
        RECT 16.250 164.140 16.390 190.600 ;
        RECT 16.710 189.220 16.850 190.600 ;
        RECT 16.650 188.900 16.910 189.220 ;
        RECT 17.170 187.180 17.310 194.000 ;
        RECT 17.110 186.860 17.370 187.180 ;
        RECT 17.630 186.500 17.770 196.040 ;
        RECT 18.090 191.600 18.230 196.040 ;
        RECT 18.490 195.020 18.750 195.340 ;
        RECT 18.030 191.280 18.290 191.600 ;
        RECT 17.570 186.180 17.830 186.500 ;
        RECT 18.090 186.160 18.230 191.280 ;
        RECT 18.550 187.180 18.690 195.020 ;
        RECT 18.950 194.000 19.210 194.320 ;
        RECT 19.010 193.640 19.150 194.000 ;
        RECT 19.470 193.640 19.610 196.040 ;
        RECT 18.950 193.320 19.210 193.640 ;
        RECT 19.410 193.320 19.670 193.640 ;
        RECT 18.950 188.560 19.210 188.880 ;
        RECT 18.490 186.860 18.750 187.180 ;
        RECT 18.030 185.900 18.290 186.160 ;
        RECT 19.010 185.900 19.150 188.560 ;
        RECT 16.710 185.840 18.290 185.900 ;
        RECT 16.710 185.760 18.230 185.840 ;
        RECT 18.550 185.760 19.150 185.900 ;
        RECT 16.710 171.880 16.850 185.760 ;
        RECT 18.030 185.160 18.290 185.480 ;
        RECT 17.570 182.440 17.830 182.760 ;
        RECT 17.630 181.740 17.770 182.440 ;
        RECT 17.110 181.420 17.370 181.740 ;
        RECT 17.570 181.420 17.830 181.740 ;
        RECT 17.170 179.020 17.310 181.420 ;
        RECT 17.110 178.700 17.370 179.020 ;
        RECT 17.170 175.280 17.310 178.700 ;
        RECT 17.110 174.960 17.370 175.280 ;
        RECT 17.630 173.540 17.770 181.420 ;
        RECT 18.090 175.280 18.230 185.160 ;
        RECT 18.550 178.000 18.690 185.760 ;
        RECT 19.470 183.180 19.610 193.320 ;
        RECT 19.930 184.460 20.070 199.440 ;
        RECT 20.330 197.060 20.590 197.380 ;
        RECT 20.390 192.280 20.530 197.060 ;
        RECT 20.850 197.040 20.990 202.840 ;
        RECT 22.160 201.965 22.440 202.335 ;
        RECT 23.150 202.220 23.290 207.940 ;
        RECT 26.830 207.920 26.970 209.640 ;
        RECT 26.770 207.600 27.030 207.920 ;
        RECT 27.290 207.580 27.430 216.100 ;
        RECT 27.750 210.980 27.890 218.820 ;
        RECT 30.910 217.975 31.170 218.120 ;
        RECT 30.900 217.605 31.180 217.975 ;
        RECT 29.070 216.100 29.330 216.420 ;
        RECT 28.150 215.080 28.410 215.400 ;
        RECT 28.210 211.320 28.350 215.080 ;
        RECT 28.150 211.000 28.410 211.320 ;
        RECT 27.690 210.660 27.950 210.980 ;
        RECT 27.230 207.260 27.490 207.580 ;
        RECT 24.010 206.920 24.270 207.240 ;
        RECT 24.470 206.920 24.730 207.240 ;
        RECT 26.310 206.920 26.570 207.240 ;
        RECT 26.770 206.920 27.030 207.240 ;
        RECT 24.070 206.220 24.210 206.920 ;
        RECT 23.550 205.900 23.810 206.220 ;
        RECT 24.010 205.900 24.270 206.220 ;
        RECT 23.610 205.620 23.750 205.900 ;
        RECT 23.610 205.480 24.210 205.620 ;
        RECT 23.550 204.880 23.810 205.200 ;
        RECT 22.690 202.080 23.290 202.220 ;
        RECT 22.170 201.820 22.430 201.965 ;
        RECT 22.230 200.100 22.370 201.820 ;
        RECT 22.690 200.440 22.830 202.080 ;
        RECT 23.090 201.480 23.350 201.800 ;
        RECT 22.630 200.120 22.890 200.440 ;
        RECT 22.170 199.780 22.430 200.100 ;
        RECT 21.415 198.225 22.955 198.595 ;
        RECT 20.790 196.720 21.050 197.040 ;
        RECT 23.150 196.780 23.290 201.480 ;
        RECT 23.610 199.080 23.750 204.880 ;
        RECT 24.070 204.860 24.210 205.480 ;
        RECT 24.010 204.540 24.270 204.860 ;
        RECT 24.530 203.500 24.670 206.920 ;
        RECT 26.370 206.220 26.510 206.920 ;
        RECT 26.310 205.900 26.570 206.220 ;
        RECT 25.390 205.450 25.650 205.540 ;
        RECT 25.390 205.310 26.510 205.450 ;
        RECT 25.390 205.220 25.650 205.310 ;
        RECT 24.930 204.200 25.190 204.520 ;
        RECT 24.990 203.500 25.130 204.200 ;
        RECT 24.470 203.180 24.730 203.500 ;
        RECT 24.930 203.180 25.190 203.500 ;
        RECT 24.930 202.730 25.190 202.820 ;
        RECT 24.930 202.590 25.590 202.730 ;
        RECT 24.930 202.500 25.190 202.590 ;
        RECT 24.010 201.480 24.270 201.800 ;
        RECT 23.550 198.760 23.810 199.080 ;
        RECT 23.610 197.720 23.750 198.760 ;
        RECT 23.550 197.400 23.810 197.720 ;
        RECT 22.690 196.700 23.290 196.780 ;
        RECT 22.630 196.640 23.290 196.700 ;
        RECT 22.630 196.380 22.890 196.640 ;
        RECT 20.790 196.040 21.050 196.360 ;
        RECT 20.330 191.960 20.590 192.280 ;
        RECT 20.390 188.880 20.530 191.960 ;
        RECT 20.330 188.560 20.590 188.880 ;
        RECT 20.330 185.160 20.590 185.480 ;
        RECT 19.870 184.140 20.130 184.460 ;
        RECT 19.010 183.040 19.610 183.180 ;
        RECT 18.490 177.680 18.750 178.000 ;
        RECT 18.030 174.960 18.290 175.280 ;
        RECT 17.630 173.400 18.230 173.540 ;
        RECT 16.650 171.560 16.910 171.880 ;
        RECT 18.090 170.860 18.230 173.400 ;
        RECT 19.010 172.900 19.150 183.040 ;
        RECT 19.410 179.720 19.670 180.040 ;
        RECT 19.470 174.940 19.610 179.720 ;
        RECT 19.410 174.620 19.670 174.940 ;
        RECT 19.870 174.620 20.130 174.940 ;
        RECT 19.470 173.580 19.610 174.620 ;
        RECT 19.410 173.260 19.670 173.580 ;
        RECT 19.930 173.240 20.070 174.620 ;
        RECT 20.390 173.240 20.530 185.160 ;
        RECT 20.850 183.440 20.990 196.040 ;
        RECT 23.550 194.340 23.810 194.660 ;
        RECT 21.415 192.785 22.955 193.155 ;
        RECT 23.090 190.600 23.350 190.920 ;
        RECT 21.415 187.345 22.955 187.715 ;
        RECT 23.150 185.480 23.290 190.600 ;
        RECT 23.610 189.980 23.750 194.340 ;
        RECT 24.070 193.640 24.210 201.480 ;
        RECT 24.470 198.760 24.730 199.080 ;
        RECT 24.010 193.320 24.270 193.640 ;
        RECT 23.610 189.840 24.210 189.980 ;
        RECT 24.070 189.220 24.210 189.840 ;
        RECT 24.010 189.130 24.270 189.220 ;
        RECT 23.610 188.990 24.270 189.130 ;
        RECT 21.250 185.160 21.510 185.480 ;
        RECT 23.090 185.160 23.350 185.480 ;
        RECT 20.790 183.120 21.050 183.440 ;
        RECT 21.310 182.670 21.450 185.160 ;
        RECT 23.610 184.460 23.750 188.990 ;
        RECT 24.010 188.900 24.270 188.990 ;
        RECT 24.010 185.500 24.270 185.820 ;
        RECT 24.070 184.460 24.210 185.500 ;
        RECT 23.550 184.140 23.810 184.460 ;
        RECT 24.010 184.140 24.270 184.460 ;
        RECT 20.850 182.530 21.450 182.670 ;
        RECT 22.630 182.670 22.890 182.760 ;
        RECT 22.630 182.530 23.290 182.670 ;
        RECT 20.850 181.740 20.990 182.530 ;
        RECT 22.630 182.440 22.890 182.530 ;
        RECT 21.415 181.905 22.955 182.275 ;
        RECT 20.790 181.420 21.050 181.740 ;
        RECT 20.790 177.680 21.050 178.000 ;
        RECT 20.850 176.300 20.990 177.680 ;
        RECT 21.415 176.465 22.955 176.835 ;
        RECT 20.790 175.980 21.050 176.300 ;
        RECT 23.150 175.620 23.290 182.530 ;
        RECT 23.610 180.040 23.750 184.140 ;
        RECT 24.530 183.860 24.670 198.760 ;
        RECT 25.450 197.575 25.590 202.590 ;
        RECT 26.370 201.800 26.510 205.310 ;
        RECT 26.830 202.480 26.970 206.920 ;
        RECT 27.230 204.880 27.490 205.200 ;
        RECT 27.290 203.500 27.430 204.880 ;
        RECT 27.230 203.180 27.490 203.500 ;
        RECT 27.290 203.015 27.430 203.180 ;
        RECT 27.220 202.645 27.500 203.015 ;
        RECT 26.770 202.160 27.030 202.480 ;
        RECT 26.310 201.480 26.570 201.800 ;
        RECT 25.380 197.205 25.660 197.575 ;
        RECT 25.450 197.040 25.590 197.205 ;
        RECT 25.390 196.720 25.650 197.040 ;
        RECT 25.850 196.720 26.110 197.040 ;
        RECT 25.910 195.340 26.050 196.720 ;
        RECT 25.850 195.020 26.110 195.340 ;
        RECT 26.370 193.980 26.510 201.480 ;
        RECT 27.290 200.180 27.430 202.645 ;
        RECT 26.830 200.040 27.430 200.180 ;
        RECT 26.310 193.660 26.570 193.980 ;
        RECT 25.850 193.320 26.110 193.640 ;
        RECT 25.910 191.940 26.050 193.320 ;
        RECT 24.930 191.620 25.190 191.940 ;
        RECT 25.850 191.620 26.110 191.940 ;
        RECT 24.990 188.200 25.130 191.620 ;
        RECT 25.850 190.600 26.110 190.920 ;
        RECT 24.930 187.880 25.190 188.200 ;
        RECT 24.070 183.720 24.670 183.860 ;
        RECT 23.550 179.720 23.810 180.040 ;
        RECT 23.610 178.680 23.750 179.720 ;
        RECT 23.550 178.360 23.810 178.680 ;
        RECT 24.070 177.910 24.210 183.720 ;
        RECT 24.470 183.120 24.730 183.440 ;
        RECT 24.530 181.740 24.670 183.120 ;
        RECT 24.470 181.420 24.730 181.740 ;
        RECT 23.610 177.770 24.210 177.910 ;
        RECT 23.090 175.300 23.350 175.620 ;
        RECT 21.250 174.960 21.510 175.280 ;
        RECT 20.790 174.280 21.050 174.600 ;
        RECT 19.870 172.920 20.130 173.240 ;
        RECT 20.330 172.920 20.590 173.240 ;
        RECT 18.950 172.580 19.210 172.900 ;
        RECT 17.110 170.540 17.370 170.860 ;
        RECT 18.030 170.540 18.290 170.860 ;
        RECT 17.170 167.120 17.310 170.540 ;
        RECT 19.930 170.260 20.070 172.920 ;
        RECT 17.570 169.860 17.830 170.180 ;
        RECT 19.930 170.120 20.530 170.260 ;
        RECT 17.110 166.800 17.370 167.120 ;
        RECT 16.250 164.060 16.850 164.140 ;
        RECT 16.250 164.000 16.910 164.060 ;
        RECT 16.650 163.740 16.910 164.000 ;
        RECT 16.180 155.725 16.460 156.095 ;
        RECT 15.730 155.240 15.990 155.560 ;
        RECT 14.810 152.860 15.070 153.180 ;
        RECT 15.270 152.860 15.530 153.180 ;
        RECT 15.790 152.840 15.930 155.240 ;
        RECT 15.730 152.520 15.990 152.840 ;
        RECT 14.340 151.645 14.620 152.015 ;
        RECT 13.890 148.440 14.150 148.760 ;
        RECT 14.410 148.080 14.550 151.645 ;
        RECT 14.810 148.440 15.070 148.760 ;
        RECT 14.350 147.760 14.610 148.080 ;
        RECT 13.890 147.420 14.150 147.740 ;
        RECT 12.970 147.080 13.230 147.400 ;
        RECT 12.510 145.720 12.770 146.040 ;
        RECT 11.590 145.040 11.850 145.360 ;
        RECT 11.130 142.210 11.390 142.300 ;
        RECT 11.130 142.070 11.790 142.210 ;
        RECT 11.130 141.980 11.390 142.070 ;
        RECT 11.650 137.540 11.790 142.070 ;
        RECT 11.590 137.220 11.850 137.540 ;
        RECT 10.670 134.840 10.930 135.160 ;
        RECT 5.610 132.460 5.870 132.780 ;
        RECT 5.150 131.780 5.410 132.100 ;
        RECT 10.210 131.780 10.470 132.100 ;
        RECT 6.990 131.100 7.250 131.420 ;
        RECT 7.050 128.700 7.190 131.100 ;
        RECT 10.270 130.060 10.410 131.780 ;
        RECT 11.650 131.670 11.790 137.220 ;
        RECT 12.050 136.880 12.310 137.200 ;
        RECT 12.110 136.520 12.250 136.880 ;
        RECT 12.050 136.200 12.310 136.520 ;
        RECT 12.110 134.820 12.250 136.200 ;
        RECT 12.050 134.500 12.310 134.820 ;
        RECT 12.050 131.670 12.310 131.760 ;
        RECT 11.650 131.530 12.310 131.670 ;
        RECT 12.050 131.440 12.310 131.530 ;
        RECT 10.210 129.740 10.470 130.060 ;
        RECT 8.370 129.060 8.630 129.380 ;
        RECT 6.990 128.380 7.250 128.700 ;
        RECT 8.430 127.340 8.570 129.060 ;
        RECT 11.590 128.720 11.850 129.040 ;
        RECT 11.650 127.340 11.790 128.720 ;
        RECT 8.370 127.020 8.630 127.340 ;
        RECT 11.590 127.020 11.850 127.340 ;
        RECT 12.570 125.980 12.710 145.720 ;
        RECT 13.030 135.500 13.170 147.080 ;
        RECT 13.950 145.700 14.090 147.420 ;
        RECT 14.870 147.310 15.010 148.440 ;
        RECT 14.410 147.170 15.010 147.310 ;
        RECT 14.410 145.700 14.550 147.170 ;
        RECT 13.890 145.380 14.150 145.700 ;
        RECT 14.350 145.380 14.610 145.700 ;
        RECT 14.410 141.960 14.550 145.380 ;
        RECT 15.790 145.360 15.930 152.520 ;
        RECT 14.810 145.040 15.070 145.360 ;
        RECT 15.270 145.040 15.530 145.360 ;
        RECT 15.730 145.040 15.990 145.360 ;
        RECT 14.870 143.660 15.010 145.040 ;
        RECT 14.810 143.340 15.070 143.660 ;
        RECT 13.890 141.640 14.150 141.960 ;
        RECT 14.350 141.640 14.610 141.960 ;
        RECT 13.430 139.940 13.690 140.260 ;
        RECT 13.490 139.150 13.630 139.940 ;
        RECT 13.950 139.920 14.090 141.640 ;
        RECT 14.870 141.020 15.010 143.340 ;
        RECT 14.410 140.940 15.010 141.020 ;
        RECT 14.350 140.880 15.010 140.940 ;
        RECT 14.350 140.620 14.610 140.880 ;
        RECT 13.890 139.600 14.150 139.920 ;
        RECT 13.490 139.010 14.550 139.150 ;
        RECT 14.410 137.880 14.550 139.010 ;
        RECT 14.350 137.560 14.610 137.880 ;
        RECT 14.350 136.200 14.610 136.520 ;
        RECT 14.410 135.500 14.550 136.200 ;
        RECT 12.970 135.180 13.230 135.500 ;
        RECT 14.350 135.180 14.610 135.500 ;
        RECT 13.430 134.840 13.690 135.160 ;
        RECT 12.970 133.480 13.230 133.800 ;
        RECT 13.030 131.670 13.170 133.480 ;
        RECT 13.490 132.180 13.630 134.840 ;
        RECT 13.890 132.180 14.150 132.440 ;
        RECT 13.490 132.120 14.150 132.180 ;
        RECT 13.490 132.040 14.090 132.120 ;
        RECT 14.350 131.780 14.610 132.100 ;
        RECT 13.890 131.670 14.150 131.760 ;
        RECT 13.030 131.530 14.150 131.670 ;
        RECT 13.890 131.440 14.150 131.530 ;
        RECT 13.950 126.660 14.090 131.440 ;
        RECT 14.410 126.660 14.550 131.780 ;
        RECT 15.330 131.760 15.470 145.040 ;
        RECT 16.250 132.100 16.390 155.725 ;
        RECT 16.710 136.520 16.850 163.740 ;
        RECT 17.170 161.680 17.310 166.800 ;
        RECT 17.630 165.080 17.770 169.860 ;
        RECT 19.410 166.800 19.670 167.120 ;
        RECT 17.570 164.760 17.830 165.080 ;
        RECT 18.490 163.400 18.750 163.720 ;
        RECT 18.550 162.700 18.690 163.400 ;
        RECT 18.490 162.380 18.750 162.700 ;
        RECT 17.110 161.360 17.370 161.680 ;
        RECT 17.570 160.680 17.830 161.000 ;
        RECT 17.630 156.580 17.770 160.680 ;
        RECT 19.470 159.980 19.610 166.800 ;
        RECT 19.870 166.120 20.130 166.440 ;
        RECT 19.410 159.660 19.670 159.980 ;
        RECT 19.930 159.740 20.070 166.120 ;
        RECT 20.390 165.420 20.530 170.120 ;
        RECT 20.330 165.100 20.590 165.420 ;
        RECT 20.320 164.565 20.600 164.935 ;
        RECT 20.390 164.400 20.530 164.565 ;
        RECT 20.850 164.400 20.990 174.280 ;
        RECT 21.310 172.900 21.450 174.960 ;
        RECT 22.630 174.620 22.890 174.940 ;
        RECT 22.690 173.240 22.830 174.620 ;
        RECT 23.150 173.240 23.290 175.300 ;
        RECT 22.630 172.920 22.890 173.240 ;
        RECT 23.090 172.920 23.350 173.240 ;
        RECT 21.250 172.580 21.510 172.900 ;
        RECT 23.150 172.560 23.290 172.920 ;
        RECT 23.090 172.240 23.350 172.560 ;
        RECT 23.090 171.560 23.350 171.880 ;
        RECT 21.415 171.025 22.955 171.395 ;
        RECT 22.630 170.540 22.890 170.860 ;
        RECT 22.170 170.200 22.430 170.520 ;
        RECT 22.230 168.140 22.370 170.200 ;
        RECT 22.170 167.820 22.430 168.140 ;
        RECT 22.690 167.540 22.830 170.540 ;
        RECT 23.150 168.140 23.290 171.560 ;
        RECT 23.090 167.820 23.350 168.140 ;
        RECT 22.690 167.400 23.290 167.540 ;
        RECT 21.415 165.585 22.955 165.955 ;
        RECT 20.330 164.080 20.590 164.400 ;
        RECT 20.790 164.080 21.050 164.400 ;
        RECT 21.415 160.145 22.955 160.515 ;
        RECT 19.470 156.920 19.610 159.660 ;
        RECT 19.930 159.600 20.990 159.740 ;
        RECT 20.850 158.620 20.990 159.600 ;
        RECT 22.630 158.640 22.890 158.960 ;
        RECT 20.790 158.300 21.050 158.620 ;
        RECT 22.690 157.260 22.830 158.640 ;
        RECT 22.630 156.940 22.890 157.260 ;
        RECT 19.410 156.600 19.670 156.920 ;
        RECT 17.570 156.260 17.830 156.580 ;
        RECT 20.790 155.920 21.050 156.240 ;
        RECT 18.030 155.580 18.290 155.900 ;
        RECT 17.110 152.520 17.370 152.840 ;
        RECT 17.170 146.380 17.310 152.520 ;
        RECT 17.570 150.480 17.830 150.800 ;
        RECT 17.110 146.060 17.370 146.380 ;
        RECT 17.110 145.610 17.370 145.700 ;
        RECT 17.630 145.610 17.770 150.480 ;
        RECT 17.110 145.470 17.770 145.610 ;
        RECT 17.110 145.380 17.370 145.470 ;
        RECT 18.090 145.020 18.230 155.580 ;
        RECT 19.870 155.240 20.130 155.560 ;
        RECT 19.930 154.540 20.070 155.240 ;
        RECT 20.850 154.540 20.990 155.920 ;
        RECT 23.150 155.560 23.290 167.400 ;
        RECT 23.610 158.960 23.750 177.770 ;
        RECT 24.470 174.620 24.730 174.940 ;
        RECT 24.010 172.240 24.270 172.560 ;
        RECT 24.070 170.860 24.210 172.240 ;
        RECT 24.010 170.540 24.270 170.860 ;
        RECT 24.070 164.400 24.210 170.540 ;
        RECT 24.530 169.160 24.670 174.620 ;
        RECT 24.470 168.840 24.730 169.160 ;
        RECT 24.470 167.140 24.730 167.460 ;
        RECT 24.530 166.780 24.670 167.140 ;
        RECT 24.470 166.460 24.730 166.780 ;
        RECT 24.470 165.100 24.730 165.420 ;
        RECT 24.010 164.080 24.270 164.400 ;
        RECT 24.010 163.400 24.270 163.720 ;
        RECT 23.550 158.640 23.810 158.960 ;
        RECT 23.550 157.960 23.810 158.280 ;
        RECT 23.610 157.455 23.750 157.960 ;
        RECT 23.540 157.085 23.820 157.455 ;
        RECT 24.070 156.240 24.210 163.400 ;
        RECT 24.530 162.020 24.670 165.100 ;
        RECT 24.990 162.700 25.130 187.880 ;
        RECT 25.910 180.720 26.050 190.600 ;
        RECT 25.850 180.400 26.110 180.720 ;
        RECT 25.840 175.445 26.120 175.815 ;
        RECT 25.910 174.600 26.050 175.445 ;
        RECT 25.850 174.280 26.110 174.600 ;
        RECT 25.390 172.580 25.650 172.900 ;
        RECT 25.450 167.030 25.590 172.580 ;
        RECT 25.850 167.710 26.110 167.800 ;
        RECT 26.370 167.710 26.510 193.660 ;
        RECT 26.830 193.640 26.970 200.040 ;
        RECT 27.230 199.615 27.490 199.760 ;
        RECT 27.220 199.245 27.500 199.615 ;
        RECT 26.770 193.320 27.030 193.640 ;
        RECT 26.760 191.765 27.040 192.135 ;
        RECT 27.750 191.940 27.890 210.660 ;
        RECT 28.150 206.920 28.410 207.240 ;
        RECT 28.210 203.500 28.350 206.920 ;
        RECT 28.610 204.880 28.870 205.200 ;
        RECT 28.670 203.500 28.810 204.880 ;
        RECT 28.150 203.180 28.410 203.500 ;
        RECT 28.610 203.180 28.870 203.500 ;
        RECT 29.130 200.780 29.270 216.100 ;
        RECT 31.430 216.080 31.570 218.820 ;
        RECT 31.890 218.120 32.030 219.500 ;
        RECT 45.170 218.820 45.430 219.140 ;
        RECT 48.850 218.820 49.110 219.140 ;
        RECT 33.210 218.480 33.470 218.800 ;
        RECT 31.830 217.800 32.090 218.120 ;
        RECT 31.370 215.760 31.630 216.080 ;
        RECT 30.450 215.080 30.710 215.400 ;
        RECT 29.990 207.600 30.250 207.920 ;
        RECT 30.050 207.240 30.190 207.600 ;
        RECT 29.990 206.920 30.250 207.240 ;
        RECT 29.520 204.685 29.800 205.055 ;
        RECT 29.070 200.460 29.330 200.780 ;
        RECT 28.150 200.120 28.410 200.440 ;
        RECT 28.210 198.060 28.350 200.120 ;
        RECT 29.590 199.500 29.730 204.685 ;
        RECT 30.050 201.800 30.190 206.920 ;
        RECT 30.510 202.480 30.650 215.080 ;
        RECT 30.910 210.320 31.170 210.640 ;
        RECT 30.970 206.130 31.110 210.320 ;
        RECT 31.430 208.260 31.570 215.760 ;
        RECT 31.890 215.255 32.030 217.800 ;
        RECT 32.280 216.925 32.560 217.295 ;
        RECT 33.270 217.100 33.410 218.480 ;
        RECT 34.590 218.140 34.850 218.460 ;
        RECT 35.050 218.140 35.310 218.460 ;
        RECT 36.430 218.140 36.690 218.460 ;
        RECT 36.890 218.140 37.150 218.460 ;
        RECT 32.290 216.780 32.550 216.925 ;
        RECT 33.210 216.780 33.470 217.100 ;
        RECT 31.820 214.885 32.100 215.255 ;
        RECT 32.350 212.680 32.490 216.780 ;
        RECT 34.650 216.420 34.790 218.140 ;
        RECT 35.110 216.760 35.250 218.140 ;
        RECT 35.970 217.800 36.230 218.120 ;
        RECT 35.050 216.440 35.310 216.760 ;
        RECT 34.590 216.100 34.850 216.420 ;
        RECT 34.650 212.680 34.790 216.100 ;
        RECT 36.030 213.700 36.170 217.800 ;
        RECT 36.490 216.080 36.630 218.140 ;
        RECT 36.430 215.760 36.690 216.080 ;
        RECT 35.970 213.380 36.230 213.700 ;
        RECT 32.290 212.360 32.550 212.680 ;
        RECT 34.590 212.360 34.850 212.680 ;
        RECT 34.650 211.320 34.790 212.360 ;
        RECT 34.590 211.000 34.850 211.320 ;
        RECT 33.210 210.320 33.470 210.640 ;
        RECT 32.740 208.765 33.020 209.135 ;
        RECT 31.370 207.940 31.630 208.260 ;
        RECT 32.810 207.240 32.950 208.765 ;
        RECT 33.270 207.775 33.410 210.320 ;
        RECT 34.650 209.960 34.790 211.000 ;
        RECT 34.590 209.640 34.850 209.960 ;
        RECT 33.200 207.405 33.480 207.775 ;
        RECT 33.210 207.260 33.470 207.405 ;
        RECT 32.750 206.920 33.010 207.240 ;
        RECT 31.370 206.130 31.630 206.220 ;
        RECT 30.970 205.990 31.630 206.130 ;
        RECT 30.970 202.480 31.110 205.990 ;
        RECT 31.370 205.900 31.630 205.990 ;
        RECT 32.290 204.200 32.550 204.520 ;
        RECT 30.450 202.160 30.710 202.480 ;
        RECT 30.910 202.160 31.170 202.480 ;
        RECT 32.350 202.335 32.490 204.200 ;
        RECT 29.990 201.480 30.250 201.800 ;
        RECT 28.670 199.360 29.730 199.500 ;
        RECT 28.150 197.740 28.410 198.060 ;
        RECT 28.150 196.040 28.410 196.360 ;
        RECT 28.210 195.000 28.350 196.040 ;
        RECT 28.150 194.680 28.410 195.000 ;
        RECT 26.830 191.600 26.970 191.765 ;
        RECT 27.690 191.620 27.950 191.940 ;
        RECT 26.770 191.280 27.030 191.600 ;
        RECT 26.830 189.900 26.970 191.280 ;
        RECT 26.770 189.580 27.030 189.900 ;
        RECT 27.750 187.180 27.890 191.620 ;
        RECT 28.150 190.940 28.410 191.260 ;
        RECT 27.690 186.860 27.950 187.180 ;
        RECT 27.750 183.780 27.890 186.860 ;
        RECT 28.210 184.460 28.350 190.940 ;
        RECT 28.150 184.140 28.410 184.460 ;
        RECT 27.690 183.460 27.950 183.780 ;
        RECT 26.770 181.420 27.030 181.740 ;
        RECT 26.830 173.580 26.970 181.420 ;
        RECT 27.750 181.060 27.890 183.460 ;
        RECT 27.690 180.740 27.950 181.060 ;
        RECT 27.750 179.020 27.890 180.740 ;
        RECT 27.690 178.700 27.950 179.020 ;
        RECT 28.150 177.680 28.410 178.000 ;
        RECT 27.230 175.640 27.490 175.960 ;
        RECT 27.290 174.940 27.430 175.640 ;
        RECT 28.210 175.280 28.350 177.680 ;
        RECT 28.150 174.960 28.410 175.280 ;
        RECT 27.230 174.620 27.490 174.940 ;
        RECT 26.770 173.260 27.030 173.580 ;
        RECT 26.760 172.725 27.040 173.095 ;
        RECT 26.830 171.880 26.970 172.725 ;
        RECT 26.770 171.560 27.030 171.880 ;
        RECT 25.850 167.570 26.510 167.710 ;
        RECT 25.850 167.480 26.110 167.570 ;
        RECT 26.770 167.480 27.030 167.800 ;
        RECT 25.450 166.890 26.050 167.030 ;
        RECT 25.390 163.400 25.650 163.720 ;
        RECT 24.930 162.380 25.190 162.700 ;
        RECT 24.470 161.700 24.730 162.020 ;
        RECT 24.530 161.340 24.670 161.700 ;
        RECT 24.470 161.020 24.730 161.340 ;
        RECT 24.010 155.920 24.270 156.240 ;
        RECT 23.090 155.240 23.350 155.560 ;
        RECT 24.010 155.240 24.270 155.560 ;
        RECT 21.415 154.705 22.955 155.075 ;
        RECT 19.870 154.220 20.130 154.540 ;
        RECT 20.790 154.220 21.050 154.540 ;
        RECT 21.250 154.220 21.510 154.540 ;
        RECT 19.410 153.540 19.670 153.860 ;
        RECT 18.490 151.500 18.750 151.820 ;
        RECT 18.030 144.700 18.290 145.020 ;
        RECT 18.550 142.980 18.690 151.500 ;
        RECT 18.950 149.800 19.210 150.120 ;
        RECT 19.010 149.100 19.150 149.800 ;
        RECT 18.950 148.780 19.210 149.100 ;
        RECT 18.950 148.330 19.210 148.420 ;
        RECT 19.470 148.330 19.610 153.540 ;
        RECT 21.310 153.180 21.450 154.220 ;
        RECT 21.250 152.860 21.510 153.180 ;
        RECT 23.550 152.860 23.810 153.180 ;
        RECT 23.090 152.520 23.350 152.840 ;
        RECT 20.320 151.645 20.600 152.015 ;
        RECT 19.870 150.140 20.130 150.460 ;
        RECT 18.950 148.190 19.610 148.330 ;
        RECT 18.950 148.100 19.210 148.190 ;
        RECT 18.490 142.660 18.750 142.980 ;
        RECT 19.010 142.890 19.150 148.100 ;
        RECT 19.410 147.080 19.670 147.400 ;
        RECT 19.470 146.575 19.610 147.080 ;
        RECT 19.400 146.205 19.680 146.575 ;
        RECT 19.930 146.380 20.070 150.140 ;
        RECT 19.870 146.060 20.130 146.380 ;
        RECT 20.390 144.680 20.530 151.645 ;
        RECT 21.415 149.265 22.955 149.635 ;
        RECT 20.790 147.760 21.050 148.080 ;
        RECT 20.330 144.360 20.590 144.680 ;
        RECT 20.390 143.320 20.530 144.360 ;
        RECT 20.330 143.000 20.590 143.320 ;
        RECT 19.410 142.890 19.670 142.980 ;
        RECT 19.010 142.750 19.670 142.890 ;
        RECT 19.410 142.660 19.670 142.750 ;
        RECT 18.550 140.850 18.690 142.660 ;
        RECT 18.950 140.850 19.210 140.940 ;
        RECT 18.550 140.710 19.210 140.850 ;
        RECT 18.950 140.620 19.210 140.710 ;
        RECT 19.470 139.920 19.610 142.660 ;
        RECT 19.860 142.125 20.140 142.495 ;
        RECT 19.870 141.980 20.130 142.125 ;
        RECT 20.850 141.960 20.990 147.760 ;
        RECT 22.630 147.420 22.890 147.740 ;
        RECT 22.690 145.360 22.830 147.420 ;
        RECT 22.630 145.215 22.890 145.360 ;
        RECT 22.620 144.845 22.900 145.215 ;
        RECT 21.415 143.825 22.955 144.195 ;
        RECT 21.250 143.340 21.510 143.660 ;
        RECT 20.790 141.640 21.050 141.960 ;
        RECT 21.310 140.260 21.450 143.340 ;
        RECT 23.150 142.640 23.290 152.520 ;
        RECT 23.610 150.120 23.750 152.860 ;
        RECT 23.550 149.800 23.810 150.120 ;
        RECT 24.070 148.760 24.210 155.240 ;
        RECT 24.530 154.540 24.670 161.020 ;
        RECT 24.930 159.320 25.190 159.640 ;
        RECT 24.990 156.580 25.130 159.320 ;
        RECT 24.930 156.260 25.190 156.580 ;
        RECT 24.930 155.240 25.190 155.560 ;
        RECT 24.470 154.220 24.730 154.540 ;
        RECT 24.470 149.800 24.730 150.120 ;
        RECT 24.530 149.100 24.670 149.800 ;
        RECT 24.470 148.780 24.730 149.100 ;
        RECT 24.010 148.440 24.270 148.760 ;
        RECT 24.010 147.760 24.270 148.080 ;
        RECT 23.550 147.080 23.810 147.400 ;
        RECT 23.090 142.320 23.350 142.640 ;
        RECT 20.330 139.940 20.590 140.260 ;
        RECT 21.250 139.940 21.510 140.260 ;
        RECT 23.090 139.940 23.350 140.260 ;
        RECT 19.410 139.600 19.670 139.920 ;
        RECT 18.950 138.920 19.210 139.240 ;
        RECT 16.650 136.200 16.910 136.520 ;
        RECT 16.710 134.480 16.850 136.200 ;
        RECT 16.650 134.160 16.910 134.480 ;
        RECT 16.190 131.780 16.450 132.100 ;
        RECT 15.270 131.440 15.530 131.760 ;
        RECT 16.710 131.080 16.850 134.160 ;
        RECT 16.190 130.760 16.450 131.080 ;
        RECT 16.650 130.760 16.910 131.080 ;
        RECT 18.490 130.760 18.750 131.080 ;
        RECT 16.250 127.340 16.390 130.760 ;
        RECT 18.550 127.340 18.690 130.760 ;
        RECT 19.010 129.040 19.150 138.920 ;
        RECT 19.470 137.540 19.610 139.600 ;
        RECT 19.410 137.220 19.670 137.540 ;
        RECT 20.390 136.520 20.530 139.940 ;
        RECT 20.790 138.920 21.050 139.240 ;
        RECT 20.850 137.540 20.990 138.920 ;
        RECT 21.415 138.385 22.955 138.755 ;
        RECT 20.790 137.220 21.050 137.540 ;
        RECT 20.330 136.200 20.590 136.520 ;
        RECT 20.390 135.160 20.530 136.200 ;
        RECT 23.150 135.500 23.290 139.940 ;
        RECT 23.610 136.860 23.750 147.080 ;
        RECT 24.070 145.610 24.210 147.760 ;
        RECT 24.470 147.650 24.730 147.740 ;
        RECT 24.990 147.650 25.130 155.240 ;
        RECT 24.470 147.510 25.130 147.650 ;
        RECT 24.470 147.420 24.730 147.510 ;
        RECT 24.070 145.470 24.670 145.610 ;
        RECT 24.010 144.700 24.270 145.020 ;
        RECT 24.070 143.060 24.210 144.700 ;
        RECT 24.530 143.570 24.670 145.470 ;
        RECT 24.930 145.380 25.190 145.700 ;
        RECT 24.990 144.535 25.130 145.380 ;
        RECT 25.450 144.680 25.590 163.400 ;
        RECT 25.910 159.495 26.050 166.890 ;
        RECT 26.300 166.605 26.580 166.975 ;
        RECT 26.370 162.700 26.510 166.605 ;
        RECT 26.830 163.720 26.970 167.480 ;
        RECT 26.770 163.400 27.030 163.720 ;
        RECT 26.310 162.380 26.570 162.700 ;
        RECT 26.830 162.020 26.970 163.400 ;
        RECT 26.770 161.700 27.030 162.020 ;
        RECT 25.840 159.125 26.120 159.495 ;
        RECT 25.910 158.960 26.050 159.125 ;
        RECT 25.850 158.640 26.110 158.960 ;
        RECT 26.310 157.960 26.570 158.280 ;
        RECT 25.850 156.260 26.110 156.580 ;
        RECT 25.910 156.095 26.050 156.260 ;
        RECT 25.840 155.725 26.120 156.095 ;
        RECT 25.850 155.240 26.110 155.560 ;
        RECT 25.910 154.540 26.050 155.240 ;
        RECT 25.850 154.220 26.110 154.540 ;
        RECT 25.850 152.520 26.110 152.840 ;
        RECT 24.920 144.165 25.200 144.535 ;
        RECT 25.390 144.360 25.650 144.680 ;
        RECT 24.530 143.430 25.130 143.570 ;
        RECT 24.070 142.920 24.670 143.060 ;
        RECT 24.010 142.320 24.270 142.640 ;
        RECT 24.070 140.940 24.210 142.320 ;
        RECT 24.010 140.620 24.270 140.940 ;
        RECT 24.530 139.660 24.670 142.920 ;
        RECT 24.070 139.520 24.670 139.660 ;
        RECT 24.990 139.580 25.130 143.430 ;
        RECT 25.910 142.640 26.050 152.520 ;
        RECT 26.370 151.140 26.510 157.960 ;
        RECT 26.830 152.840 26.970 161.700 ;
        RECT 27.290 158.620 27.430 174.620 ;
        RECT 28.150 167.140 28.410 167.460 ;
        RECT 27.690 166.120 27.950 166.440 ;
        RECT 27.750 165.420 27.890 166.120 ;
        RECT 27.690 165.100 27.950 165.420 ;
        RECT 27.230 158.300 27.490 158.620 ;
        RECT 27.690 157.170 27.950 157.260 ;
        RECT 28.210 157.170 28.350 167.140 ;
        RECT 27.690 157.030 28.350 157.170 ;
        RECT 27.690 156.940 27.950 157.030 ;
        RECT 27.750 153.180 27.890 156.940 ;
        RECT 28.670 156.775 28.810 199.360 ;
        RECT 29.530 198.760 29.790 199.080 ;
        RECT 29.590 198.060 29.730 198.760 ;
        RECT 29.530 197.740 29.790 198.060 ;
        RECT 30.970 197.380 31.110 202.160 ;
        RECT 32.280 201.965 32.560 202.335 ;
        RECT 32.290 199.440 32.550 199.760 ;
        RECT 30.910 197.060 31.170 197.380 ;
        RECT 30.450 190.940 30.710 191.260 ;
        RECT 30.510 189.900 30.650 190.940 ;
        RECT 30.970 189.900 31.110 197.060 ;
        RECT 30.450 189.580 30.710 189.900 ;
        RECT 30.910 189.580 31.170 189.900 ;
        RECT 31.370 185.160 31.630 185.480 ;
        RECT 30.450 184.140 30.710 184.460 ;
        RECT 29.070 180.060 29.330 180.380 ;
        RECT 29.130 179.020 29.270 180.060 ;
        RECT 29.070 178.700 29.330 179.020 ;
        RECT 29.990 171.560 30.250 171.880 ;
        RECT 30.050 170.180 30.190 171.560 ;
        RECT 29.990 169.860 30.250 170.180 ;
        RECT 29.070 168.840 29.330 169.160 ;
        RECT 29.130 167.460 29.270 168.840 ;
        RECT 29.070 167.370 29.330 167.460 ;
        RECT 29.070 167.230 29.730 167.370 ;
        RECT 29.070 167.140 29.330 167.230 ;
        RECT 29.070 166.460 29.330 166.780 ;
        RECT 28.600 156.405 28.880 156.775 ;
        RECT 28.150 155.920 28.410 156.240 ;
        RECT 28.210 153.375 28.350 155.920 ;
        RECT 27.690 152.860 27.950 153.180 ;
        RECT 28.140 153.005 28.420 153.375 ;
        RECT 26.770 152.520 27.030 152.840 ;
        RECT 26.310 150.820 26.570 151.140 ;
        RECT 26.770 150.820 27.030 151.140 ;
        RECT 27.230 150.820 27.490 151.140 ;
        RECT 26.310 150.140 26.570 150.460 ;
        RECT 26.370 146.380 26.510 150.140 ;
        RECT 26.310 146.060 26.570 146.380 ;
        RECT 26.310 145.380 26.570 145.700 ;
        RECT 26.370 144.680 26.510 145.380 ;
        RECT 26.310 144.360 26.570 144.680 ;
        RECT 26.830 143.660 26.970 150.820 ;
        RECT 27.290 150.655 27.430 150.820 ;
        RECT 27.220 150.285 27.500 150.655 ;
        RECT 27.230 149.975 27.490 150.120 ;
        RECT 27.220 149.605 27.500 149.975 ;
        RECT 27.230 148.100 27.490 148.420 ;
        RECT 27.290 147.255 27.430 148.100 ;
        RECT 27.220 146.885 27.500 147.255 ;
        RECT 27.290 145.895 27.430 146.885 ;
        RECT 27.750 146.380 27.890 152.860 ;
        RECT 28.670 151.140 28.810 156.405 ;
        RECT 29.130 151.140 29.270 166.460 ;
        RECT 29.590 165.420 29.730 167.230 ;
        RECT 29.530 165.100 29.790 165.420 ;
        RECT 30.510 158.815 30.650 184.140 ;
        RECT 31.430 183.780 31.570 185.160 ;
        RECT 31.370 183.460 31.630 183.780 ;
        RECT 31.830 180.740 32.090 181.060 ;
        RECT 31.890 178.340 32.030 180.740 ;
        RECT 31.370 178.020 31.630 178.340 ;
        RECT 31.830 178.020 32.090 178.340 ;
        RECT 31.430 176.300 31.570 178.020 ;
        RECT 31.370 175.980 31.630 176.300 ;
        RECT 32.350 175.700 32.490 199.440 ;
        RECT 32.810 188.620 32.950 206.920 ;
        RECT 34.650 205.200 34.790 209.640 ;
        RECT 36.950 207.920 37.090 218.140 ;
        RECT 44.710 217.800 44.970 218.120 ;
        RECT 40.850 217.265 42.390 217.635 ;
        RECT 44.770 217.100 44.910 217.800 ;
        RECT 45.230 217.100 45.370 218.820 ;
        RECT 48.390 218.480 48.650 218.800 ;
        RECT 45.630 217.800 45.890 218.120 ;
        RECT 44.710 216.780 44.970 217.100 ;
        RECT 45.170 216.780 45.430 217.100 ;
        RECT 45.170 215.760 45.430 216.080 ;
        RECT 39.640 214.205 39.920 214.575 ;
        RECT 43.320 214.205 43.600 214.575 ;
        RECT 39.180 213.525 39.460 213.895 ;
        RECT 39.190 213.380 39.450 213.525 ;
        RECT 39.190 212.360 39.450 212.680 ;
        RECT 37.350 211.000 37.610 211.320 ;
        RECT 36.890 207.600 37.150 207.920 ;
        RECT 37.410 207.240 37.550 211.000 ;
        RECT 39.250 210.980 39.390 212.360 ;
        RECT 39.190 210.660 39.450 210.980 ;
        RECT 39.710 208.600 39.850 214.205 ;
        RECT 43.330 214.060 43.590 214.205 ;
        RECT 40.110 213.720 40.370 214.040 ;
        RECT 39.650 208.280 39.910 208.600 ;
        RECT 40.170 207.920 40.310 213.720 ;
        RECT 45.230 213.020 45.370 215.760 ;
        RECT 44.250 212.700 44.510 213.020 ;
        RECT 45.170 212.700 45.430 213.020 ;
        RECT 42.870 212.360 43.130 212.680 ;
        RECT 40.850 211.825 42.390 212.195 ;
        RECT 40.110 207.600 40.370 207.920 ;
        RECT 39.650 207.260 39.910 207.580 ;
        RECT 37.350 206.920 37.610 207.240 ;
        RECT 34.590 204.880 34.850 205.200 ;
        RECT 34.130 200.460 34.390 200.780 ;
        RECT 33.670 198.760 33.930 199.080 ;
        RECT 33.200 194.485 33.480 194.855 ;
        RECT 33.270 189.900 33.410 194.485 ;
        RECT 33.210 189.580 33.470 189.900 ;
        RECT 33.730 189.220 33.870 198.760 ;
        RECT 34.190 189.220 34.330 200.460 ;
        RECT 34.650 197.040 34.790 204.880 ;
        RECT 36.890 204.200 37.150 204.520 ;
        RECT 35.970 201.480 36.230 201.800 ;
        RECT 36.030 200.440 36.170 201.480 ;
        RECT 35.970 200.120 36.230 200.440 ;
        RECT 35.510 199.440 35.770 199.760 ;
        RECT 34.590 196.720 34.850 197.040 ;
        RECT 35.570 194.320 35.710 199.440 ;
        RECT 35.510 194.000 35.770 194.320 ;
        RECT 33.670 188.900 33.930 189.220 ;
        RECT 34.130 188.900 34.390 189.220 ;
        RECT 35.050 189.130 35.310 189.220 ;
        RECT 35.570 189.130 35.710 194.000 ;
        RECT 35.050 188.990 35.710 189.130 ;
        RECT 35.050 188.900 35.310 188.990 ;
        RECT 32.810 188.480 33.870 188.620 ;
        RECT 31.430 175.560 32.490 175.700 ;
        RECT 31.430 173.580 31.570 175.560 ;
        RECT 32.750 174.280 33.010 174.600 ;
        RECT 31.370 173.260 31.630 173.580 ;
        RECT 30.910 166.800 31.170 167.120 ;
        RECT 30.970 164.740 31.110 166.800 ;
        RECT 31.430 165.330 31.570 173.260 ;
        RECT 31.830 172.920 32.090 173.240 ;
        RECT 31.890 170.180 32.030 172.920 ;
        RECT 31.830 170.090 32.090 170.180 ;
        RECT 31.830 169.950 32.490 170.090 ;
        RECT 31.830 169.860 32.090 169.950 ;
        RECT 31.430 165.190 32.030 165.330 ;
        RECT 30.910 164.420 31.170 164.740 ;
        RECT 31.370 164.420 31.630 164.740 ;
        RECT 31.430 159.980 31.570 164.420 ;
        RECT 31.370 159.660 31.630 159.980 ;
        RECT 30.900 159.125 31.180 159.495 ;
        RECT 30.440 158.700 30.720 158.815 ;
        RECT 30.050 158.560 30.720 158.700 ;
        RECT 28.610 150.820 28.870 151.140 ;
        RECT 29.070 150.820 29.330 151.140 ;
        RECT 29.520 150.965 29.800 151.335 ;
        RECT 28.610 149.800 28.870 150.120 ;
        RECT 28.150 147.420 28.410 147.740 ;
        RECT 27.690 146.060 27.950 146.380 ;
        RECT 27.220 145.525 27.500 145.895 ;
        RECT 27.220 144.845 27.500 145.215 ;
        RECT 27.690 145.040 27.950 145.360 ;
        RECT 27.230 144.700 27.490 144.845 ;
        RECT 27.750 143.660 27.890 145.040 ;
        RECT 26.770 143.340 27.030 143.660 ;
        RECT 27.690 143.340 27.950 143.660 ;
        RECT 28.210 142.640 28.350 147.420 ;
        RECT 28.670 145.020 28.810 149.800 ;
        RECT 29.590 149.100 29.730 150.965 ;
        RECT 29.530 148.780 29.790 149.100 ;
        RECT 29.070 147.760 29.330 148.080 ;
        RECT 29.130 146.040 29.270 147.760 ;
        RECT 29.070 145.720 29.330 146.040 ;
        RECT 29.070 145.040 29.330 145.360 ;
        RECT 28.610 144.700 28.870 145.020 ;
        RECT 29.130 143.855 29.270 145.040 ;
        RECT 29.060 143.485 29.340 143.855 ;
        RECT 25.850 142.320 26.110 142.640 ;
        RECT 28.150 142.320 28.410 142.640 ;
        RECT 25.850 141.640 26.110 141.960 ;
        RECT 25.910 140.940 26.050 141.640 ;
        RECT 25.850 140.620 26.110 140.940 ;
        RECT 26.310 139.940 26.570 140.260 ;
        RECT 24.070 138.220 24.210 139.520 ;
        RECT 24.930 139.260 25.190 139.580 ;
        RECT 24.470 138.920 24.730 139.240 ;
        RECT 24.010 137.900 24.270 138.220 ;
        RECT 24.010 137.220 24.270 137.540 ;
        RECT 23.550 136.540 23.810 136.860 ;
        RECT 23.090 135.180 23.350 135.500 ;
        RECT 20.330 134.840 20.590 135.160 ;
        RECT 19.410 133.820 19.670 134.140 ;
        RECT 19.470 132.440 19.610 133.820 ;
        RECT 19.410 132.120 19.670 132.440 ;
        RECT 19.470 129.380 19.610 132.120 ;
        RECT 20.390 131.760 20.530 134.840 ;
        RECT 23.090 133.480 23.350 133.800 ;
        RECT 21.415 132.945 22.955 133.315 ;
        RECT 23.150 132.780 23.290 133.480 ;
        RECT 23.090 132.460 23.350 132.780 ;
        RECT 20.330 131.440 20.590 131.760 ;
        RECT 22.630 131.440 22.890 131.760 ;
        RECT 20.390 129.720 20.530 131.440 ;
        RECT 21.250 130.760 21.510 131.080 ;
        RECT 21.310 129.720 21.450 130.760 ;
        RECT 22.690 130.060 22.830 131.440 ;
        RECT 24.070 130.060 24.210 137.220 ;
        RECT 24.530 131.420 24.670 138.920 ;
        RECT 26.370 135.500 26.510 139.940 ;
        RECT 26.310 135.180 26.570 135.500 ;
        RECT 24.470 131.100 24.730 131.420 ;
        RECT 22.630 129.740 22.890 130.060 ;
        RECT 24.010 129.740 24.270 130.060 ;
        RECT 20.330 129.400 20.590 129.720 ;
        RECT 21.250 129.400 21.510 129.720 ;
        RECT 19.410 129.060 19.670 129.380 ;
        RECT 28.210 129.040 28.350 142.320 ;
        RECT 30.050 140.940 30.190 158.560 ;
        RECT 30.440 158.445 30.720 158.560 ;
        RECT 30.440 155.045 30.720 155.415 ;
        RECT 30.510 148.080 30.650 155.045 ;
        RECT 30.970 148.080 31.110 159.125 ;
        RECT 31.890 156.920 32.030 165.190 ;
        RECT 32.350 159.640 32.490 169.950 ;
        RECT 32.810 169.500 32.950 174.280 ;
        RECT 32.750 169.180 33.010 169.500 ;
        RECT 32.810 167.800 32.950 169.180 ;
        RECT 32.750 167.480 33.010 167.800 ;
        RECT 32.740 163.885 33.020 164.255 ;
        RECT 32.810 159.640 32.950 163.885 ;
        RECT 32.290 159.320 32.550 159.640 ;
        RECT 32.750 159.320 33.010 159.640 ;
        RECT 32.290 158.640 32.550 158.960 ;
        RECT 31.830 156.600 32.090 156.920 ;
        RECT 32.350 156.580 32.490 158.640 ;
        RECT 32.290 156.260 32.550 156.580 ;
        RECT 31.370 155.920 31.630 156.240 ;
        RECT 31.830 155.920 32.090 156.240 ;
        RECT 31.430 154.540 31.570 155.920 ;
        RECT 31.370 154.220 31.630 154.540 ;
        RECT 31.890 150.540 32.030 155.920 ;
        RECT 32.350 152.015 32.490 156.260 ;
        RECT 33.730 155.980 33.870 188.480 ;
        RECT 34.190 186.500 34.330 188.900 ;
        RECT 34.130 186.180 34.390 186.500 ;
        RECT 34.590 185.840 34.850 186.160 ;
        RECT 34.650 180.720 34.790 185.840 ;
        RECT 35.110 182.760 35.250 188.900 ;
        RECT 35.510 185.160 35.770 185.480 ;
        RECT 35.570 184.460 35.710 185.160 ;
        RECT 35.510 184.140 35.770 184.460 ;
        RECT 35.510 183.460 35.770 183.780 ;
        RECT 35.050 182.440 35.310 182.760 ;
        RECT 35.570 181.820 35.710 183.460 ;
        RECT 35.110 181.680 35.710 181.820 ;
        RECT 34.590 180.400 34.850 180.720 ;
        RECT 34.650 178.680 34.790 180.400 ;
        RECT 34.590 178.360 34.850 178.680 ;
        RECT 34.590 175.300 34.850 175.620 ;
        RECT 34.130 168.840 34.390 169.160 ;
        RECT 34.190 166.440 34.330 168.840 ;
        RECT 34.130 166.120 34.390 166.440 ;
        RECT 34.190 164.400 34.330 166.120 ;
        RECT 34.650 164.740 34.790 175.300 ;
        RECT 34.590 164.420 34.850 164.740 ;
        RECT 34.130 164.080 34.390 164.400 ;
        RECT 34.650 161.535 34.790 164.420 ;
        RECT 35.110 162.700 35.250 181.680 ;
        RECT 35.510 174.620 35.770 174.940 ;
        RECT 35.570 169.695 35.710 174.620 ;
        RECT 35.500 169.325 35.780 169.695 ;
        RECT 36.030 167.540 36.170 200.120 ;
        RECT 36.950 200.010 37.090 204.200 ;
        RECT 37.410 202.140 37.550 206.920 ;
        RECT 39.190 205.560 39.450 205.880 ;
        RECT 38.260 202.645 38.540 203.015 ;
        RECT 37.350 201.820 37.610 202.140 ;
        RECT 37.350 200.010 37.610 200.100 ;
        RECT 36.950 199.870 37.610 200.010 ;
        RECT 37.350 199.780 37.610 199.870 ;
        RECT 36.430 199.440 36.690 199.760 ;
        RECT 36.490 191.940 36.630 199.440 ;
        RECT 36.890 194.680 37.150 195.000 ;
        RECT 36.430 191.620 36.690 191.940 ;
        RECT 36.950 191.600 37.090 194.680 ;
        RECT 36.890 191.280 37.150 191.600 ;
        RECT 36.950 186.160 37.090 191.280 ;
        RECT 36.890 185.840 37.150 186.160 ;
        RECT 37.410 183.780 37.550 199.780 ;
        RECT 38.330 197.380 38.470 202.645 ;
        RECT 38.730 201.820 38.990 202.140 ;
        RECT 38.790 200.780 38.930 201.820 ;
        RECT 39.250 201.800 39.390 205.560 ;
        RECT 39.190 201.480 39.450 201.800 ;
        RECT 38.730 200.460 38.990 200.780 ;
        RECT 39.190 198.935 39.450 199.080 ;
        RECT 39.180 198.565 39.460 198.935 ;
        RECT 38.270 197.060 38.530 197.380 ;
        RECT 37.810 183.800 38.070 184.120 ;
        RECT 37.350 183.460 37.610 183.780 ;
        RECT 36.430 183.120 36.690 183.440 ;
        RECT 35.570 167.400 36.170 167.540 ;
        RECT 35.050 162.380 35.310 162.700 ;
        RECT 35.050 161.700 35.310 162.020 ;
        RECT 34.580 161.165 34.860 161.535 ;
        RECT 34.590 160.680 34.850 161.000 ;
        RECT 33.270 155.840 33.870 155.980 ;
        RECT 32.280 151.645 32.560 152.015 ;
        RECT 32.290 150.820 32.550 151.140 ;
        RECT 31.430 150.400 32.030 150.540 ;
        RECT 32.350 150.540 32.490 150.820 ;
        RECT 33.270 150.540 33.410 155.840 ;
        RECT 34.130 155.580 34.390 155.900 ;
        RECT 34.190 154.540 34.330 155.580 ;
        RECT 34.130 154.220 34.390 154.540 ;
        RECT 33.660 153.685 33.940 154.055 ;
        RECT 33.730 152.840 33.870 153.685 ;
        RECT 34.650 153.520 34.790 160.680 ;
        RECT 35.110 159.980 35.250 161.700 ;
        RECT 35.050 159.660 35.310 159.980 ;
        RECT 35.050 158.870 35.310 158.960 ;
        RECT 35.570 158.870 35.710 167.400 ;
        RECT 35.970 166.460 36.230 166.780 ;
        RECT 36.030 158.960 36.170 166.460 ;
        RECT 35.050 158.730 35.710 158.870 ;
        RECT 35.050 158.640 35.310 158.730 ;
        RECT 35.970 158.640 36.230 158.960 ;
        RECT 36.490 158.190 36.630 183.120 ;
        RECT 37.350 182.440 37.610 182.760 ;
        RECT 37.410 181.060 37.550 182.440 ;
        RECT 37.350 180.740 37.610 181.060 ;
        RECT 37.870 180.040 38.010 183.800 ;
        RECT 38.330 183.440 38.470 197.060 ;
        RECT 39.710 197.040 39.850 207.260 ;
        RECT 40.850 206.385 42.390 206.755 ;
        RECT 41.950 206.130 42.210 206.220 ;
        RECT 42.930 206.130 43.070 212.360 ;
        RECT 43.330 206.920 43.590 207.240 ;
        RECT 43.390 206.220 43.530 206.920 ;
        RECT 41.950 205.990 43.070 206.130 ;
        RECT 41.950 205.900 42.210 205.990 ;
        RECT 43.330 205.900 43.590 206.220 ;
        RECT 42.010 205.540 42.150 205.900 ;
        RECT 41.950 205.220 42.210 205.540 ;
        RECT 43.330 205.220 43.590 205.540 ;
        RECT 41.490 202.840 41.750 203.160 ;
        RECT 41.550 202.050 41.690 202.840 ;
        RECT 42.010 202.820 42.150 205.220 ;
        RECT 43.390 204.520 43.530 205.220 ;
        RECT 43.330 204.200 43.590 204.520 ;
        RECT 41.950 202.500 42.210 202.820 ;
        RECT 40.170 201.910 41.690 202.050 ;
        RECT 40.170 200.780 40.310 201.910 ;
        RECT 42.870 201.820 43.130 202.140 ;
        RECT 42.930 201.655 43.070 201.820 ;
        RECT 40.850 200.945 42.390 201.315 ;
        RECT 42.860 201.285 43.140 201.655 ;
        RECT 40.110 200.460 40.370 200.780 ;
        RECT 43.330 200.460 43.590 200.780 ;
        RECT 40.560 199.925 40.840 200.295 ;
        RECT 41.490 200.120 41.750 200.440 ;
        RECT 40.630 198.060 40.770 199.925 ;
        RECT 41.030 198.760 41.290 199.080 ;
        RECT 41.090 198.060 41.230 198.760 ;
        RECT 40.570 197.740 40.830 198.060 ;
        RECT 41.030 197.740 41.290 198.060 ;
        RECT 41.550 197.040 41.690 200.120 ;
        RECT 43.390 199.670 43.530 200.460 ;
        RECT 43.790 199.780 44.050 200.100 ;
        RECT 42.930 199.530 43.530 199.670 ;
        RECT 42.410 199.100 42.670 199.420 ;
        RECT 39.650 196.720 39.910 197.040 ;
        RECT 41.490 196.950 41.750 197.040 ;
        RECT 40.170 196.810 41.750 196.950 ;
        RECT 42.470 196.895 42.610 199.100 ;
        RECT 38.730 196.040 38.990 196.360 ;
        RECT 39.190 196.040 39.450 196.360 ;
        RECT 38.790 195.340 38.930 196.040 ;
        RECT 38.730 195.020 38.990 195.340 ;
        RECT 39.250 194.660 39.390 196.040 ;
        RECT 39.190 194.340 39.450 194.660 ;
        RECT 38.730 191.620 38.990 191.940 ;
        RECT 38.270 183.120 38.530 183.440 ;
        RECT 38.330 180.575 38.470 183.120 ;
        RECT 38.260 180.205 38.540 180.575 ;
        RECT 36.890 179.720 37.150 180.040 ;
        RECT 37.810 179.720 38.070 180.040 ;
        RECT 36.950 177.320 37.090 179.720 ;
        RECT 36.890 177.000 37.150 177.320 ;
        RECT 36.890 172.580 37.150 172.900 ;
        RECT 36.950 170.520 37.090 172.580 ;
        RECT 37.350 172.240 37.610 172.560 ;
        RECT 36.890 170.200 37.150 170.520 ;
        RECT 36.950 166.780 37.090 170.200 ;
        RECT 36.890 166.460 37.150 166.780 ;
        RECT 37.410 165.420 37.550 172.240 ;
        RECT 37.350 165.100 37.610 165.420 ;
        RECT 37.870 163.720 38.010 179.720 ;
        RECT 38.270 175.980 38.530 176.300 ;
        RECT 38.330 175.620 38.470 175.980 ;
        RECT 38.790 175.620 38.930 191.620 ;
        RECT 38.270 175.300 38.530 175.620 ;
        RECT 38.730 175.300 38.990 175.620 ;
        RECT 38.730 172.240 38.990 172.560 ;
        RECT 38.790 170.860 38.930 172.240 ;
        RECT 38.730 170.540 38.990 170.860 ;
        RECT 39.250 167.460 39.390 194.340 ;
        RECT 39.710 189.560 39.850 196.720 ;
        RECT 40.170 191.600 40.310 196.810 ;
        RECT 41.490 196.720 41.750 196.810 ;
        RECT 42.400 196.525 42.680 196.895 ;
        RECT 42.930 196.700 43.070 199.530 ;
        RECT 43.330 198.760 43.590 199.080 ;
        RECT 42.870 196.380 43.130 196.700 ;
        RECT 40.850 195.505 42.390 195.875 ;
        RECT 42.870 195.020 43.130 195.340 ;
        RECT 42.400 193.125 42.680 193.495 ;
        RECT 42.470 191.600 42.610 193.125 ;
        RECT 40.110 191.280 40.370 191.600 ;
        RECT 42.410 191.280 42.670 191.600 ;
        RECT 39.650 189.240 39.910 189.560 ;
        RECT 40.170 189.220 40.310 191.280 ;
        RECT 42.930 190.920 43.070 195.020 ;
        RECT 43.390 192.280 43.530 198.760 ;
        RECT 43.850 198.060 43.990 199.780 ;
        RECT 43.790 197.740 44.050 198.060 ;
        RECT 43.790 196.380 44.050 196.700 ;
        RECT 43.850 194.320 43.990 196.380 ;
        RECT 43.790 194.000 44.050 194.320 ;
        RECT 43.850 192.620 43.990 194.000 ;
        RECT 43.790 192.300 44.050 192.620 ;
        RECT 43.330 191.960 43.590 192.280 ;
        RECT 42.870 190.600 43.130 190.920 ;
        RECT 40.850 190.065 42.390 190.435 ;
        RECT 42.930 189.810 43.070 190.600 ;
        RECT 42.010 189.670 43.070 189.810 ;
        RECT 40.110 188.900 40.370 189.220 ;
        RECT 42.010 187.375 42.150 189.670 ;
        RECT 42.410 188.900 42.670 189.220 ;
        RECT 41.940 187.005 42.220 187.375 ;
        RECT 39.650 185.840 39.910 186.160 ;
        RECT 39.710 184.460 39.850 185.840 ;
        RECT 42.470 185.820 42.610 188.900 ;
        RECT 43.330 187.880 43.590 188.200 ;
        RECT 42.860 187.005 43.140 187.375 ;
        RECT 42.930 186.500 43.070 187.005 ;
        RECT 42.870 186.180 43.130 186.500 ;
        RECT 40.110 185.500 40.370 185.820 ;
        RECT 42.410 185.500 42.670 185.820 ;
        RECT 39.650 184.140 39.910 184.460 ;
        RECT 39.650 179.720 39.910 180.040 ;
        RECT 39.710 176.300 39.850 179.720 ;
        RECT 39.650 175.980 39.910 176.300 ;
        RECT 39.710 175.135 39.850 175.980 ;
        RECT 39.640 174.765 39.920 175.135 ;
        RECT 39.650 174.280 39.910 174.600 ;
        RECT 39.710 169.840 39.850 174.280 ;
        RECT 39.650 169.520 39.910 169.840 ;
        RECT 38.270 167.140 38.530 167.460 ;
        RECT 39.190 167.140 39.450 167.460 ;
        RECT 39.650 167.140 39.910 167.460 ;
        RECT 38.330 164.400 38.470 167.140 ;
        RECT 39.190 166.120 39.450 166.440 ;
        RECT 38.730 164.935 38.990 165.080 ;
        RECT 38.720 164.565 39.000 164.935 ;
        RECT 38.270 164.080 38.530 164.400 ;
        RECT 37.810 163.400 38.070 163.720 ;
        RECT 37.810 162.380 38.070 162.700 ;
        RECT 37.350 161.360 37.610 161.680 ;
        RECT 36.890 160.680 37.150 161.000 ;
        RECT 36.950 159.495 37.090 160.680 ;
        RECT 36.880 159.125 37.160 159.495 ;
        RECT 36.950 158.960 37.090 159.125 ;
        RECT 36.890 158.640 37.150 158.960 ;
        RECT 35.570 158.050 36.630 158.190 ;
        RECT 35.050 156.490 35.310 156.580 ;
        RECT 35.570 156.490 35.710 158.050 ;
        RECT 35.960 157.085 36.240 157.455 ;
        RECT 35.050 156.350 35.710 156.490 ;
        RECT 35.050 156.260 35.310 156.350 ;
        RECT 35.500 155.725 35.780 156.095 ;
        RECT 35.510 155.580 35.770 155.725 ;
        RECT 35.510 154.220 35.770 154.540 ;
        RECT 34.590 153.200 34.850 153.520 ;
        RECT 33.670 152.520 33.930 152.840 ;
        RECT 33.730 151.140 33.870 152.520 ;
        RECT 33.670 150.820 33.930 151.140 ;
        RECT 34.130 150.820 34.390 151.140 ;
        RECT 32.350 150.400 32.950 150.540 ;
        RECT 33.270 150.400 33.870 150.540 ;
        RECT 30.450 147.760 30.710 148.080 ;
        RECT 30.910 147.760 31.170 148.080 ;
        RECT 31.430 147.310 31.570 150.400 ;
        RECT 32.810 147.820 32.950 150.400 ;
        RECT 33.210 149.800 33.470 150.120 ;
        RECT 33.270 148.760 33.410 149.800 ;
        RECT 33.730 149.100 33.870 150.400 ;
        RECT 33.670 148.780 33.930 149.100 ;
        RECT 33.210 148.440 33.470 148.760 ;
        RECT 33.730 147.935 33.870 148.780 ;
        RECT 32.810 147.680 33.410 147.820 ;
        RECT 30.970 147.170 31.570 147.310 ;
        RECT 30.450 144.360 30.710 144.680 ;
        RECT 29.990 140.620 30.250 140.940 ;
        RECT 30.050 140.260 30.190 140.620 ;
        RECT 30.510 140.455 30.650 144.360 ;
        RECT 29.990 139.940 30.250 140.260 ;
        RECT 30.440 140.085 30.720 140.455 ;
        RECT 30.970 140.260 31.110 147.170 ;
        RECT 32.750 147.080 33.010 147.400 ;
        RECT 32.810 146.380 32.950 147.080 ;
        RECT 32.750 146.060 33.010 146.380 ;
        RECT 31.370 144.360 31.630 144.680 ;
        RECT 31.430 140.940 31.570 144.360 ;
        RECT 31.370 140.620 31.630 140.940 ;
        RECT 30.910 139.940 31.170 140.260 ;
        RECT 30.450 139.260 30.710 139.580 ;
        RECT 29.990 136.880 30.250 137.200 ;
        RECT 30.050 135.160 30.190 136.880 ;
        RECT 29.990 134.840 30.250 135.160 ;
        RECT 29.070 134.500 29.330 134.820 ;
        RECT 18.950 128.720 19.210 129.040 ;
        RECT 28.150 128.720 28.410 129.040 ;
        RECT 16.190 127.020 16.450 127.340 ;
        RECT 18.490 127.020 18.750 127.340 ;
        RECT 19.010 126.660 19.150 128.720 ;
        RECT 21.415 127.505 22.955 127.875 ;
        RECT 29.130 127.340 29.270 134.500 ;
        RECT 30.510 132.100 30.650 139.260 ;
        RECT 30.910 136.540 31.170 136.860 ;
        RECT 30.970 133.800 31.110 136.540 ;
        RECT 32.810 135.160 32.950 146.060 ;
        RECT 33.270 144.535 33.410 147.680 ;
        RECT 33.660 147.565 33.940 147.935 ;
        RECT 34.190 145.780 34.330 150.820 ;
        RECT 33.730 145.640 34.330 145.780 ;
        RECT 33.200 144.165 33.480 144.535 ;
        RECT 32.750 134.840 33.010 135.160 ;
        RECT 33.210 134.160 33.470 134.480 ;
        RECT 30.910 133.480 31.170 133.800 ;
        RECT 30.450 131.780 30.710 132.100 ;
        RECT 29.530 131.440 29.790 131.760 ;
        RECT 29.590 129.720 29.730 131.440 ;
        RECT 30.910 131.100 31.170 131.420 ;
        RECT 30.970 129.720 31.110 131.100 ;
        RECT 29.530 129.400 29.790 129.720 ;
        RECT 30.910 129.400 31.170 129.720 ;
        RECT 33.270 128.360 33.410 134.160 ;
        RECT 33.730 132.780 33.870 145.640 ;
        RECT 34.650 145.360 34.790 153.200 ;
        RECT 35.050 152.860 35.310 153.180 ;
        RECT 35.110 151.820 35.250 152.860 ;
        RECT 35.050 151.500 35.310 151.820 ;
        RECT 35.040 150.965 35.320 151.335 ;
        RECT 35.050 150.820 35.310 150.965 ;
        RECT 35.570 150.540 35.710 154.220 ;
        RECT 36.030 151.220 36.170 157.085 ;
        RECT 37.410 156.580 37.550 161.360 ;
        RECT 37.870 159.640 38.010 162.380 ;
        RECT 37.810 159.320 38.070 159.640 ;
        RECT 37.810 157.960 38.070 158.280 ;
        RECT 36.430 156.260 36.690 156.580 ;
        RECT 37.350 156.260 37.610 156.580 ;
        RECT 36.490 153.375 36.630 156.260 ;
        RECT 37.350 155.240 37.610 155.560 ;
        RECT 36.420 153.005 36.700 153.375 ;
        RECT 37.410 151.730 37.550 155.240 ;
        RECT 37.870 154.540 38.010 157.960 ;
        RECT 38.330 157.260 38.470 164.080 ;
        RECT 38.270 156.940 38.530 157.260 ;
        RECT 38.270 156.260 38.530 156.580 ;
        RECT 37.810 154.220 38.070 154.540 ;
        RECT 38.330 153.520 38.470 156.260 ;
        RECT 38.270 153.200 38.530 153.520 ;
        RECT 38.270 152.520 38.530 152.840 ;
        RECT 36.950 151.590 37.550 151.730 ;
        RECT 36.030 151.080 36.630 151.220 ;
        RECT 35.050 150.140 35.310 150.460 ;
        RECT 35.570 150.400 36.170 150.540 ;
        RECT 35.110 149.100 35.250 150.140 ;
        RECT 35.510 149.800 35.770 150.120 ;
        RECT 35.050 148.780 35.310 149.100 ;
        RECT 35.570 148.420 35.710 149.800 ;
        RECT 35.510 148.100 35.770 148.420 ;
        RECT 36.030 147.820 36.170 150.400 ;
        RECT 36.490 148.420 36.630 151.080 ;
        RECT 36.950 150.800 37.090 151.590 ;
        RECT 37.810 151.500 38.070 151.820 ;
        RECT 36.890 150.480 37.150 150.800 ;
        RECT 37.350 150.480 37.610 150.800 ;
        RECT 36.890 149.800 37.150 150.120 ;
        RECT 36.430 148.100 36.690 148.420 ;
        RECT 35.570 147.680 36.170 147.820 ;
        RECT 34.130 145.040 34.390 145.360 ;
        RECT 34.590 145.040 34.850 145.360 ;
        RECT 34.190 138.220 34.330 145.040 ;
        RECT 34.650 142.980 34.790 145.040 ;
        RECT 34.590 142.660 34.850 142.980 ;
        RECT 34.580 140.765 34.860 141.135 ;
        RECT 34.590 140.620 34.850 140.765 ;
        RECT 35.050 139.940 35.310 140.260 ;
        RECT 34.130 137.900 34.390 138.220 ;
        RECT 35.110 134.480 35.250 139.940 ;
        RECT 35.050 134.160 35.310 134.480 ;
        RECT 35.050 133.480 35.310 133.800 ;
        RECT 33.670 132.460 33.930 132.780 ;
        RECT 33.210 128.040 33.470 128.360 ;
        RECT 29.070 127.020 29.330 127.340 ;
        RECT 33.730 126.660 33.870 132.460 ;
        RECT 34.130 129.740 34.390 130.060 ;
        RECT 34.190 127.340 34.330 129.740 ;
        RECT 35.110 129.720 35.250 133.480 ;
        RECT 35.570 131.760 35.710 147.680 ;
        RECT 35.970 147.080 36.230 147.400 ;
        RECT 36.490 147.255 36.630 148.100 ;
        RECT 36.030 142.640 36.170 147.080 ;
        RECT 36.420 146.885 36.700 147.255 ;
        RECT 36.430 146.060 36.690 146.380 ;
        RECT 36.490 143.660 36.630 146.060 ;
        RECT 36.430 143.340 36.690 143.660 ;
        RECT 35.970 142.320 36.230 142.640 ;
        RECT 36.030 136.860 36.170 142.320 ;
        RECT 36.950 140.940 37.090 149.800 ;
        RECT 37.410 147.740 37.550 150.480 ;
        RECT 37.870 148.080 38.010 151.500 ;
        RECT 38.330 151.480 38.470 152.520 ;
        RECT 38.270 151.160 38.530 151.480 ;
        RECT 37.810 147.760 38.070 148.080 ;
        RECT 37.350 147.420 37.610 147.740 ;
        RECT 37.410 146.380 37.550 147.420 ;
        RECT 38.330 147.400 38.470 151.160 ;
        RECT 37.810 147.080 38.070 147.400 ;
        RECT 38.270 147.080 38.530 147.400 ;
        RECT 37.870 146.380 38.010 147.080 ;
        RECT 37.350 146.060 37.610 146.380 ;
        RECT 37.810 146.060 38.070 146.380 ;
        RECT 38.790 145.780 38.930 164.565 ;
        RECT 39.250 148.760 39.390 166.120 ;
        RECT 39.710 161.680 39.850 167.140 ;
        RECT 40.170 164.060 40.310 185.500 ;
        RECT 40.850 184.625 42.390 184.995 ;
        RECT 41.950 183.460 42.210 183.780 ;
        RECT 42.410 183.460 42.670 183.780 ;
        RECT 41.490 183.120 41.750 183.440 ;
        RECT 41.550 181.400 41.690 183.120 ;
        RECT 41.490 181.080 41.750 181.400 ;
        RECT 42.010 179.950 42.150 183.460 ;
        RECT 42.470 182.760 42.610 183.460 ;
        RECT 42.930 183.180 43.070 186.180 ;
        RECT 43.390 184.460 43.530 187.880 ;
        RECT 43.850 186.160 43.990 192.300 ;
        RECT 44.310 187.180 44.450 212.700 ;
        RECT 45.230 211.660 45.370 212.700 ;
        RECT 45.170 211.340 45.430 211.660 ;
        RECT 44.710 210.320 44.970 210.640 ;
        RECT 44.770 198.060 44.910 210.320 ;
        RECT 45.170 208.620 45.430 208.940 ;
        RECT 45.230 207.580 45.370 208.620 ;
        RECT 45.170 207.260 45.430 207.580 ;
        RECT 45.170 204.880 45.430 205.200 ;
        RECT 45.690 205.055 45.830 217.800 ;
        RECT 47.010 216.780 47.270 217.100 ;
        RECT 47.070 213.360 47.210 216.780 ;
        RECT 48.450 216.080 48.590 218.480 ;
        RECT 48.390 215.760 48.650 216.080 ;
        RECT 48.910 215.740 49.050 218.820 ;
        RECT 49.770 215.760 50.030 216.080 ;
        RECT 48.850 215.420 49.110 215.740 ;
        RECT 49.830 213.700 49.970 215.760 ;
        RECT 49.770 213.380 50.030 213.700 ;
        RECT 47.010 213.040 47.270 213.360 ;
        RECT 50.750 212.680 50.890 220.860 ;
        RECT 51.670 216.420 51.810 220.860 ;
        RECT 60.285 219.985 61.825 220.355 ;
        RECT 62.710 219.820 62.850 221.005 ;
        RECT 62.650 219.500 62.910 219.820 ;
        RECT 66.780 219.645 67.060 220.015 ;
        RECT 61.730 219.160 61.990 219.480 ;
        RECT 52.530 218.480 52.790 218.800 ;
        RECT 51.610 216.100 51.870 216.420 ;
        RECT 52.060 216.245 52.340 216.615 ;
        RECT 51.670 215.255 51.810 216.100 ;
        RECT 51.600 214.885 51.880 215.255 ;
        RECT 50.690 212.360 50.950 212.680 ;
        RECT 50.230 210.660 50.490 210.980 ;
        RECT 47.470 209.980 47.730 210.300 ;
        RECT 47.530 208.455 47.670 209.980 ;
        RECT 50.290 208.940 50.430 210.660 ;
        RECT 50.750 209.815 50.890 212.360 ;
        RECT 52.130 211.660 52.270 216.245 ;
        RECT 52.590 214.380 52.730 218.480 ;
        RECT 61.790 218.460 61.930 219.160 ;
        RECT 65.870 218.820 66.130 219.140 ;
        RECT 56.210 218.140 56.470 218.460 ;
        RECT 56.670 218.140 56.930 218.460 ;
        RECT 58.510 218.140 58.770 218.460 ;
        RECT 61.730 218.140 61.990 218.460 ;
        RECT 64.950 218.140 65.210 218.460 ;
        RECT 56.270 216.420 56.410 218.140 ;
        RECT 52.990 216.100 53.250 216.420 ;
        RECT 53.910 216.100 54.170 216.420 ;
        RECT 56.210 216.100 56.470 216.420 ;
        RECT 52.530 214.060 52.790 214.380 ;
        RECT 53.050 212.680 53.190 216.100 ;
        RECT 53.970 215.400 54.110 216.100 ;
        RECT 54.430 215.740 55.490 215.820 ;
        RECT 54.370 215.680 55.490 215.740 ;
        RECT 54.370 215.420 54.630 215.680 ;
        RECT 53.910 215.080 54.170 215.400 ;
        RECT 54.830 215.080 55.090 215.400 ;
        RECT 53.910 213.380 54.170 213.700 ;
        RECT 52.990 212.360 53.250 212.680 ;
        RECT 52.070 211.340 52.330 211.660 ;
        RECT 53.970 211.175 54.110 213.380 ;
        RECT 53.900 210.805 54.180 211.175 ;
        RECT 54.890 210.980 55.030 215.080 ;
        RECT 54.830 210.660 55.090 210.980 ;
        RECT 51.150 209.980 51.410 210.300 ;
        RECT 50.680 209.445 50.960 209.815 ;
        RECT 51.210 208.940 51.350 209.980 ;
        RECT 55.350 209.960 55.490 215.680 ;
        RECT 55.750 210.660 56.010 210.980 ;
        RECT 52.990 209.640 53.250 209.960 ;
        RECT 54.830 209.640 55.090 209.960 ;
        RECT 55.290 209.640 55.550 209.960 ;
        RECT 50.230 208.620 50.490 208.940 ;
        RECT 51.150 208.620 51.410 208.940 ;
        RECT 47.460 208.085 47.740 208.455 ;
        RECT 49.770 207.940 50.030 208.260 ;
        RECT 50.220 208.085 50.500 208.455 ;
        RECT 49.310 207.260 49.570 207.580 ;
        RECT 49.370 206.220 49.510 207.260 ;
        RECT 48.850 205.900 49.110 206.220 ;
        RECT 49.310 205.900 49.570 206.220 ;
        RECT 45.230 203.015 45.370 204.880 ;
        RECT 45.620 204.685 45.900 205.055 ;
        RECT 45.630 204.200 45.890 204.520 ;
        RECT 45.160 202.645 45.440 203.015 ;
        RECT 45.170 200.460 45.430 200.780 ;
        RECT 44.710 197.740 44.970 198.060 ;
        RECT 44.710 194.000 44.970 194.320 ;
        RECT 44.770 190.920 44.910 194.000 ;
        RECT 44.710 190.600 44.970 190.920 ;
        RECT 44.250 186.860 44.510 187.180 ;
        RECT 44.770 186.580 44.910 190.600 ;
        RECT 44.310 186.440 44.910 186.580 ;
        RECT 43.790 185.840 44.050 186.160 ;
        RECT 43.330 184.140 43.590 184.460 ;
        RECT 43.390 183.690 43.530 184.140 ;
        RECT 43.390 183.550 43.990 183.690 ;
        RECT 42.930 183.040 43.530 183.180 ;
        RECT 42.410 182.440 42.670 182.760 ;
        RECT 42.860 180.885 43.140 181.255 ;
        RECT 42.930 180.720 43.070 180.885 ;
        RECT 42.870 180.400 43.130 180.720 ;
        RECT 42.010 179.810 43.070 179.950 ;
        RECT 40.850 179.185 42.390 179.555 ;
        RECT 41.950 178.700 42.210 179.020 ;
        RECT 42.930 178.930 43.070 179.810 ;
        RECT 42.470 178.790 43.070 178.930 ;
        RECT 42.010 177.855 42.150 178.700 ;
        RECT 41.940 177.485 42.220 177.855 ;
        RECT 42.470 177.320 42.610 178.790 ;
        RECT 42.870 178.020 43.130 178.340 ;
        RECT 42.930 177.320 43.070 178.020 ;
        RECT 43.390 177.660 43.530 183.040 ;
        RECT 43.850 178.680 43.990 183.550 ;
        RECT 43.790 178.360 44.050 178.680 ;
        RECT 43.330 177.340 43.590 177.660 ;
        RECT 40.560 176.805 40.840 177.175 ;
        RECT 41.490 177.000 41.750 177.320 ;
        RECT 42.410 177.000 42.670 177.320 ;
        RECT 42.870 177.000 43.130 177.320 ;
        RECT 40.630 175.620 40.770 176.805 ;
        RECT 40.570 175.300 40.830 175.620 ;
        RECT 41.550 174.940 41.690 177.000 ;
        RECT 42.470 176.380 42.610 177.000 ;
        RECT 42.470 176.240 43.530 176.380 ;
        RECT 41.490 174.620 41.750 174.940 ;
        RECT 40.850 173.745 42.390 174.115 ;
        RECT 42.410 172.920 42.670 173.240 ;
        RECT 42.470 169.070 42.610 172.920 ;
        RECT 42.470 168.930 43.070 169.070 ;
        RECT 40.850 168.305 42.390 168.675 ;
        RECT 42.930 167.540 43.070 168.930 ;
        RECT 43.390 168.900 43.530 176.240 ;
        RECT 44.310 175.280 44.450 186.440 ;
        RECT 44.710 186.015 44.970 186.160 ;
        RECT 44.700 185.645 44.980 186.015 ;
        RECT 45.230 185.480 45.370 200.460 ;
        RECT 45.690 197.040 45.830 204.200 ;
        RECT 48.390 201.480 48.650 201.800 ;
        RECT 47.010 200.350 47.270 200.440 ;
        RECT 46.610 200.210 47.270 200.350 ;
        RECT 46.090 199.780 46.350 200.100 ;
        RECT 46.150 198.255 46.290 199.780 ;
        RECT 46.080 197.885 46.360 198.255 ;
        RECT 45.630 196.720 45.890 197.040 ;
        RECT 45.630 193.320 45.890 193.640 ;
        RECT 45.690 189.220 45.830 193.320 ;
        RECT 45.630 188.900 45.890 189.220 ;
        RECT 45.630 186.520 45.890 186.840 ;
        RECT 45.170 185.160 45.430 185.480 ;
        RECT 45.170 183.460 45.430 183.780 ;
        RECT 44.710 180.740 44.970 181.060 ;
        RECT 44.250 174.960 44.510 175.280 ;
        RECT 43.790 174.280 44.050 174.600 ;
        RECT 43.850 173.580 43.990 174.280 ;
        RECT 43.790 173.260 44.050 173.580 ;
        RECT 43.850 169.500 43.990 173.260 ;
        RECT 44.250 169.520 44.510 169.840 ;
        RECT 43.790 169.180 44.050 169.500 ;
        RECT 43.390 168.760 43.990 168.900 ;
        RECT 42.930 167.400 43.530 167.540 ;
        RECT 42.870 166.460 43.130 166.780 ;
        RECT 40.110 163.740 40.370 164.060 ;
        RECT 40.170 162.270 40.310 163.740 ;
        RECT 40.850 162.865 42.390 163.235 ;
        RECT 41.490 162.380 41.750 162.700 ;
        RECT 41.030 162.270 41.290 162.360 ;
        RECT 40.170 162.215 41.290 162.270 ;
        RECT 40.170 162.130 41.300 162.215 ;
        RECT 41.020 161.845 41.300 162.130 ;
        RECT 39.650 161.360 39.910 161.680 ;
        RECT 41.550 161.535 41.690 162.380 ;
        RECT 41.480 161.165 41.760 161.535 ;
        RECT 40.110 159.660 40.370 159.980 ;
        RECT 39.650 158.980 39.910 159.300 ;
        RECT 39.710 155.415 39.850 158.980 ;
        RECT 40.170 158.280 40.310 159.660 ;
        RECT 41.550 158.960 41.690 161.165 ;
        RECT 41.490 158.640 41.750 158.960 ;
        RECT 40.110 157.960 40.370 158.280 ;
        RECT 40.170 157.455 40.310 157.960 ;
        RECT 40.100 157.085 40.380 157.455 ;
        RECT 40.850 157.425 42.390 157.795 ;
        RECT 42.410 156.940 42.670 157.260 ;
        RECT 42.470 156.095 42.610 156.940 ;
        RECT 42.930 156.920 43.070 166.460 ;
        RECT 43.390 164.935 43.530 167.400 ;
        RECT 43.320 164.565 43.600 164.935 ;
        RECT 43.390 162.020 43.530 164.565 ;
        RECT 43.850 164.400 43.990 168.760 ;
        RECT 43.790 164.080 44.050 164.400 ;
        RECT 43.790 163.400 44.050 163.720 ;
        RECT 43.330 161.700 43.590 162.020 ;
        RECT 43.850 161.680 43.990 163.400 ;
        RECT 43.790 161.360 44.050 161.680 ;
        RECT 43.330 157.960 43.590 158.280 ;
        RECT 42.870 156.600 43.130 156.920 ;
        RECT 40.110 155.580 40.370 155.900 ;
        RECT 40.560 155.725 40.840 156.095 ;
        RECT 42.400 155.725 42.680 156.095 ;
        RECT 40.570 155.580 40.830 155.725 ;
        RECT 39.640 155.045 39.920 155.415 ;
        RECT 39.640 154.365 39.920 154.735 ;
        RECT 40.170 154.540 40.310 155.580 ;
        RECT 41.950 155.240 42.210 155.560 ;
        RECT 42.010 154.540 42.150 155.240 ;
        RECT 39.710 150.460 39.850 154.365 ;
        RECT 40.110 154.220 40.370 154.540 ;
        RECT 41.950 154.220 42.210 154.540 ;
        RECT 40.170 151.140 40.310 154.220 ;
        RECT 41.940 153.685 42.220 154.055 ;
        RECT 41.950 153.540 42.210 153.685 ;
        RECT 41.940 153.005 42.220 153.375 ;
        RECT 41.950 152.860 42.210 153.005 ;
        RECT 42.470 152.840 42.610 155.725 ;
        RECT 42.870 155.580 43.130 155.900 ;
        RECT 42.410 152.520 42.670 152.840 ;
        RECT 40.850 151.985 42.390 152.355 ;
        RECT 41.490 151.160 41.750 151.480 ;
        RECT 42.930 151.335 43.070 155.580 ;
        RECT 43.390 153.860 43.530 157.960 ;
        RECT 43.850 155.900 43.990 161.360 ;
        RECT 44.310 159.640 44.450 169.520 ;
        RECT 44.770 167.460 44.910 180.740 ;
        RECT 45.230 178.340 45.370 183.460 ;
        RECT 45.690 182.760 45.830 186.520 ;
        RECT 46.150 184.460 46.290 197.885 ;
        RECT 46.610 196.215 46.750 200.210 ;
        RECT 47.010 200.120 47.270 200.210 ;
        RECT 47.930 199.780 48.190 200.100 ;
        RECT 47.470 199.100 47.730 199.420 ;
        RECT 47.010 196.720 47.270 197.040 ;
        RECT 46.540 195.845 46.820 196.215 ;
        RECT 47.070 195.535 47.210 196.720 ;
        RECT 47.000 195.165 47.280 195.535 ;
        RECT 46.550 194.000 46.810 194.320 ;
        RECT 46.610 192.620 46.750 194.000 ;
        RECT 47.010 193.320 47.270 193.640 ;
        RECT 47.070 192.620 47.210 193.320 ;
        RECT 46.550 192.300 46.810 192.620 ;
        RECT 47.010 192.300 47.270 192.620 ;
        RECT 46.550 191.280 46.810 191.600 ;
        RECT 46.610 189.900 46.750 191.280 ;
        RECT 47.010 190.940 47.270 191.260 ;
        RECT 47.070 189.900 47.210 190.940 ;
        RECT 47.530 189.900 47.670 199.100 ;
        RECT 47.990 195.340 48.130 199.780 ;
        RECT 48.450 198.060 48.590 201.480 ;
        RECT 48.910 200.350 49.050 205.900 ;
        RECT 49.830 205.200 49.970 207.940 ;
        RECT 49.770 204.880 50.030 205.200 ;
        RECT 49.830 203.015 49.970 204.880 ;
        RECT 49.760 202.645 50.040 203.015 ;
        RECT 49.770 202.390 50.030 202.480 ;
        RECT 50.290 202.390 50.430 208.085 ;
        RECT 53.050 207.920 53.190 209.640 ;
        RECT 53.450 208.620 53.710 208.940 ;
        RECT 52.990 207.600 53.250 207.920 ;
        RECT 53.510 207.775 53.650 208.620 ;
        RECT 54.890 207.920 55.030 209.640 ;
        RECT 50.690 205.560 50.950 205.880 ;
        RECT 49.770 202.250 50.430 202.390 ;
        RECT 49.770 202.160 50.030 202.250 ;
        RECT 50.750 200.975 50.890 205.560 ;
        RECT 51.610 205.220 51.870 205.540 ;
        RECT 51.670 203.160 51.810 205.220 ;
        RECT 53.050 205.110 53.190 207.600 ;
        RECT 53.440 207.405 53.720 207.775 ;
        RECT 54.830 207.600 55.090 207.920 ;
        RECT 55.350 205.540 55.490 209.640 ;
        RECT 55.810 209.135 55.950 210.660 ;
        RECT 55.740 208.765 56.020 209.135 ;
        RECT 56.270 208.040 56.410 216.100 ;
        RECT 55.810 207.900 56.410 208.040 ;
        RECT 55.810 206.415 55.950 207.900 ;
        RECT 56.210 206.920 56.470 207.240 ;
        RECT 55.740 206.045 56.020 206.415 ;
        RECT 56.270 206.220 56.410 206.920 ;
        RECT 56.210 205.900 56.470 206.220 ;
        RECT 55.290 205.220 55.550 205.540 ;
        RECT 53.450 205.110 53.710 205.200 ;
        RECT 53.050 204.970 53.710 205.110 ;
        RECT 53.450 204.880 53.710 204.970 ;
        RECT 52.530 203.180 52.790 203.500 ;
        RECT 51.610 202.840 51.870 203.160 ;
        RECT 51.670 202.480 51.810 202.840 ;
        RECT 51.610 202.160 51.870 202.480 ;
        RECT 49.770 200.460 50.030 200.780 ;
        RECT 50.680 200.605 50.960 200.975 ;
        RECT 49.310 200.350 49.570 200.440 ;
        RECT 48.910 200.210 49.570 200.350 ;
        RECT 49.310 200.120 49.570 200.210 ;
        RECT 49.830 199.500 49.970 200.460 ;
        RECT 50.680 199.925 50.960 200.295 ;
        RECT 50.690 199.780 50.950 199.925 ;
        RECT 48.910 199.360 49.970 199.500 ;
        RECT 48.390 197.740 48.650 198.060 ;
        RECT 48.910 197.380 49.050 199.360 ;
        RECT 50.750 198.060 50.890 199.780 ;
        RECT 51.150 199.100 51.410 199.420 ;
        RECT 50.690 197.740 50.950 198.060 ;
        RECT 51.210 197.720 51.350 199.100 ;
        RECT 49.310 197.400 49.570 197.720 ;
        RECT 51.150 197.400 51.410 197.720 ;
        RECT 48.850 197.060 49.110 197.380 ;
        RECT 49.370 196.780 49.510 197.400 ;
        RECT 51.670 197.040 51.810 202.160 ;
        RECT 52.070 201.480 52.330 201.800 ;
        RECT 52.130 200.780 52.270 201.480 ;
        RECT 52.070 200.460 52.330 200.780 ;
        RECT 52.590 200.100 52.730 203.180 ;
        RECT 53.510 202.480 53.650 204.880 ;
        RECT 54.830 204.540 55.090 204.860 ;
        RECT 55.280 204.685 55.560 205.055 ;
        RECT 55.290 204.540 55.550 204.685 ;
        RECT 54.890 203.500 55.030 204.540 ;
        RECT 54.830 203.180 55.090 203.500 ;
        RECT 55.290 203.180 55.550 203.500 ;
        RECT 53.450 202.160 53.710 202.480 ;
        RECT 52.990 201.480 53.250 201.800 ;
        RECT 53.050 200.780 53.190 201.480 ;
        RECT 52.990 200.460 53.250 200.780 ;
        RECT 52.530 199.780 52.790 200.100 ;
        RECT 52.990 199.780 53.250 200.100 ;
        RECT 52.520 198.140 52.800 198.255 ;
        RECT 53.050 198.140 53.190 199.780 ;
        RECT 53.510 199.420 53.650 202.160 ;
        RECT 54.360 201.285 54.640 201.655 ;
        RECT 54.830 201.480 55.090 201.800 ;
        RECT 53.910 199.780 54.170 200.100 ;
        RECT 53.450 199.100 53.710 199.420 ;
        RECT 52.070 197.740 52.330 198.060 ;
        RECT 52.520 198.000 53.190 198.140 ;
        RECT 52.520 197.885 52.800 198.000 ;
        RECT 49.770 196.780 50.030 197.040 ;
        RECT 49.370 196.720 50.030 196.780 ;
        RECT 50.690 196.720 50.950 197.040 ;
        RECT 51.150 196.720 51.410 197.040 ;
        RECT 51.610 196.720 51.870 197.040 ;
        RECT 48.850 196.380 49.110 196.700 ;
        RECT 49.370 196.640 49.970 196.720 ;
        RECT 48.910 195.340 49.050 196.380 ;
        RECT 47.930 195.020 48.190 195.340 ;
        RECT 48.850 195.020 49.110 195.340 ;
        RECT 48.910 194.320 49.050 195.020 ;
        RECT 48.390 194.000 48.650 194.320 ;
        RECT 48.850 194.000 49.110 194.320 ;
        RECT 48.450 192.620 48.590 194.000 ;
        RECT 48.390 192.300 48.650 192.620 ;
        RECT 47.930 191.510 48.190 191.600 ;
        RECT 47.930 191.370 48.590 191.510 ;
        RECT 47.930 191.280 48.190 191.370 ;
        RECT 46.550 189.580 46.810 189.900 ;
        RECT 47.010 189.580 47.270 189.900 ;
        RECT 47.470 189.580 47.730 189.900 ;
        RECT 47.930 189.580 48.190 189.900 ;
        RECT 47.990 189.300 48.130 189.580 ;
        RECT 48.450 189.415 48.590 191.370 ;
        RECT 46.610 189.160 48.130 189.300 ;
        RECT 46.610 188.540 46.750 189.160 ;
        RECT 46.550 188.220 46.810 188.540 ;
        RECT 47.010 188.220 47.270 188.540 ;
        RECT 46.540 187.005 46.820 187.375 ;
        RECT 46.610 186.160 46.750 187.005 ;
        RECT 46.550 185.840 46.810 186.160 ;
        RECT 46.550 185.160 46.810 185.480 ;
        RECT 46.610 184.460 46.750 185.160 ;
        RECT 46.090 184.140 46.350 184.460 ;
        RECT 46.550 184.140 46.810 184.460 ;
        RECT 46.150 182.760 46.290 184.140 ;
        RECT 47.070 183.100 47.210 188.220 ;
        RECT 47.530 186.580 47.670 189.160 ;
        RECT 48.380 189.045 48.660 189.415 ;
        RECT 48.910 188.880 49.050 194.000 ;
        RECT 49.370 192.620 49.510 196.640 ;
        RECT 50.230 195.250 50.490 195.340 ;
        RECT 50.750 195.250 50.890 196.720 ;
        RECT 50.230 195.110 50.890 195.250 ;
        RECT 50.230 195.020 50.490 195.110 ;
        RECT 49.770 194.570 50.030 194.660 ;
        RECT 49.770 194.430 50.890 194.570 ;
        RECT 49.770 194.340 50.030 194.430 ;
        RECT 49.310 192.300 49.570 192.620 ;
        RECT 48.850 188.560 49.110 188.880 ;
        RECT 47.530 186.500 48.130 186.580 ;
        RECT 47.530 186.440 48.190 186.500 ;
        RECT 47.930 186.180 48.190 186.440 ;
        RECT 48.910 186.160 49.050 188.560 ;
        RECT 49.370 188.540 49.510 192.300 ;
        RECT 49.770 190.940 50.030 191.260 ;
        RECT 49.830 189.560 49.970 190.940 ;
        RECT 49.770 189.240 50.030 189.560 ;
        RECT 49.310 188.220 49.570 188.540 ;
        RECT 49.760 188.365 50.040 188.735 ;
        RECT 49.370 186.160 49.510 188.220 ;
        RECT 49.830 186.500 49.970 188.365 ;
        RECT 49.770 186.180 50.030 186.500 ;
        RECT 47.470 185.840 47.730 186.160 ;
        RECT 48.850 185.840 49.110 186.160 ;
        RECT 49.310 185.840 49.570 186.160 ;
        RECT 50.230 185.840 50.490 186.160 ;
        RECT 47.530 184.460 47.670 185.840 ;
        RECT 48.840 184.965 49.120 185.335 ;
        RECT 47.470 184.140 47.730 184.460 ;
        RECT 47.930 183.800 48.190 184.120 ;
        RECT 47.010 182.780 47.270 183.100 ;
        RECT 45.630 182.440 45.890 182.760 ;
        RECT 46.090 182.440 46.350 182.760 ;
        RECT 45.690 180.720 45.830 182.440 ;
        RECT 47.070 180.720 47.210 182.780 ;
        RECT 47.470 181.080 47.730 181.400 ;
        RECT 47.530 180.720 47.670 181.080 ;
        RECT 47.990 180.720 48.130 183.800 ;
        RECT 48.910 183.440 49.050 184.965 ;
        RECT 49.370 183.860 49.510 185.840 ;
        RECT 50.290 184.460 50.430 185.840 ;
        RECT 50.230 184.140 50.490 184.460 ;
        RECT 49.370 183.720 49.970 183.860 ;
        RECT 48.850 183.120 49.110 183.440 ;
        RECT 49.310 183.120 49.570 183.440 ;
        RECT 49.830 183.295 49.970 183.720 ;
        RECT 50.230 183.460 50.490 183.780 ;
        RECT 48.390 182.440 48.650 182.760 ;
        RECT 48.450 181.060 48.590 182.440 ;
        RECT 49.370 181.400 49.510 183.120 ;
        RECT 49.760 182.925 50.040 183.295 ;
        RECT 49.310 181.080 49.570 181.400 ;
        RECT 48.390 180.740 48.650 181.060 ;
        RECT 45.630 180.630 45.890 180.720 ;
        RECT 45.630 180.490 46.290 180.630 ;
        RECT 45.630 180.400 45.890 180.490 ;
        RECT 45.630 179.720 45.890 180.040 ;
        RECT 45.690 178.680 45.830 179.720 ;
        RECT 45.630 178.360 45.890 178.680 ;
        RECT 45.170 178.020 45.430 178.340 ;
        RECT 46.150 177.660 46.290 180.490 ;
        RECT 47.010 180.400 47.270 180.720 ;
        RECT 47.470 180.400 47.730 180.720 ;
        RECT 47.930 180.400 48.190 180.720 ;
        RECT 45.170 177.340 45.430 177.660 ;
        RECT 46.090 177.340 46.350 177.660 ;
        RECT 45.230 174.600 45.370 177.340 ;
        RECT 46.090 175.980 46.350 176.300 ;
        RECT 45.630 175.300 45.890 175.620 ;
        RECT 45.170 174.280 45.430 174.600 ;
        RECT 45.690 173.240 45.830 175.300 ;
        RECT 45.630 172.920 45.890 173.240 ;
        RECT 45.620 172.045 45.900 172.415 ;
        RECT 45.690 170.860 45.830 172.045 ;
        RECT 45.630 170.540 45.890 170.860 ;
        RECT 45.170 169.860 45.430 170.180 ;
        RECT 45.230 169.695 45.370 169.860 ;
        RECT 45.160 169.325 45.440 169.695 ;
        RECT 46.150 169.160 46.290 175.980 ;
        RECT 46.550 174.280 46.810 174.600 ;
        RECT 46.610 172.900 46.750 174.280 ;
        RECT 47.070 173.580 47.210 180.400 ;
        RECT 47.470 178.360 47.730 178.680 ;
        RECT 47.530 176.300 47.670 178.360 ;
        RECT 47.930 178.250 48.190 178.340 ;
        RECT 48.450 178.250 48.590 180.740 ;
        RECT 49.770 180.575 50.030 180.720 ;
        RECT 49.760 180.205 50.040 180.575 ;
        RECT 49.760 179.525 50.040 179.895 ;
        RECT 48.850 178.930 49.110 179.020 ;
        RECT 48.850 178.790 49.510 178.930 ;
        RECT 48.850 178.700 49.110 178.790 ;
        RECT 47.930 178.110 48.590 178.250 ;
        RECT 47.930 178.020 48.190 178.110 ;
        RECT 47.470 175.980 47.730 176.300 ;
        RECT 47.990 175.960 48.130 178.020 ;
        RECT 47.930 175.640 48.190 175.960 ;
        RECT 47.470 174.960 47.730 175.280 ;
        RECT 47.010 173.260 47.270 173.580 ;
        RECT 46.550 172.580 46.810 172.900 ;
        RECT 47.010 172.580 47.270 172.900 ;
        RECT 46.610 169.840 46.750 172.580 ;
        RECT 46.550 169.520 46.810 169.840 ;
        RECT 45.170 168.840 45.430 169.160 ;
        RECT 46.090 168.840 46.350 169.160 ;
        RECT 44.710 167.140 44.970 167.460 ;
        RECT 44.710 166.460 44.970 166.780 ;
        RECT 44.770 166.295 44.910 166.460 ;
        RECT 44.700 165.925 44.980 166.295 ;
        RECT 44.710 164.080 44.970 164.400 ;
        RECT 44.770 159.980 44.910 164.080 ;
        RECT 45.230 162.700 45.370 168.840 ;
        RECT 47.070 168.050 47.210 172.580 ;
        RECT 47.530 170.860 47.670 174.960 ;
        RECT 47.990 173.240 48.130 175.640 ;
        RECT 49.370 174.510 49.510 178.790 ;
        RECT 49.830 175.135 49.970 179.525 ;
        RECT 50.290 178.340 50.430 183.460 ;
        RECT 50.750 183.100 50.890 194.430 ;
        RECT 51.210 193.980 51.350 196.720 ;
        RECT 52.130 195.250 52.270 197.740 ;
        RECT 53.050 195.340 53.190 198.000 ;
        RECT 53.970 197.460 54.110 199.780 ;
        RECT 54.430 199.080 54.570 201.285 ;
        RECT 54.890 200.440 55.030 201.480 ;
        RECT 54.830 200.120 55.090 200.440 ;
        RECT 54.370 198.760 54.630 199.080 ;
        RECT 54.890 198.935 55.030 200.120 ;
        RECT 54.820 198.565 55.100 198.935 ;
        RECT 54.360 197.460 54.640 197.575 ;
        RECT 53.450 197.060 53.710 197.380 ;
        RECT 53.970 197.320 54.640 197.460 ;
        RECT 54.890 197.380 55.030 198.565 ;
        RECT 55.350 198.060 55.490 203.180 ;
        RECT 55.740 200.605 56.020 200.975 ;
        RECT 55.290 197.740 55.550 198.060 ;
        RECT 54.360 197.205 54.640 197.320 ;
        RECT 54.830 197.060 55.090 197.380 ;
        RECT 51.670 195.110 52.270 195.250 ;
        RECT 51.670 194.660 51.810 195.110 ;
        RECT 52.990 195.020 53.250 195.340 ;
        RECT 51.610 194.340 51.870 194.660 ;
        RECT 52.070 194.340 52.330 194.660 ;
        RECT 52.530 194.340 52.790 194.660 ;
        RECT 52.980 194.485 53.260 194.855 ;
        RECT 52.990 194.340 53.250 194.485 ;
        RECT 51.150 193.660 51.410 193.980 ;
        RECT 51.150 188.560 51.410 188.880 ;
        RECT 51.210 187.180 51.350 188.560 ;
        RECT 51.150 186.860 51.410 187.180 ;
        RECT 51.670 184.460 51.810 194.340 ;
        RECT 52.130 192.135 52.270 194.340 ;
        RECT 52.590 194.060 52.730 194.340 ;
        RECT 53.510 194.060 53.650 197.060 ;
        RECT 53.910 196.380 54.170 196.700 ;
        RECT 54.830 196.380 55.090 196.700 ;
        RECT 52.590 193.920 53.650 194.060 ;
        RECT 53.440 193.380 53.720 193.495 ;
        RECT 53.970 193.380 54.110 196.380 ;
        RECT 54.890 196.215 55.030 196.380 ;
        RECT 54.820 195.845 55.100 196.215 ;
        RECT 55.290 196.040 55.550 196.360 ;
        RECT 55.350 194.660 55.490 196.040 ;
        RECT 55.290 194.340 55.550 194.660 ;
        RECT 54.830 193.660 55.090 193.980 ;
        RECT 53.440 193.240 54.570 193.380 ;
        RECT 53.440 193.125 53.720 193.240 ;
        RECT 54.430 192.620 54.570 193.240 ;
        RECT 54.370 192.300 54.630 192.620 ;
        RECT 52.060 191.765 52.340 192.135 ;
        RECT 54.370 189.240 54.630 189.560 ;
        RECT 53.910 188.560 54.170 188.880 ;
        RECT 52.530 188.220 52.790 188.540 ;
        RECT 51.610 184.370 51.870 184.460 ;
        RECT 51.610 184.230 52.270 184.370 ;
        RECT 51.610 184.140 51.870 184.230 ;
        RECT 51.610 183.120 51.870 183.440 ;
        RECT 50.690 182.780 50.950 183.100 ;
        RECT 50.750 181.255 50.890 182.780 ;
        RECT 51.150 182.440 51.410 182.760 ;
        RECT 50.680 180.885 50.960 181.255 ;
        RECT 51.210 178.340 51.350 182.440 ;
        RECT 51.670 180.040 51.810 183.120 ;
        RECT 52.130 180.720 52.270 184.230 ;
        RECT 52.070 180.400 52.330 180.720 ;
        RECT 52.590 180.575 52.730 188.220 ;
        RECT 53.450 187.880 53.710 188.200 ;
        RECT 53.510 186.500 53.650 187.880 ;
        RECT 53.450 186.180 53.710 186.500 ;
        RECT 53.970 186.015 54.110 188.560 ;
        RECT 52.990 185.500 53.250 185.820 ;
        RECT 53.900 185.645 54.180 186.015 ;
        RECT 54.430 185.820 54.570 189.240 ;
        RECT 54.890 186.695 55.030 193.660 ;
        RECT 55.350 191.940 55.490 194.340 ;
        RECT 55.290 191.620 55.550 191.940 ;
        RECT 55.810 190.830 55.950 200.605 ;
        RECT 56.200 199.925 56.480 200.295 ;
        RECT 56.270 199.420 56.410 199.925 ;
        RECT 56.210 199.100 56.470 199.420 ;
        RECT 56.210 197.740 56.470 198.060 ;
        RECT 56.270 192.020 56.410 197.740 ;
        RECT 56.730 192.620 56.870 218.140 ;
        RECT 57.130 215.935 57.390 216.080 ;
        RECT 57.120 215.565 57.400 215.935 ;
        RECT 57.590 215.760 57.850 216.080 ;
        RECT 57.650 210.640 57.790 215.760 ;
        RECT 58.050 215.080 58.310 215.400 ;
        RECT 58.110 213.360 58.250 215.080 ;
        RECT 58.050 213.040 58.310 213.360 ;
        RECT 58.050 212.360 58.310 212.680 ;
        RECT 58.110 210.980 58.250 212.360 ;
        RECT 58.050 210.660 58.310 210.980 ;
        RECT 57.130 210.320 57.390 210.640 ;
        RECT 57.590 210.320 57.850 210.640 ;
        RECT 57.190 208.940 57.330 210.320 ;
        RECT 57.130 208.620 57.390 208.940 ;
        RECT 57.130 207.775 57.390 207.920 ;
        RECT 57.120 207.405 57.400 207.775 ;
        RECT 57.650 207.150 57.790 210.320 ;
        RECT 58.050 207.260 58.310 207.580 ;
        RECT 57.190 207.010 57.790 207.150 ;
        RECT 58.110 207.095 58.250 207.260 ;
        RECT 57.190 203.160 57.330 207.010 ;
        RECT 58.040 206.725 58.320 207.095 ;
        RECT 57.580 205.365 57.860 205.735 ;
        RECT 57.130 202.840 57.390 203.160 ;
        RECT 57.130 202.160 57.390 202.480 ;
        RECT 57.190 200.440 57.330 202.160 ;
        RECT 57.130 200.120 57.390 200.440 ;
        RECT 57.650 197.040 57.790 205.365 ;
        RECT 58.050 205.220 58.310 205.540 ;
        RECT 58.110 203.500 58.250 205.220 ;
        RECT 58.050 203.180 58.310 203.500 ;
        RECT 58.050 202.160 58.310 202.480 ;
        RECT 57.590 196.720 57.850 197.040 ;
        RECT 58.110 196.360 58.250 202.160 ;
        RECT 57.130 196.040 57.390 196.360 ;
        RECT 58.050 196.040 58.310 196.360 ;
        RECT 57.190 195.000 57.330 196.040 ;
        RECT 57.130 194.680 57.390 195.000 ;
        RECT 56.670 192.300 56.930 192.620 ;
        RECT 58.110 192.135 58.250 196.040 ;
        RECT 56.270 191.880 56.870 192.020 ;
        RECT 56.210 190.830 56.470 190.920 ;
        RECT 55.810 190.690 56.470 190.830 ;
        RECT 55.290 189.580 55.550 189.900 ;
        RECT 55.350 188.540 55.490 189.580 ;
        RECT 55.810 189.220 55.950 190.690 ;
        RECT 56.210 190.600 56.470 190.690 ;
        RECT 55.750 188.900 56.010 189.220 ;
        RECT 55.290 188.220 55.550 188.540 ;
        RECT 55.280 187.260 55.560 187.375 ;
        RECT 55.810 187.260 55.950 188.900 ;
        RECT 55.280 187.120 55.950 187.260 ;
        RECT 55.280 187.005 55.560 187.120 ;
        RECT 54.820 186.325 55.100 186.695 ;
        RECT 55.290 186.180 55.550 186.500 ;
        RECT 54.370 185.500 54.630 185.820 ;
        RECT 52.520 180.205 52.800 180.575 ;
        RECT 51.610 179.720 51.870 180.040 ;
        RECT 52.070 179.720 52.330 180.040 ;
        RECT 52.530 179.720 52.790 180.040 ;
        RECT 52.130 179.020 52.270 179.720 ;
        RECT 52.070 178.700 52.330 179.020 ;
        RECT 52.590 178.680 52.730 179.720 ;
        RECT 52.530 178.360 52.790 178.680 ;
        RECT 50.230 178.020 50.490 178.340 ;
        RECT 51.150 178.020 51.410 178.340 ;
        RECT 49.760 174.765 50.040 175.135 ;
        RECT 50.290 174.940 50.430 178.020 ;
        RECT 50.690 177.855 50.950 178.000 ;
        RECT 50.680 177.485 50.960 177.855 ;
        RECT 51.150 177.000 51.410 177.320 ;
        RECT 52.530 177.175 52.790 177.320 ;
        RECT 50.230 174.620 50.490 174.940 ;
        RECT 49.770 174.510 50.030 174.600 ;
        RECT 49.370 174.370 50.030 174.510 ;
        RECT 49.770 174.280 50.030 174.370 ;
        RECT 48.390 173.260 48.650 173.580 ;
        RECT 47.930 172.920 48.190 173.240 ;
        RECT 47.470 170.540 47.730 170.860 ;
        RECT 47.990 169.840 48.130 172.920 ;
        RECT 47.930 169.520 48.190 169.840 ;
        RECT 47.470 168.050 47.730 168.140 ;
        RECT 47.070 167.910 47.730 168.050 ;
        RECT 47.470 167.820 47.730 167.910 ;
        RECT 45.630 167.140 45.890 167.460 ;
        RECT 47.930 167.370 48.190 167.460 ;
        RECT 48.450 167.370 48.590 173.260 ;
        RECT 49.830 173.240 49.970 174.280 ;
        RECT 49.770 172.920 50.030 173.240 ;
        RECT 48.850 172.580 49.110 172.900 ;
        RECT 47.930 167.230 48.590 167.370 ;
        RECT 47.930 167.140 48.190 167.230 ;
        RECT 45.690 166.440 45.830 167.140 ;
        RECT 46.090 166.460 46.350 166.780 ;
        RECT 45.630 166.120 45.890 166.440 ;
        RECT 45.630 163.400 45.890 163.720 ;
        RECT 45.170 162.380 45.430 162.700 ;
        RECT 44.710 159.660 44.970 159.980 ;
        RECT 44.250 159.320 44.510 159.640 ;
        RECT 45.170 158.980 45.430 159.300 ;
        RECT 44.240 158.445 44.520 158.815 ;
        RECT 44.250 158.300 44.510 158.445 ;
        RECT 44.710 157.960 44.970 158.280 ;
        RECT 44.770 155.900 44.910 157.960 ;
        RECT 45.230 156.920 45.370 158.980 ;
        RECT 45.170 156.600 45.430 156.920 ;
        RECT 43.790 155.580 44.050 155.900 ;
        RECT 44.710 155.580 44.970 155.900 ;
        RECT 43.330 153.540 43.590 153.860 ;
        RECT 44.240 153.685 44.520 154.055 ;
        RECT 44.310 152.580 44.450 153.685 ;
        RECT 43.850 152.440 44.450 152.580 ;
        RECT 43.850 151.730 43.990 152.440 ;
        RECT 43.390 151.590 43.990 151.730 ;
        RECT 44.250 151.730 44.510 151.820 ;
        RECT 44.770 151.730 44.910 155.580 ;
        RECT 45.170 154.220 45.430 154.540 ;
        RECT 45.230 152.015 45.370 154.220 ;
        RECT 44.250 151.590 44.910 151.730 ;
        RECT 45.160 151.645 45.440 152.015 ;
        RECT 40.110 150.820 40.370 151.140 ;
        RECT 39.650 150.140 39.910 150.460 ;
        RECT 40.100 150.285 40.380 150.655 ;
        RECT 41.020 150.285 41.300 150.655 ;
        RECT 39.190 148.440 39.450 148.760 ;
        RECT 40.170 148.080 40.310 150.285 ;
        RECT 40.570 149.800 40.830 150.120 ;
        RECT 39.650 147.760 39.910 148.080 ;
        RECT 40.110 147.760 40.370 148.080 ;
        RECT 37.410 145.640 38.930 145.780 ;
        RECT 36.890 140.620 37.150 140.940 ;
        RECT 37.410 139.920 37.550 145.640 ;
        RECT 37.810 145.040 38.070 145.360 ;
        RECT 37.870 142.980 38.010 145.040 ;
        RECT 38.730 144.360 38.990 144.680 ;
        RECT 38.790 143.060 38.930 144.360 ;
        RECT 37.810 142.660 38.070 142.980 ;
        RECT 38.330 142.920 38.930 143.060 ;
        RECT 37.350 139.600 37.610 139.920 ;
        RECT 35.970 136.540 36.230 136.860 ;
        RECT 36.030 135.160 36.170 136.540 ;
        RECT 37.410 135.500 37.550 139.600 ;
        RECT 37.870 138.220 38.010 142.660 ;
        RECT 38.330 140.940 38.470 142.920 ;
        RECT 39.180 142.805 39.460 143.175 ;
        RECT 39.250 142.640 39.390 142.805 ;
        RECT 38.730 142.320 38.990 142.640 ;
        RECT 39.190 142.320 39.450 142.640 ;
        RECT 38.790 141.815 38.930 142.320 ;
        RECT 38.720 141.445 39.000 141.815 ;
        RECT 38.270 140.620 38.530 140.940 ;
        RECT 39.710 139.660 39.850 147.760 ;
        RECT 40.630 147.650 40.770 149.800 ;
        RECT 41.090 148.760 41.230 150.285 ;
        RECT 41.030 148.440 41.290 148.760 ;
        RECT 41.550 148.080 41.690 151.160 ;
        RECT 42.410 150.820 42.670 151.140 ;
        RECT 42.860 150.965 43.140 151.335 ;
        RECT 43.390 151.140 43.530 151.590 ;
        RECT 44.250 151.500 44.510 151.590 ;
        RECT 43.330 150.820 43.590 151.140 ;
        RECT 43.790 151.050 44.050 151.140 ;
        RECT 43.790 150.910 44.450 151.050 ;
        RECT 44.700 150.965 44.980 151.335 ;
        RECT 43.790 150.820 44.050 150.910 ;
        RECT 41.490 147.760 41.750 148.080 ;
        RECT 42.470 147.820 42.610 150.820 ;
        RECT 42.870 150.480 43.130 150.800 ;
        RECT 42.930 149.010 43.070 150.480 ;
        RECT 43.320 150.285 43.600 150.655 ;
        RECT 44.310 150.540 44.450 150.910 ;
        RECT 43.850 150.400 44.450 150.540 ;
        RECT 43.330 150.140 43.590 150.285 ;
        RECT 43.850 149.180 43.990 150.400 ;
        RECT 44.770 150.120 44.910 150.965 ;
        RECT 44.710 149.800 44.970 150.120 ;
        RECT 43.850 149.040 44.910 149.180 ;
        RECT 42.930 148.870 43.530 149.010 ;
        RECT 43.390 148.670 43.530 148.870 ;
        RECT 44.250 148.670 44.510 148.760 ;
        RECT 43.390 148.530 44.510 148.670 ;
        RECT 44.250 148.440 44.510 148.530 ;
        RECT 42.470 147.680 43.530 147.820 ;
        RECT 43.790 147.760 44.050 148.080 ;
        RECT 40.625 147.510 40.770 147.650 ;
        RECT 40.625 147.310 40.765 147.510 ;
        RECT 40.350 147.170 40.765 147.310 ;
        RECT 40.350 147.140 40.490 147.170 ;
        RECT 40.170 147.000 40.490 147.140 ;
        RECT 42.870 147.080 43.130 147.400 ;
        RECT 40.170 142.640 40.310 147.000 ;
        RECT 40.850 146.545 42.390 146.915 ;
        RECT 40.570 145.950 40.830 146.040 ;
        RECT 40.570 145.810 41.230 145.950 ;
        RECT 40.570 145.720 40.830 145.810 ;
        RECT 41.090 145.215 41.230 145.810 ;
        RECT 41.020 144.845 41.300 145.215 ;
        RECT 42.400 144.845 42.680 145.215 ;
        RECT 42.470 143.660 42.610 144.845 ;
        RECT 42.930 143.660 43.070 147.080 ;
        RECT 42.410 143.340 42.670 143.660 ;
        RECT 42.870 143.340 43.130 143.660 ;
        RECT 42.870 142.660 43.130 142.980 ;
        RECT 40.110 142.320 40.370 142.640 ;
        RECT 40.110 141.640 40.370 141.960 ;
        RECT 39.250 139.520 39.850 139.660 ;
        RECT 38.730 138.920 38.990 139.240 ;
        RECT 37.810 137.900 38.070 138.220 ;
        RECT 37.350 135.180 37.610 135.500 ;
        RECT 37.810 135.180 38.070 135.500 ;
        RECT 35.970 134.840 36.230 135.160 ;
        RECT 36.030 132.780 36.170 134.840 ;
        RECT 37.410 132.780 37.550 135.180 ;
        RECT 35.970 132.460 36.230 132.780 ;
        RECT 37.350 132.460 37.610 132.780 ;
        RECT 37.870 132.100 38.010 135.180 ;
        RECT 37.810 131.780 38.070 132.100 ;
        RECT 35.510 131.440 35.770 131.760 ;
        RECT 35.050 129.400 35.310 129.720 ;
        RECT 34.130 127.020 34.390 127.340 ;
        RECT 13.890 126.340 14.150 126.660 ;
        RECT 14.350 126.340 14.610 126.660 ;
        RECT 18.950 126.340 19.210 126.660 ;
        RECT 33.670 126.340 33.930 126.660 ;
        RECT 35.570 126.320 35.710 131.440 ;
        RECT 38.790 126.660 38.930 138.920 ;
        RECT 39.250 138.220 39.390 139.520 ;
        RECT 39.650 138.920 39.910 139.240 ;
        RECT 39.190 137.900 39.450 138.220 ;
        RECT 39.190 136.540 39.450 136.860 ;
        RECT 39.250 127.340 39.390 136.540 ;
        RECT 39.190 127.020 39.450 127.340 ;
        RECT 38.730 126.340 38.990 126.660 ;
        RECT 39.710 126.320 39.850 138.920 ;
        RECT 40.170 136.860 40.310 141.640 ;
        RECT 40.850 141.105 42.390 141.475 ;
        RECT 42.930 140.940 43.070 142.660 ;
        RECT 42.870 140.620 43.130 140.940 ;
        RECT 42.870 138.920 43.130 139.240 ;
        RECT 40.110 136.540 40.370 136.860 ;
        RECT 40.170 129.040 40.310 136.540 ;
        RECT 40.850 135.665 42.390 136.035 ;
        RECT 42.930 132.100 43.070 138.920 ;
        RECT 42.870 131.780 43.130 132.100 ;
        RECT 42.870 130.760 43.130 131.080 ;
        RECT 40.850 130.225 42.390 130.595 ;
        RECT 41.950 129.400 42.210 129.720 ;
        RECT 42.410 129.400 42.670 129.720 ;
        RECT 40.110 128.720 40.370 129.040 ;
        RECT 42.010 127.340 42.150 129.400 ;
        RECT 41.950 127.020 42.210 127.340 ;
        RECT 42.470 126.660 42.610 129.400 ;
        RECT 42.930 127.340 43.070 130.760 ;
        RECT 43.390 128.270 43.530 147.680 ;
        RECT 43.850 146.575 43.990 147.760 ;
        RECT 43.780 146.205 44.060 146.575 ;
        RECT 43.850 145.360 43.990 146.205 ;
        RECT 43.790 145.040 44.050 145.360 ;
        RECT 44.310 143.320 44.450 148.440 ;
        RECT 44.250 143.000 44.510 143.320 ;
        RECT 43.790 141.640 44.050 141.960 ;
        RECT 43.850 140.940 43.990 141.640 ;
        RECT 43.790 140.620 44.050 140.940 ;
        RECT 43.850 140.260 43.990 140.620 ;
        RECT 43.790 139.940 44.050 140.260 ;
        RECT 44.250 136.540 44.510 136.860 ;
        RECT 43.790 133.820 44.050 134.140 ;
        RECT 43.850 131.420 43.990 133.820 ;
        RECT 44.310 132.780 44.450 136.540 ;
        RECT 44.770 135.500 44.910 149.040 ;
        RECT 45.170 147.760 45.430 148.080 ;
        RECT 45.230 147.400 45.370 147.760 ;
        RECT 45.170 147.080 45.430 147.400 ;
        RECT 45.690 146.290 45.830 163.400 ;
        RECT 46.150 148.420 46.290 166.460 ;
        RECT 47.990 166.180 48.130 167.140 ;
        RECT 48.380 166.605 48.660 166.975 ;
        RECT 48.390 166.460 48.650 166.605 ;
        RECT 47.990 166.040 48.590 166.180 ;
        RECT 46.550 164.420 46.810 164.740 ;
        RECT 46.610 154.540 46.750 164.420 ;
        RECT 47.930 163.740 48.190 164.060 ;
        RECT 47.470 163.400 47.730 163.720 ;
        RECT 47.010 158.300 47.270 158.620 ;
        RECT 46.550 154.220 46.810 154.540 ;
        RECT 47.070 153.260 47.210 158.300 ;
        RECT 47.530 156.660 47.670 163.400 ;
        RECT 47.990 157.260 48.130 163.740 ;
        RECT 47.930 156.940 48.190 157.260 ;
        RECT 47.530 156.520 48.130 156.660 ;
        RECT 47.470 155.415 47.730 155.560 ;
        RECT 47.460 155.045 47.740 155.415 ;
        RECT 47.990 153.520 48.130 156.520 ;
        RECT 48.450 155.560 48.590 166.040 ;
        RECT 48.910 165.080 49.050 172.580 ;
        RECT 49.830 171.735 49.970 172.920 ;
        RECT 50.290 172.810 50.430 174.620 ;
        RECT 51.210 173.580 51.350 177.000 ;
        RECT 52.520 176.805 52.800 177.175 ;
        RECT 52.070 175.640 52.330 175.960 ;
        RECT 51.610 174.850 51.870 174.940 ;
        RECT 52.130 174.850 52.270 175.640 ;
        RECT 53.050 175.280 53.190 185.500 ;
        RECT 53.910 180.575 54.170 180.720 ;
        RECT 53.900 180.460 54.180 180.575 ;
        RECT 53.510 180.320 54.180 180.460 ;
        RECT 54.430 180.460 54.570 185.500 ;
        RECT 55.350 183.440 55.490 186.180 ;
        RECT 55.750 183.460 56.010 183.780 ;
        RECT 56.210 183.460 56.470 183.780 ;
        RECT 55.290 183.120 55.550 183.440 ;
        RECT 55.810 181.740 55.950 183.460 ;
        RECT 55.750 181.420 56.010 181.740 ;
        RECT 56.270 181.255 56.410 183.460 ;
        RECT 56.200 180.885 56.480 181.255 ;
        RECT 54.430 180.320 55.030 180.460 ;
        RECT 53.510 179.020 53.650 180.320 ;
        RECT 53.900 180.205 54.180 180.320 ;
        RECT 54.890 180.040 55.030 180.320 ;
        RECT 53.910 179.720 54.170 180.040 ;
        RECT 54.830 179.720 55.090 180.040 ;
        RECT 56.210 179.720 56.470 180.040 ;
        RECT 56.730 179.895 56.870 191.880 ;
        RECT 58.040 191.765 58.320 192.135 ;
        RECT 58.570 189.900 58.710 218.140 ;
        RECT 61.270 217.800 61.530 218.120 ;
        RECT 61.330 216.760 61.470 217.800 ;
        RECT 61.270 216.440 61.530 216.760 ;
        RECT 61.720 216.245 62.000 216.615 ;
        RECT 61.730 216.100 61.990 216.245 ;
        RECT 64.030 216.100 64.290 216.420 ;
        RECT 59.890 215.420 60.150 215.740 ;
        RECT 58.960 214.205 59.240 214.575 ;
        RECT 58.970 214.060 59.230 214.205 ;
        RECT 59.950 210.980 60.090 215.420 ;
        RECT 61.960 215.080 62.220 215.400 ;
        RECT 60.285 214.545 61.825 214.915 ;
        RECT 62.020 214.290 62.160 215.080 ;
        RECT 61.330 214.150 62.160 214.290 ;
        RECT 61.330 213.020 61.470 214.150 ;
        RECT 61.270 212.700 61.530 213.020 ;
        RECT 61.330 211.660 61.470 212.700 ;
        RECT 61.270 211.340 61.530 211.660 ;
        RECT 64.090 211.320 64.230 216.100 ;
        RECT 65.010 213.700 65.150 218.140 ;
        RECT 65.930 217.100 66.070 218.820 ;
        RECT 66.330 218.140 66.590 218.460 ;
        RECT 66.390 217.975 66.530 218.140 ;
        RECT 66.850 218.120 66.990 219.645 ;
        RECT 68.230 219.480 68.370 221.800 ;
        RECT 68.620 221.685 68.900 221.800 ;
        RECT 68.620 221.005 68.900 221.375 ;
        RECT 75.990 221.200 76.250 221.520 ;
        RECT 122.910 221.200 123.170 221.520 ;
        RECT 67.700 218.965 67.980 219.335 ;
        RECT 68.170 219.160 68.430 219.480 ;
        RECT 67.770 218.800 67.910 218.965 ;
        RECT 67.710 218.710 67.970 218.800 ;
        RECT 67.310 218.570 67.970 218.710 ;
        RECT 66.320 217.605 66.600 217.975 ;
        RECT 66.790 217.800 67.050 218.120 ;
        RECT 65.410 216.780 65.670 217.100 ;
        RECT 65.870 216.780 66.130 217.100 ;
        RECT 65.470 216.080 65.610 216.780 ;
        RECT 66.330 216.100 66.590 216.420 ;
        RECT 65.410 215.760 65.670 216.080 ;
        RECT 64.950 213.380 65.210 213.700 ;
        RECT 64.490 213.040 64.750 213.360 ;
        RECT 65.870 213.040 66.130 213.360 ;
        RECT 64.030 211.000 64.290 211.320 ;
        RECT 59.890 210.660 60.150 210.980 ;
        RECT 61.270 210.660 61.530 210.980 ;
        RECT 58.970 210.550 59.230 210.640 ;
        RECT 58.970 210.410 59.630 210.550 ;
        RECT 58.970 210.320 59.230 210.410 ;
        RECT 59.490 207.920 59.630 210.410 ;
        RECT 59.430 207.600 59.690 207.920 ;
        RECT 59.430 205.220 59.690 205.540 ;
        RECT 58.970 204.200 59.230 204.520 ;
        RECT 59.030 203.160 59.170 204.200 ;
        RECT 58.970 202.840 59.230 203.160 ;
        RECT 58.970 202.160 59.230 202.480 ;
        RECT 59.030 201.655 59.170 202.160 ;
        RECT 58.960 201.285 59.240 201.655 ;
        RECT 58.970 199.780 59.230 200.100 ;
        RECT 59.030 197.720 59.170 199.780 ;
        RECT 58.970 197.400 59.230 197.720 ;
        RECT 58.970 196.720 59.230 197.040 ;
        RECT 59.030 194.855 59.170 196.720 ;
        RECT 59.490 195.000 59.630 205.220 ;
        RECT 59.950 201.800 60.090 210.660 ;
        RECT 61.330 210.380 61.470 210.660 ;
        RECT 61.330 210.240 62.390 210.380 ;
        RECT 62.650 210.320 62.910 210.640 ;
        RECT 63.110 210.320 63.370 210.640 ;
        RECT 60.285 209.105 61.825 209.475 ;
        RECT 60.285 203.665 61.825 204.035 ;
        RECT 61.730 201.820 61.990 202.140 ;
        RECT 59.890 201.480 60.150 201.800 ;
        RECT 59.880 200.605 60.160 200.975 ;
        RECT 61.790 200.780 61.930 201.820 ;
        RECT 59.950 200.100 60.090 200.605 ;
        RECT 61.730 200.460 61.990 200.780 ;
        RECT 62.250 200.100 62.390 210.240 ;
        RECT 62.710 206.220 62.850 210.320 ;
        RECT 63.170 208.260 63.310 210.320 ;
        RECT 64.030 208.620 64.290 208.940 ;
        RECT 63.110 207.940 63.370 208.260 ;
        RECT 62.650 205.900 62.910 206.220 ;
        RECT 62.710 200.860 62.850 205.900 ;
        RECT 63.110 204.200 63.370 204.520 ;
        RECT 63.170 203.160 63.310 204.200 ;
        RECT 63.110 202.840 63.370 203.160 ;
        RECT 62.710 200.720 63.770 200.860 ;
        RECT 63.110 200.120 63.370 200.440 ;
        RECT 59.890 199.780 60.150 200.100 ;
        RECT 62.190 199.780 62.450 200.100 ;
        RECT 59.890 198.760 60.150 199.080 ;
        RECT 59.950 197.970 60.090 198.760 ;
        RECT 60.285 198.225 61.825 198.595 ;
        RECT 59.950 197.830 60.550 197.970 ;
        RECT 59.880 196.525 60.160 196.895 ;
        RECT 59.890 196.380 60.150 196.525 ;
        RECT 59.880 195.845 60.160 196.215 ;
        RECT 58.960 194.485 59.240 194.855 ;
        RECT 59.430 194.680 59.690 195.000 ;
        RECT 59.950 192.620 60.090 195.845 ;
        RECT 60.410 194.660 60.550 197.830 ;
        RECT 62.650 197.630 62.910 197.720 ;
        RECT 62.250 197.490 62.910 197.630 ;
        RECT 60.810 196.040 61.070 196.360 ;
        RECT 60.870 195.000 61.010 196.040 ;
        RECT 60.810 194.680 61.070 195.000 ;
        RECT 60.350 194.340 60.610 194.660 ;
        RECT 60.410 194.175 60.550 194.340 ;
        RECT 60.340 193.805 60.620 194.175 ;
        RECT 60.285 192.785 61.825 193.155 ;
        RECT 59.890 192.300 60.150 192.620 ;
        RECT 59.430 191.620 59.690 191.940 ;
        RECT 58.510 189.580 58.770 189.900 ;
        RECT 58.970 189.240 59.230 189.560 ;
        RECT 58.050 188.900 58.310 189.220 ;
        RECT 57.590 188.560 57.850 188.880 ;
        RECT 57.650 185.335 57.790 188.560 ;
        RECT 58.110 186.500 58.250 188.900 ;
        RECT 59.030 186.840 59.170 189.240 ;
        RECT 59.490 188.540 59.630 191.620 ;
        RECT 59.430 188.220 59.690 188.540 ;
        RECT 59.890 188.220 60.150 188.540 ;
        RECT 59.490 187.180 59.630 188.220 ;
        RECT 59.430 186.860 59.690 187.180 ;
        RECT 58.970 186.520 59.230 186.840 ;
        RECT 58.050 186.180 58.310 186.500 ;
        RECT 59.420 185.645 59.700 186.015 ;
        RECT 59.490 185.480 59.630 185.645 ;
        RECT 57.580 184.965 57.860 185.335 ;
        RECT 59.430 185.160 59.690 185.480 ;
        RECT 59.950 184.120 60.090 188.220 ;
        RECT 60.285 187.345 61.825 187.715 ;
        RECT 62.250 186.840 62.390 197.490 ;
        RECT 62.650 197.400 62.910 197.490 ;
        RECT 62.650 196.720 62.910 197.040 ;
        RECT 62.710 189.900 62.850 196.720 ;
        RECT 63.170 194.320 63.310 200.120 ;
        RECT 63.630 198.990 63.770 200.720 ;
        RECT 64.090 199.760 64.230 208.620 ;
        RECT 64.030 199.440 64.290 199.760 ;
        RECT 63.630 198.850 64.230 198.990 ;
        RECT 64.090 196.700 64.230 198.850 ;
        RECT 64.030 196.380 64.290 196.700 ;
        RECT 63.570 196.040 63.830 196.360 ;
        RECT 63.630 194.320 63.770 196.040 ;
        RECT 63.110 194.000 63.370 194.320 ;
        RECT 63.570 194.000 63.830 194.320 ;
        RECT 64.090 192.280 64.230 196.380 ;
        RECT 64.030 191.960 64.290 192.280 ;
        RECT 63.570 190.600 63.830 190.920 ;
        RECT 63.630 189.900 63.770 190.600 ;
        RECT 62.650 189.580 62.910 189.900 ;
        RECT 63.570 189.580 63.830 189.900 ;
        RECT 63.570 188.900 63.830 189.220 ;
        RECT 62.190 186.520 62.450 186.840 ;
        RECT 63.630 186.750 63.770 188.900 ;
        RECT 64.030 186.750 64.290 186.840 ;
        RECT 63.630 186.610 64.290 186.750 ;
        RECT 64.030 186.520 64.290 186.610 ;
        RECT 62.190 185.840 62.450 186.160 ;
        RECT 59.890 183.800 60.150 184.120 ;
        RECT 58.510 183.460 58.770 183.780 ;
        RECT 58.050 182.440 58.310 182.760 ;
        RECT 57.590 180.740 57.850 181.060 ;
        RECT 53.450 178.700 53.710 179.020 ;
        RECT 53.450 178.020 53.710 178.340 ;
        RECT 52.990 174.960 53.250 175.280 ;
        RECT 51.610 174.710 52.270 174.850 ;
        RECT 51.610 174.620 51.870 174.710 ;
        RECT 51.150 173.260 51.410 173.580 ;
        RECT 53.510 173.095 53.650 178.020 ;
        RECT 53.970 175.960 54.110 179.720 ;
        RECT 56.270 178.340 56.410 179.720 ;
        RECT 56.660 179.525 56.940 179.895 ;
        RECT 56.210 178.020 56.470 178.340 ;
        RECT 56.670 178.020 56.930 178.340 ;
        RECT 54.830 175.980 55.090 176.300 ;
        RECT 53.910 175.640 54.170 175.960 ;
        RECT 54.360 175.445 54.640 175.815 ;
        RECT 53.910 175.135 54.170 175.280 ;
        RECT 53.900 174.765 54.180 175.135 ;
        RECT 50.290 172.670 50.890 172.810 ;
        RECT 50.750 172.220 50.890 172.670 ;
        RECT 52.070 172.580 52.330 172.900 ;
        RECT 53.440 172.725 53.720 173.095 ;
        RECT 50.230 171.900 50.490 172.220 ;
        RECT 50.690 171.900 50.950 172.220 ;
        RECT 49.760 171.365 50.040 171.735 ;
        RECT 49.310 169.520 49.570 169.840 ;
        RECT 49.370 167.120 49.510 169.520 ;
        RECT 49.830 169.160 49.970 171.365 ;
        RECT 50.290 170.375 50.430 171.900 ;
        RECT 50.750 170.520 50.890 171.900 ;
        RECT 50.220 170.005 50.500 170.375 ;
        RECT 50.690 170.200 50.950 170.520 ;
        RECT 49.770 168.840 50.030 169.160 ;
        RECT 49.770 167.480 50.030 167.800 ;
        RECT 49.310 166.800 49.570 167.120 ;
        RECT 48.850 164.760 49.110 165.080 ;
        RECT 48.910 159.300 49.050 164.760 ;
        RECT 49.830 161.000 49.970 167.480 ;
        RECT 50.290 165.420 50.430 170.005 ;
        RECT 51.150 169.520 51.410 169.840 ;
        RECT 50.690 167.140 50.950 167.460 ;
        RECT 50.750 165.420 50.890 167.140 ;
        RECT 50.230 165.100 50.490 165.420 ;
        RECT 50.690 165.100 50.950 165.420 ;
        RECT 50.750 164.400 50.890 165.100 ;
        RECT 50.690 164.080 50.950 164.400 ;
        RECT 50.680 163.205 50.960 163.575 ;
        RECT 50.750 162.020 50.890 163.205 ;
        RECT 51.210 162.700 51.350 169.520 ;
        RECT 51.600 165.925 51.880 166.295 ;
        RECT 51.150 162.380 51.410 162.700 ;
        RECT 50.690 161.700 50.950 162.020 ;
        RECT 49.770 160.680 50.030 161.000 ;
        RECT 48.850 158.980 49.110 159.300 ;
        RECT 49.310 158.300 49.570 158.620 ;
        RECT 49.370 156.240 49.510 158.300 ;
        RECT 49.310 155.920 49.570 156.240 ;
        RECT 49.830 156.095 49.970 160.680 ;
        RECT 50.230 158.640 50.490 158.960 ;
        RECT 48.390 155.240 48.650 155.560 ;
        RECT 47.070 153.120 47.670 153.260 ;
        RECT 47.930 153.200 48.190 153.520 ;
        RECT 48.450 153.430 48.590 155.240 ;
        RECT 49.370 154.540 49.510 155.920 ;
        RECT 49.760 155.725 50.040 156.095 ;
        RECT 49.830 155.560 49.970 155.725 ;
        RECT 49.770 155.240 50.030 155.560 ;
        RECT 49.310 154.220 49.570 154.540 ;
        RECT 48.850 153.430 49.110 153.520 ;
        RECT 48.450 153.290 49.110 153.430 ;
        RECT 48.850 153.200 49.110 153.290 ;
        RECT 49.770 153.200 50.030 153.520 ;
        RECT 46.550 152.520 46.810 152.840 ;
        RECT 47.010 152.520 47.270 152.840 ;
        RECT 46.610 151.140 46.750 152.520 ;
        RECT 46.550 150.820 46.810 151.140 ;
        RECT 46.550 149.800 46.810 150.120 ;
        RECT 46.610 149.100 46.750 149.800 ;
        RECT 46.550 148.780 46.810 149.100 ;
        RECT 46.090 148.100 46.350 148.420 ;
        RECT 46.550 147.080 46.810 147.400 ;
        RECT 45.690 146.150 46.290 146.290 ;
        RECT 45.630 145.380 45.890 145.700 ;
        RECT 45.170 145.040 45.430 145.360 ;
        RECT 45.230 142.980 45.370 145.040 ;
        RECT 45.170 142.660 45.430 142.980 ;
        RECT 45.690 137.450 45.830 145.380 ;
        RECT 46.150 142.640 46.290 146.150 ;
        RECT 46.090 142.320 46.350 142.640 ;
        RECT 46.080 141.445 46.360 141.815 ;
        RECT 46.150 140.940 46.290 141.445 ;
        RECT 46.090 140.620 46.350 140.940 ;
        RECT 46.090 137.450 46.350 137.540 ;
        RECT 45.690 137.310 46.350 137.450 ;
        RECT 46.090 137.220 46.350 137.310 ;
        RECT 44.710 135.180 44.970 135.500 ;
        RECT 46.150 135.160 46.290 137.220 ;
        RECT 46.090 135.070 46.350 135.160 ;
        RECT 45.690 134.930 46.350 135.070 ;
        RECT 44.250 132.460 44.510 132.780 ;
        RECT 43.790 131.100 44.050 131.420 ;
        RECT 45.170 131.100 45.430 131.420 ;
        RECT 44.250 128.720 44.510 129.040 ;
        RECT 43.790 128.270 44.050 128.360 ;
        RECT 43.390 128.130 44.050 128.270 ;
        RECT 42.870 127.020 43.130 127.340 ;
        RECT 42.410 126.340 42.670 126.660 ;
        RECT 35.510 126.000 35.770 126.320 ;
        RECT 39.650 126.000 39.910 126.320 ;
        RECT 12.510 125.660 12.770 125.980 ;
        RECT 37.350 125.320 37.610 125.640 ;
        RECT 37.410 124.620 37.550 125.320 ;
        RECT 40.850 124.785 42.390 125.155 ;
        RECT 37.350 124.300 37.610 124.620 ;
        RECT 43.390 123.940 43.530 128.130 ;
        RECT 43.790 128.040 44.050 128.130 ;
        RECT 44.310 127.000 44.450 128.720 ;
        RECT 45.230 128.360 45.370 131.100 ;
        RECT 45.690 129.720 45.830 134.930 ;
        RECT 46.090 134.840 46.350 134.930 ;
        RECT 46.610 133.710 46.750 147.080 ;
        RECT 47.070 140.600 47.210 152.520 ;
        RECT 47.530 144.680 47.670 153.120 ;
        RECT 47.920 151.645 48.200 152.015 ;
        RECT 49.300 151.645 49.580 152.015 ;
        RECT 47.470 144.360 47.730 144.680 ;
        RECT 47.470 143.340 47.730 143.660 ;
        RECT 47.530 141.960 47.670 143.340 ;
        RECT 47.470 141.640 47.730 141.960 ;
        RECT 47.010 140.280 47.270 140.600 ;
        RECT 47.990 140.455 48.130 151.645 ;
        RECT 48.390 150.820 48.650 151.140 ;
        RECT 48.840 150.965 49.120 151.335 ;
        RECT 48.450 145.360 48.590 150.820 ;
        RECT 48.910 149.975 49.050 150.965 ;
        RECT 49.370 150.800 49.510 151.645 ;
        RECT 49.830 151.220 49.970 153.200 ;
        RECT 50.290 151.820 50.430 158.640 ;
        RECT 50.690 158.135 50.950 158.280 ;
        RECT 50.680 157.765 50.960 158.135 ;
        RECT 50.750 153.430 50.890 157.765 ;
        RECT 51.150 156.600 51.410 156.920 ;
        RECT 51.210 154.540 51.350 156.600 ;
        RECT 51.670 156.580 51.810 165.925 ;
        RECT 52.130 162.700 52.270 172.580 ;
        RECT 52.530 172.240 52.790 172.560 ;
        RECT 52.590 170.260 52.730 172.240 ;
        RECT 53.450 171.900 53.710 172.220 ;
        RECT 52.990 170.260 53.250 170.520 ;
        RECT 52.590 170.200 53.250 170.260 ;
        RECT 52.590 170.120 53.190 170.200 ;
        RECT 52.590 166.295 52.730 170.120 ;
        RECT 53.510 169.840 53.650 171.900 ;
        RECT 53.910 171.560 54.170 171.880 ;
        RECT 53.970 170.860 54.110 171.560 ;
        RECT 53.910 170.540 54.170 170.860 ;
        RECT 54.430 169.840 54.570 175.445 ;
        RECT 54.890 170.860 55.030 175.980 ;
        RECT 55.750 175.300 56.010 175.620 ;
        RECT 55.290 174.280 55.550 174.600 ;
        RECT 55.810 174.455 55.950 175.300 ;
        RECT 55.350 172.560 55.490 174.280 ;
        RECT 55.740 174.085 56.020 174.455 ;
        RECT 55.290 172.240 55.550 172.560 ;
        RECT 55.750 171.900 56.010 172.220 ;
        RECT 55.280 171.365 55.560 171.735 ;
        RECT 54.830 170.540 55.090 170.860 ;
        RECT 53.450 169.520 53.710 169.840 ;
        RECT 54.370 169.520 54.630 169.840 ;
        RECT 54.830 169.520 55.090 169.840 ;
        RECT 53.450 167.140 53.710 167.460 ;
        RECT 52.990 166.460 53.250 166.780 ;
        RECT 52.520 165.925 52.800 166.295 ;
        RECT 52.530 164.420 52.790 164.740 ;
        RECT 52.590 163.575 52.730 164.420 ;
        RECT 52.520 163.205 52.800 163.575 ;
        RECT 52.070 162.380 52.330 162.700 ;
        RECT 52.530 162.040 52.790 162.360 ;
        RECT 52.590 158.280 52.730 162.040 ;
        RECT 52.530 157.960 52.790 158.280 ;
        RECT 52.530 156.940 52.790 157.260 ;
        RECT 51.610 156.260 51.870 156.580 ;
        RECT 51.670 154.540 51.810 156.260 ;
        RECT 52.060 155.725 52.340 156.095 ;
        RECT 51.150 154.220 51.410 154.540 ;
        RECT 51.610 154.220 51.870 154.540 ;
        RECT 51.210 153.770 51.350 154.220 ;
        RECT 51.210 153.630 51.810 153.770 ;
        RECT 50.750 153.290 51.350 153.430 ;
        RECT 50.690 152.520 50.950 152.840 ;
        RECT 51.210 152.580 51.350 153.290 ;
        RECT 51.670 153.180 51.810 153.630 ;
        RECT 51.610 152.860 51.870 153.180 ;
        RECT 50.230 151.500 50.490 151.820 ;
        RECT 49.830 151.080 50.430 151.220 ;
        RECT 49.310 150.480 49.570 150.800 ;
        RECT 49.770 150.480 50.030 150.800 ;
        RECT 48.840 149.605 49.120 149.975 ;
        RECT 49.310 149.800 49.570 150.120 ;
        RECT 48.850 148.440 49.110 148.760 ;
        RECT 49.370 148.670 49.510 149.800 ;
        RECT 49.830 149.295 49.970 150.480 ;
        RECT 49.760 148.925 50.040 149.295 ;
        RECT 49.370 148.530 49.970 148.670 ;
        RECT 48.910 145.700 49.050 148.440 ;
        RECT 49.830 148.080 49.970 148.530 ;
        RECT 50.290 148.080 50.430 151.080 ;
        RECT 50.750 148.420 50.890 152.520 ;
        RECT 51.210 152.440 51.810 152.580 ;
        RECT 51.140 151.645 51.420 152.015 ;
        RECT 51.210 149.100 51.350 151.645 ;
        RECT 51.670 150.800 51.810 152.440 ;
        RECT 51.610 150.480 51.870 150.800 ;
        RECT 51.150 148.780 51.410 149.100 ;
        RECT 50.690 148.100 50.950 148.420 ;
        RECT 49.310 147.760 49.570 148.080 ;
        RECT 49.770 147.760 50.030 148.080 ;
        RECT 50.230 147.760 50.490 148.080 ;
        RECT 48.850 145.380 49.110 145.700 ;
        RECT 48.390 145.040 48.650 145.360 ;
        RECT 48.450 142.980 48.590 145.040 ;
        RECT 48.840 144.845 49.120 145.215 ;
        RECT 48.910 144.680 49.050 144.845 ;
        RECT 48.850 144.360 49.110 144.680 ;
        RECT 49.370 143.660 49.510 147.760 ;
        RECT 49.770 147.080 50.030 147.400 ;
        RECT 49.310 143.340 49.570 143.660 ;
        RECT 48.390 142.660 48.650 142.980 ;
        RECT 48.840 141.445 49.120 141.815 ;
        RECT 47.920 140.085 48.200 140.455 ;
        RECT 47.470 137.900 47.730 138.220 ;
        RECT 47.010 133.710 47.270 133.800 ;
        RECT 46.610 133.570 47.270 133.710 ;
        RECT 47.010 133.480 47.270 133.570 ;
        RECT 46.550 132.120 46.810 132.440 ;
        RECT 46.090 131.780 46.350 132.100 ;
        RECT 46.150 130.060 46.290 131.780 ;
        RECT 46.610 130.060 46.750 132.120 ;
        RECT 46.090 129.740 46.350 130.060 ;
        RECT 46.550 129.740 46.810 130.060 ;
        RECT 45.630 129.400 45.890 129.720 ;
        RECT 47.070 129.040 47.210 133.480 ;
        RECT 47.530 131.080 47.670 137.900 ;
        RECT 47.990 132.780 48.130 140.085 ;
        RECT 47.930 132.460 48.190 132.780 ;
        RECT 48.910 131.420 49.050 141.445 ;
        RECT 48.850 131.100 49.110 131.420 ;
        RECT 47.470 130.760 47.730 131.080 ;
        RECT 49.830 129.040 49.970 147.080 ;
        RECT 50.230 146.060 50.490 146.380 ;
        RECT 50.290 145.700 50.430 146.060 ;
        RECT 50.230 145.380 50.490 145.700 ;
        RECT 50.750 144.680 50.890 148.100 ;
        RECT 51.150 147.935 51.410 148.080 ;
        RECT 51.140 147.565 51.420 147.935 ;
        RECT 52.130 146.380 52.270 155.725 ;
        RECT 52.590 153.860 52.730 156.940 ;
        RECT 52.530 153.540 52.790 153.860 ;
        RECT 52.530 152.860 52.790 153.180 ;
        RECT 52.070 146.060 52.330 146.380 ;
        RECT 52.060 145.525 52.340 145.895 ;
        RECT 50.690 144.360 50.950 144.680 ;
        RECT 51.600 144.165 51.880 144.535 ;
        RECT 51.150 142.660 51.410 142.980 ;
        RECT 51.210 140.260 51.350 142.660 ;
        RECT 51.670 141.135 51.810 144.165 ;
        RECT 51.600 140.765 51.880 141.135 ;
        RECT 51.670 140.260 51.810 140.765 ;
        RECT 52.130 140.260 52.270 145.525 ;
        RECT 51.150 139.940 51.410 140.260 ;
        RECT 51.610 139.940 51.870 140.260 ;
        RECT 52.070 139.940 52.330 140.260 ;
        RECT 51.600 138.725 51.880 139.095 ;
        RECT 51.670 138.220 51.810 138.725 ;
        RECT 51.610 137.900 51.870 138.220 ;
        RECT 51.610 136.540 51.870 136.860 ;
        RECT 51.670 136.375 51.810 136.540 ;
        RECT 51.600 136.005 51.880 136.375 ;
        RECT 47.010 128.720 47.270 129.040 ;
        RECT 49.770 128.720 50.030 129.040 ;
        RECT 45.170 128.040 45.430 128.360 ;
        RECT 44.250 126.680 44.510 127.000 ;
        RECT 45.230 126.320 45.370 128.040 ;
        RECT 45.170 126.000 45.430 126.320 ;
        RECT 46.090 125.320 46.350 125.640 ;
        RECT 46.150 124.620 46.290 125.320 ;
        RECT 49.830 125.240 49.970 128.720 ;
        RECT 51.670 125.640 51.810 136.005 ;
        RECT 52.130 135.695 52.270 139.940 ;
        RECT 52.060 135.325 52.340 135.695 ;
        RECT 52.070 134.500 52.330 134.820 ;
        RECT 52.130 132.780 52.270 134.500 ;
        RECT 52.070 132.460 52.330 132.780 ;
        RECT 52.590 131.420 52.730 152.860 ;
        RECT 53.050 148.080 53.190 166.460 ;
        RECT 53.510 157.455 53.650 167.140 ;
        RECT 54.890 167.120 55.030 169.520 ;
        RECT 55.350 167.800 55.490 171.365 ;
        RECT 55.290 167.480 55.550 167.800 ;
        RECT 55.810 167.710 55.950 171.900 ;
        RECT 56.270 170.180 56.410 178.020 ;
        RECT 56.210 169.860 56.470 170.180 ;
        RECT 56.730 169.840 56.870 178.020 ;
        RECT 57.650 178.000 57.790 180.740 ;
        RECT 57.590 177.680 57.850 178.000 ;
        RECT 57.130 177.000 57.390 177.320 ;
        RECT 57.590 177.000 57.850 177.320 ;
        RECT 57.190 176.300 57.330 177.000 ;
        RECT 57.130 175.980 57.390 176.300 ;
        RECT 57.650 172.900 57.790 177.000 ;
        RECT 57.590 172.580 57.850 172.900 ;
        RECT 58.110 170.860 58.250 182.440 ;
        RECT 58.570 174.940 58.710 183.460 ;
        RECT 59.430 183.120 59.690 183.440 ;
        RECT 59.490 181.740 59.630 183.120 ;
        RECT 59.890 182.780 60.150 183.100 ;
        RECT 59.950 181.740 60.090 182.780 ;
        RECT 60.285 181.905 61.825 182.275 ;
        RECT 59.430 181.420 59.690 181.740 ;
        RECT 59.890 181.420 60.150 181.740 ;
        RECT 59.950 180.970 60.090 181.420 ;
        RECT 59.490 180.830 60.090 180.970 ;
        RECT 59.490 180.575 59.630 180.830 ;
        RECT 59.420 180.205 59.700 180.575 ;
        RECT 59.890 180.060 60.150 180.380 ;
        RECT 58.960 179.525 59.240 179.895 ;
        RECT 59.030 177.855 59.170 179.525 ;
        RECT 59.950 179.100 60.090 180.060 ;
        RECT 59.950 178.960 61.470 179.100 ;
        RECT 61.330 178.680 61.470 178.960 ;
        RECT 61.730 178.930 61.990 179.020 ;
        RECT 62.250 178.930 62.390 185.840 ;
        RECT 62.640 185.645 62.920 186.015 ;
        RECT 62.710 184.120 62.850 185.645 ;
        RECT 62.650 183.800 62.910 184.120 ;
        RECT 64.090 183.780 64.230 186.520 ;
        RECT 64.030 183.460 64.290 183.780 ;
        RECT 63.560 182.925 63.840 183.295 ;
        RECT 61.730 178.790 62.390 178.930 ;
        RECT 61.730 178.700 61.990 178.790 ;
        RECT 60.350 178.360 60.610 178.680 ;
        RECT 61.270 178.420 61.530 178.680 ;
        RECT 61.270 178.360 61.930 178.420 ;
        RECT 60.410 178.000 60.550 178.360 ;
        RECT 61.330 178.280 61.930 178.360 ;
        RECT 59.890 177.910 60.150 178.000 ;
        RECT 58.960 177.485 59.240 177.855 ;
        RECT 59.490 177.770 60.150 177.910 ;
        RECT 58.510 174.620 58.770 174.940 ;
        RECT 58.570 172.900 58.710 174.620 ;
        RECT 59.490 173.580 59.630 177.770 ;
        RECT 59.890 177.680 60.150 177.770 ;
        RECT 60.350 177.680 60.610 178.000 ;
        RECT 61.790 177.740 61.930 178.280 ;
        RECT 61.790 177.600 62.160 177.740 ;
        RECT 59.890 177.000 60.150 177.320 ;
        RECT 59.950 175.620 60.090 177.000 ;
        RECT 60.285 176.465 61.825 176.835 ;
        RECT 62.020 175.700 62.160 177.600 ;
        RECT 59.890 175.300 60.150 175.620 ;
        RECT 61.790 175.560 62.160 175.700 ;
        RECT 59.430 173.260 59.690 173.580 ;
        RECT 58.510 172.580 58.770 172.900 ;
        RECT 58.970 172.240 59.230 172.560 ;
        RECT 59.430 172.240 59.690 172.560 ;
        RECT 58.050 170.540 58.310 170.860 ;
        RECT 59.030 170.180 59.170 172.240 ;
        RECT 59.490 170.860 59.630 172.240 ;
        RECT 59.430 170.540 59.690 170.860 ;
        RECT 58.970 169.860 59.230 170.180 ;
        RECT 56.670 169.520 56.930 169.840 ;
        RECT 58.510 169.695 58.770 169.840 ;
        RECT 58.500 169.325 58.780 169.695 ;
        RECT 59.430 169.520 59.690 169.840 ;
        RECT 57.590 168.840 57.850 169.160 ;
        RECT 56.210 167.710 56.470 167.800 ;
        RECT 55.810 167.570 56.470 167.710 ;
        RECT 54.830 166.800 55.090 167.120 ;
        RECT 53.910 166.120 54.170 166.440 ;
        RECT 53.970 160.060 54.110 166.120 ;
        RECT 54.360 165.245 54.640 165.615 ;
        RECT 54.430 161.680 54.570 165.245 ;
        RECT 54.830 163.575 55.090 163.720 ;
        RECT 54.820 163.205 55.100 163.575 ;
        RECT 55.290 161.700 55.550 162.020 ;
        RECT 54.370 161.360 54.630 161.680 ;
        RECT 54.430 160.855 54.570 161.360 ;
        RECT 55.350 161.000 55.490 161.700 ;
        RECT 55.810 161.680 55.950 167.570 ;
        RECT 56.210 167.480 56.470 167.570 ;
        RECT 56.670 167.480 56.930 167.800 ;
        RECT 57.650 167.655 57.790 168.840 ;
        RECT 59.490 167.800 59.630 169.520 ;
        RECT 56.730 167.120 56.870 167.480 ;
        RECT 57.130 167.140 57.390 167.460 ;
        RECT 57.580 167.285 57.860 167.655 ;
        RECT 59.430 167.480 59.690 167.800 ;
        RECT 57.590 167.140 57.850 167.285 ;
        RECT 58.510 167.140 58.770 167.460 ;
        RECT 56.670 166.975 56.930 167.120 ;
        RECT 56.660 166.860 56.940 166.975 ;
        RECT 56.270 166.720 56.940 166.860 ;
        RECT 56.270 162.020 56.410 166.720 ;
        RECT 56.660 166.605 56.940 166.720 ;
        RECT 56.660 164.565 56.940 164.935 ;
        RECT 56.730 164.060 56.870 164.565 ;
        RECT 56.670 163.740 56.930 164.060 ;
        RECT 56.210 161.700 56.470 162.020 ;
        RECT 55.750 161.360 56.010 161.680 ;
        RECT 56.730 161.420 56.870 163.740 ;
        RECT 57.190 162.020 57.330 167.140 ;
        RECT 57.650 162.020 57.790 167.140 ;
        RECT 58.050 166.460 58.310 166.780 ;
        RECT 58.110 164.740 58.250 166.460 ;
        RECT 58.050 164.420 58.310 164.740 ;
        RECT 57.130 161.700 57.390 162.020 ;
        RECT 57.590 161.700 57.850 162.020 ;
        RECT 56.730 161.280 57.330 161.420 ;
        RECT 58.050 161.360 58.310 161.680 ;
        RECT 54.360 160.485 54.640 160.855 ;
        RECT 55.290 160.680 55.550 161.000 ;
        RECT 55.750 160.680 56.010 161.000 ;
        RECT 55.810 160.060 55.950 160.680 ;
        RECT 53.970 159.920 55.950 160.060 ;
        RECT 57.190 158.530 57.330 161.280 ;
        RECT 58.110 160.740 58.250 161.360 ;
        RECT 57.650 160.600 58.250 160.740 ;
        RECT 57.650 159.980 57.790 160.600 ;
        RECT 57.590 159.660 57.850 159.980 ;
        RECT 58.050 159.660 58.310 159.980 ;
        RECT 58.110 159.300 58.250 159.660 ;
        RECT 58.050 158.980 58.310 159.300 ;
        RECT 58.570 158.620 58.710 167.140 ;
        RECT 59.950 167.120 60.090 175.300 ;
        RECT 61.790 174.940 61.930 175.560 ;
        RECT 61.730 174.620 61.990 174.940 ;
        RECT 62.650 171.560 62.910 171.880 ;
        RECT 60.285 171.025 61.825 171.395 ;
        RECT 60.340 170.005 60.620 170.375 ;
        RECT 59.890 166.800 60.150 167.120 ;
        RECT 58.960 165.925 59.240 166.295 ;
        RECT 59.430 166.120 59.690 166.440 ;
        RECT 60.410 166.350 60.550 170.005 ;
        RECT 62.180 168.645 62.460 169.015 ;
        RECT 60.810 167.480 61.070 167.800 ;
        RECT 60.870 167.030 61.010 167.480 ;
        RECT 61.270 167.030 61.530 167.120 ;
        RECT 60.870 166.890 61.530 167.030 ;
        RECT 61.270 166.800 61.530 166.890 ;
        RECT 59.950 166.210 60.550 166.350 ;
        RECT 59.030 163.720 59.170 165.925 ;
        RECT 58.970 163.400 59.230 163.720 ;
        RECT 59.490 162.700 59.630 166.120 ;
        RECT 58.970 162.380 59.230 162.700 ;
        RECT 59.430 162.380 59.690 162.700 ;
        RECT 59.030 159.980 59.170 162.380 ;
        RECT 59.430 161.020 59.690 161.340 ;
        RECT 59.490 160.855 59.630 161.020 ;
        RECT 59.420 160.485 59.700 160.855 ;
        RECT 59.950 159.980 60.090 166.210 ;
        RECT 60.285 165.585 61.825 165.955 ;
        RECT 62.250 164.740 62.390 168.645 ;
        RECT 62.710 167.800 62.850 171.560 ;
        RECT 63.630 170.180 63.770 182.925 ;
        RECT 64.550 177.740 64.690 213.040 ;
        RECT 65.930 211.660 66.070 213.040 ;
        RECT 65.870 211.340 66.130 211.660 ;
        RECT 64.950 211.000 65.210 211.320 ;
        RECT 65.410 211.000 65.670 211.320 ;
        RECT 65.010 207.920 65.150 211.000 ;
        RECT 64.950 207.600 65.210 207.920 ;
        RECT 65.010 205.880 65.150 207.600 ;
        RECT 64.950 205.560 65.210 205.880 ;
        RECT 65.470 204.520 65.610 211.000 ;
        RECT 66.390 208.455 66.530 216.100 ;
        RECT 66.320 208.085 66.600 208.455 ;
        RECT 66.790 205.220 67.050 205.540 ;
        RECT 65.410 204.200 65.670 204.520 ;
        RECT 64.940 203.325 65.220 203.695 ;
        RECT 65.010 203.160 65.150 203.325 ;
        RECT 64.950 202.840 65.210 203.160 ;
        RECT 66.850 203.015 66.990 205.220 ;
        RECT 65.010 191.940 65.150 202.840 ;
        RECT 66.780 202.645 67.060 203.015 ;
        RECT 66.330 202.160 66.590 202.480 ;
        RECT 66.780 202.220 67.060 202.335 ;
        RECT 67.310 202.220 67.450 218.570 ;
        RECT 67.710 218.480 67.970 218.570 ;
        RECT 68.230 208.940 68.370 219.160 ;
        RECT 68.690 217.100 68.830 221.005 ;
        RECT 69.080 220.325 69.360 220.695 ;
        RECT 69.150 219.820 69.290 220.325 ;
        RECT 69.090 219.500 69.350 219.820 ;
        RECT 69.550 218.820 69.810 219.140 ;
        RECT 73.680 218.965 73.960 219.335 ;
        RECT 69.610 218.120 69.750 218.820 ;
        RECT 72.770 218.140 73.030 218.460 ;
        RECT 69.550 217.800 69.810 218.120 ;
        RECT 70.930 217.975 71.190 218.120 ;
        RECT 68.630 216.780 68.890 217.100 ;
        RECT 69.610 216.420 69.750 217.800 ;
        RECT 70.920 217.605 71.200 217.975 ;
        RECT 71.850 217.800 72.110 218.120 ;
        RECT 71.910 217.100 72.050 217.800 ;
        RECT 71.850 216.780 72.110 217.100 ;
        RECT 69.550 216.100 69.810 216.420 ;
        RECT 70.470 216.100 70.730 216.420 ;
        RECT 69.090 215.760 69.350 216.080 ;
        RECT 68.630 215.080 68.890 215.400 ;
        RECT 68.690 214.575 68.830 215.080 ;
        RECT 68.620 214.205 68.900 214.575 ;
        RECT 69.150 214.040 69.290 215.760 ;
        RECT 70.010 214.060 70.270 214.380 ;
        RECT 69.090 213.720 69.350 214.040 ;
        RECT 68.170 208.620 68.430 208.940 ;
        RECT 68.170 207.600 68.430 207.920 ;
        RECT 69.550 207.775 69.810 207.920 ;
        RECT 68.230 205.540 68.370 207.600 ;
        RECT 68.630 207.260 68.890 207.580 ;
        RECT 69.540 207.405 69.820 207.775 ;
        RECT 68.690 206.415 68.830 207.260 ;
        RECT 69.090 206.920 69.350 207.240 ;
        RECT 68.620 206.045 68.900 206.415 ;
        RECT 68.690 205.540 68.830 206.045 ;
        RECT 68.170 205.220 68.430 205.540 ;
        RECT 68.630 205.220 68.890 205.540 ;
        RECT 65.410 196.720 65.670 197.040 ;
        RECT 65.870 196.720 66.130 197.040 ;
        RECT 65.470 195.340 65.610 196.720 ;
        RECT 65.930 196.360 66.070 196.720 ;
        RECT 65.870 196.040 66.130 196.360 ;
        RECT 65.410 195.020 65.670 195.340 ;
        RECT 65.410 194.000 65.670 194.320 ;
        RECT 64.950 191.620 65.210 191.940 ;
        RECT 65.470 190.920 65.610 194.000 ;
        RECT 65.870 193.320 66.130 193.640 ;
        RECT 65.410 190.600 65.670 190.920 ;
        RECT 65.930 189.220 66.070 193.320 ;
        RECT 65.870 188.900 66.130 189.220 ;
        RECT 66.390 189.130 66.530 202.160 ;
        RECT 66.780 202.080 67.450 202.220 ;
        RECT 66.780 201.965 67.060 202.080 ;
        RECT 67.250 201.480 67.510 201.800 ;
        RECT 66.790 199.440 67.050 199.760 ;
        RECT 66.850 194.660 66.990 199.440 ;
        RECT 67.310 196.360 67.450 201.480 ;
        RECT 67.700 199.925 67.980 200.295 ;
        RECT 67.710 199.780 67.970 199.925 ;
        RECT 68.170 199.780 68.430 200.100 ;
        RECT 68.230 197.380 68.370 199.780 ;
        RECT 68.170 197.060 68.430 197.380 ;
        RECT 67.250 196.040 67.510 196.360 ;
        RECT 66.790 194.340 67.050 194.660 ;
        RECT 66.790 193.660 67.050 193.980 ;
        RECT 66.850 192.620 66.990 193.660 ;
        RECT 66.790 192.300 67.050 192.620 ;
        RECT 66.850 189.980 66.990 192.300 ;
        RECT 67.310 190.920 67.450 196.040 ;
        RECT 67.700 194.485 67.980 194.855 ;
        RECT 67.250 190.600 67.510 190.920 ;
        RECT 66.850 189.840 67.450 189.980 ;
        RECT 66.790 189.130 67.050 189.220 ;
        RECT 66.390 188.990 67.050 189.130 ;
        RECT 66.790 188.900 67.050 188.990 ;
        RECT 64.950 187.880 65.210 188.200 ;
        RECT 65.010 186.160 65.150 187.880 ;
        RECT 66.850 186.840 66.990 188.900 ;
        RECT 66.790 186.520 67.050 186.840 ;
        RECT 64.950 185.840 65.210 186.160 ;
        RECT 65.010 181.060 65.150 185.840 ;
        RECT 67.310 183.440 67.450 189.840 ;
        RECT 67.250 183.120 67.510 183.440 ;
        RECT 67.250 182.440 67.510 182.760 ;
        RECT 67.310 181.740 67.450 182.440 ;
        RECT 67.250 181.420 67.510 181.740 ;
        RECT 64.950 180.740 65.210 181.060 ;
        RECT 65.870 180.400 66.130 180.720 ;
        RECT 64.550 177.660 65.150 177.740 ;
        RECT 64.550 177.600 65.210 177.660 ;
        RECT 64.950 177.340 65.210 177.600 ;
        RECT 65.410 175.640 65.670 175.960 ;
        RECT 65.470 174.455 65.610 175.640 ;
        RECT 65.400 174.085 65.680 174.455 ;
        RECT 64.950 172.240 65.210 172.560 ;
        RECT 65.010 170.860 65.150 172.240 ;
        RECT 65.410 171.560 65.670 171.880 ;
        RECT 64.950 170.540 65.210 170.860 ;
        RECT 65.470 170.520 65.610 171.560 ;
        RECT 63.570 169.860 63.830 170.180 ;
        RECT 64.490 170.090 64.750 170.180 ;
        RECT 64.940 170.090 65.220 170.375 ;
        RECT 65.410 170.200 65.670 170.520 ;
        RECT 64.490 170.005 65.220 170.090 ;
        RECT 64.490 169.950 65.150 170.005 ;
        RECT 64.490 169.860 64.750 169.950 ;
        RECT 64.030 169.520 64.290 169.840 ;
        RECT 63.560 167.965 63.840 168.335 ;
        RECT 63.630 167.800 63.770 167.965 ;
        RECT 62.650 167.480 62.910 167.800 ;
        RECT 63.570 167.480 63.830 167.800 ;
        RECT 62.190 164.650 62.450 164.740 ;
        RECT 61.790 164.510 62.450 164.650 ;
        RECT 60.800 162.525 61.080 162.895 ;
        RECT 60.870 161.535 61.010 162.525 ;
        RECT 61.790 162.020 61.930 164.510 ;
        RECT 62.190 164.420 62.450 164.510 ;
        RECT 63.110 162.040 63.370 162.360 ;
        RECT 61.730 161.700 61.990 162.020 ;
        RECT 60.800 161.165 61.080 161.535 ;
        RECT 61.720 161.165 62.000 161.535 ;
        RECT 62.650 161.360 62.910 161.680 ;
        RECT 61.730 161.020 61.990 161.165 ;
        RECT 60.285 160.145 61.825 160.515 ;
        RECT 58.970 159.660 59.230 159.980 ;
        RECT 59.890 159.740 60.150 159.980 ;
        RECT 59.490 159.660 60.150 159.740 ;
        RECT 59.490 159.600 60.090 159.660 ;
        RECT 62.710 159.640 62.850 161.360 ;
        RECT 57.590 158.530 57.850 158.620 ;
        RECT 57.190 158.390 57.850 158.530 ;
        RECT 57.590 158.300 57.850 158.390 ;
        RECT 58.510 158.300 58.770 158.620 ;
        RECT 55.280 158.020 55.560 158.135 ;
        RECT 54.890 157.880 55.560 158.020 ;
        RECT 53.440 157.170 53.720 157.455 ;
        RECT 53.910 157.170 54.170 157.260 ;
        RECT 53.440 157.085 54.170 157.170 ;
        RECT 53.510 157.030 54.170 157.085 ;
        RECT 53.910 156.940 54.170 157.030 ;
        RECT 53.450 155.415 53.710 155.560 ;
        RECT 53.440 155.045 53.720 155.415 ;
        RECT 53.450 154.055 53.710 154.200 ;
        RECT 53.440 153.685 53.720 154.055 ;
        RECT 53.910 152.750 54.170 152.840 ;
        RECT 53.510 152.610 54.170 152.750 ;
        RECT 53.510 151.820 53.650 152.610 ;
        RECT 53.910 152.520 54.170 152.610 ;
        RECT 53.450 151.500 53.710 151.820 ;
        RECT 54.890 151.140 55.030 157.880 ;
        RECT 55.280 157.765 55.560 157.880 ;
        RECT 56.210 156.940 56.470 157.260 ;
        RECT 55.750 156.260 56.010 156.580 ;
        RECT 55.290 155.920 55.550 156.240 ;
        RECT 55.350 155.415 55.490 155.920 ;
        RECT 55.280 155.045 55.560 155.415 ;
        RECT 55.280 154.365 55.560 154.735 ;
        RECT 55.350 151.820 55.490 154.365 ;
        RECT 55.290 151.500 55.550 151.820 ;
        RECT 53.910 150.820 54.170 151.140 ;
        RECT 54.830 150.820 55.090 151.140 ;
        RECT 53.450 150.480 53.710 150.800 ;
        RECT 53.510 149.010 53.650 150.480 ;
        RECT 53.970 149.975 54.110 150.820 ;
        RECT 55.290 150.140 55.550 150.460 ;
        RECT 53.900 149.605 54.180 149.975 ;
        RECT 54.820 149.605 55.100 149.975 ;
        RECT 54.890 149.100 55.030 149.605 ;
        RECT 53.510 148.870 54.110 149.010 ;
        RECT 53.440 148.245 53.720 148.615 ;
        RECT 53.510 148.080 53.650 148.245 ;
        RECT 52.990 147.760 53.250 148.080 ;
        RECT 53.450 147.760 53.710 148.080 ;
        RECT 53.440 142.125 53.720 142.495 ;
        RECT 53.450 141.980 53.710 142.125 ;
        RECT 53.450 140.280 53.710 140.600 ;
        RECT 53.970 140.455 54.110 148.870 ;
        RECT 54.830 148.780 55.090 149.100 ;
        RECT 54.830 147.760 55.090 148.080 ;
        RECT 54.370 147.420 54.630 147.740 ;
        RECT 54.430 145.610 54.570 147.420 ;
        RECT 54.890 147.400 55.030 147.760 ;
        RECT 54.830 147.080 55.090 147.400 ;
        RECT 54.830 145.610 55.090 145.700 ;
        RECT 54.430 145.470 55.090 145.610 ;
        RECT 54.830 145.380 55.090 145.470 ;
        RECT 52.980 136.685 53.260 137.055 ;
        RECT 53.050 132.100 53.190 136.685 ;
        RECT 53.510 135.500 53.650 140.280 ;
        RECT 53.900 140.085 54.180 140.455 ;
        RECT 54.370 140.170 54.630 140.260 ;
        RECT 55.350 140.170 55.490 150.140 ;
        RECT 55.810 149.100 55.950 156.260 ;
        RECT 56.270 153.375 56.410 156.940 ;
        RECT 56.670 155.240 56.930 155.560 ;
        RECT 56.730 154.540 56.870 155.240 ;
        RECT 57.120 155.045 57.400 155.415 ;
        RECT 56.670 154.220 56.930 154.540 ;
        RECT 56.200 153.005 56.480 153.375 ;
        RECT 56.670 152.860 56.930 153.180 ;
        RECT 56.210 149.800 56.470 150.120 ;
        RECT 55.750 148.780 56.010 149.100 ;
        RECT 55.750 147.080 56.010 147.400 ;
        RECT 54.370 140.030 55.490 140.170 ;
        RECT 54.370 139.940 54.630 140.030 ;
        RECT 54.830 139.260 55.090 139.580 ;
        RECT 53.910 138.920 54.170 139.240 ;
        RECT 53.450 135.180 53.710 135.500 ;
        RECT 53.970 134.820 54.110 138.920 ;
        RECT 54.890 137.880 55.030 139.260 ;
        RECT 54.830 137.560 55.090 137.880 ;
        RECT 54.890 135.500 55.030 137.560 ;
        RECT 55.810 136.520 55.950 147.080 ;
        RECT 56.270 146.380 56.410 149.800 ;
        RECT 56.210 146.060 56.470 146.380 ;
        RECT 56.730 145.360 56.870 152.860 ;
        RECT 57.190 148.420 57.330 155.045 ;
        RECT 57.650 154.540 57.790 158.300 ;
        RECT 59.490 156.150 59.630 159.600 ;
        RECT 61.260 159.125 61.540 159.495 ;
        RECT 62.650 159.320 62.910 159.640 ;
        RECT 59.890 157.960 60.150 158.280 ;
        RECT 59.950 156.580 60.090 157.960 ;
        RECT 61.330 156.580 61.470 159.125 ;
        RECT 61.730 158.640 61.990 158.960 ;
        RECT 62.650 158.640 62.910 158.960 ;
        RECT 61.790 157.260 61.930 158.640 ;
        RECT 62.710 158.280 62.850 158.640 ;
        RECT 62.650 157.960 62.910 158.280 ;
        RECT 61.730 156.940 61.990 157.260 ;
        RECT 59.890 156.260 60.150 156.580 ;
        RECT 60.350 156.260 60.610 156.580 ;
        RECT 61.270 156.260 61.530 156.580 ;
        RECT 58.570 156.010 59.630 156.150 ;
        RECT 60.410 156.095 60.550 156.260 ;
        RECT 58.570 154.620 58.710 156.010 ;
        RECT 60.340 155.725 60.620 156.095 ;
        RECT 60.285 154.705 61.825 155.075 ;
        RECT 63.170 154.620 63.310 162.040 ;
        RECT 63.570 160.680 63.830 161.000 ;
        RECT 64.090 160.855 64.230 169.520 ;
        RECT 64.950 167.820 65.210 168.140 ;
        RECT 63.630 159.980 63.770 160.680 ;
        RECT 64.020 160.485 64.300 160.855 ;
        RECT 63.570 159.660 63.830 159.980 ;
        RECT 64.490 158.980 64.750 159.300 ;
        RECT 64.030 157.960 64.290 158.280 ;
        RECT 63.560 157.085 63.840 157.455 ;
        RECT 63.570 156.940 63.830 157.085 ;
        RECT 63.630 155.900 63.770 156.940 ;
        RECT 63.570 155.580 63.830 155.900 ;
        RECT 64.090 155.470 64.230 157.960 ;
        RECT 64.550 156.240 64.690 158.980 ;
        RECT 65.010 158.280 65.150 167.820 ;
        RECT 65.930 165.420 66.070 180.400 ;
        RECT 67.310 178.680 67.450 181.420 ;
        RECT 67.250 178.360 67.510 178.680 ;
        RECT 67.770 178.340 67.910 194.485 ;
        RECT 68.230 191.940 68.370 197.060 ;
        RECT 69.150 196.780 69.290 206.920 ;
        RECT 69.610 205.540 69.750 207.405 ;
        RECT 69.550 205.220 69.810 205.540 ;
        RECT 69.550 202.160 69.810 202.480 ;
        RECT 69.610 198.060 69.750 202.160 ;
        RECT 70.070 199.420 70.210 214.060 ;
        RECT 70.530 199.615 70.670 216.100 ;
        RECT 70.930 213.040 71.190 213.360 ;
        RECT 71.850 213.040 72.110 213.360 ;
        RECT 70.990 209.960 71.130 213.040 ;
        RECT 70.930 209.640 71.190 209.960 ;
        RECT 71.910 208.940 72.050 213.040 ;
        RECT 72.830 210.300 72.970 218.140 ;
        RECT 73.750 216.760 73.890 218.965 ;
        RECT 75.520 218.285 75.800 218.655 ;
        RECT 75.530 218.140 75.790 218.285 ;
        RECT 73.690 216.440 73.950 216.760 ;
        RECT 76.050 216.420 76.190 221.200 ;
        RECT 79.210 220.520 79.470 220.840 ;
        RECT 76.450 218.480 76.710 218.800 ;
        RECT 73.230 216.100 73.490 216.420 ;
        RECT 75.990 216.100 76.250 216.420 ;
        RECT 72.770 209.980 73.030 210.300 ;
        RECT 71.850 208.620 72.110 208.940 ;
        RECT 72.310 208.280 72.570 208.600 ;
        RECT 73.290 208.340 73.430 216.100 ;
        RECT 75.520 215.565 75.800 215.935 ;
        RECT 75.590 213.360 75.730 215.565 ;
        RECT 73.690 213.040 73.950 213.360 ;
        RECT 74.150 213.040 74.410 213.360 ;
        RECT 75.070 213.040 75.330 213.360 ;
        RECT 75.530 213.040 75.790 213.360 ;
        RECT 73.750 208.940 73.890 213.040 ;
        RECT 74.210 211.320 74.350 213.040 ;
        RECT 74.610 212.360 74.870 212.680 ;
        RECT 74.150 211.000 74.410 211.320 ;
        RECT 73.690 208.620 73.950 208.940 ;
        RECT 71.850 207.600 72.110 207.920 ;
        RECT 71.910 204.520 72.050 207.600 ;
        RECT 70.930 204.200 71.190 204.520 ;
        RECT 70.010 199.100 70.270 199.420 ;
        RECT 70.460 199.245 70.740 199.615 ;
        RECT 69.550 197.740 69.810 198.060 ;
        RECT 69.550 197.290 69.810 197.380 ;
        RECT 70.070 197.290 70.210 199.100 ;
        RECT 70.470 198.760 70.730 199.080 ;
        RECT 69.550 197.150 70.210 197.290 ;
        RECT 69.550 197.060 69.810 197.150 ;
        RECT 69.150 196.640 69.750 196.780 ;
        RECT 69.610 195.000 69.750 196.640 ;
        RECT 69.550 194.680 69.810 195.000 ;
        RECT 70.530 193.640 70.670 198.760 ;
        RECT 70.470 193.320 70.730 193.640 ;
        RECT 70.010 191.960 70.270 192.280 ;
        RECT 68.170 191.620 68.430 191.940 ;
        RECT 69.550 185.160 69.810 185.480 ;
        RECT 68.170 184.140 68.430 184.460 ;
        RECT 67.710 178.020 67.970 178.340 ;
        RECT 68.230 173.540 68.370 184.140 ;
        RECT 69.610 183.780 69.750 185.160 ;
        RECT 69.550 183.460 69.810 183.780 ;
        RECT 69.090 179.720 69.350 180.040 ;
        RECT 69.150 174.940 69.290 179.720 ;
        RECT 69.090 174.620 69.350 174.940 ;
        RECT 68.230 173.400 68.830 173.540 ;
        RECT 67.250 172.920 67.510 173.240 ;
        RECT 66.330 167.820 66.590 168.140 ;
        RECT 66.390 166.780 66.530 167.820 ;
        RECT 66.330 166.460 66.590 166.780 ;
        RECT 67.310 166.295 67.450 172.920 ;
        RECT 68.170 172.580 68.430 172.900 ;
        RECT 68.230 172.415 68.370 172.580 ;
        RECT 68.160 172.045 68.440 172.415 ;
        RECT 67.710 171.560 67.970 171.880 ;
        RECT 67.770 170.520 67.910 171.560 ;
        RECT 67.710 170.200 67.970 170.520 ;
        RECT 67.710 169.520 67.970 169.840 ;
        RECT 67.770 166.440 67.910 169.520 ;
        RECT 68.690 169.015 68.830 173.400 ;
        RECT 69.150 172.900 69.290 174.620 ;
        RECT 69.090 172.580 69.350 172.900 ;
        RECT 69.090 169.180 69.350 169.500 ;
        RECT 68.620 168.645 68.900 169.015 ;
        RECT 68.620 168.220 68.900 168.335 ;
        RECT 69.150 168.220 69.290 169.180 ;
        RECT 68.620 168.080 69.290 168.220 ;
        RECT 69.610 168.140 69.750 183.460 ;
        RECT 70.070 181.820 70.210 191.960 ;
        RECT 70.990 189.900 71.130 204.200 ;
        RECT 71.380 204.005 71.660 204.375 ;
        RECT 71.850 204.200 72.110 204.520 ;
        RECT 70.930 189.580 71.190 189.900 ;
        RECT 70.930 188.900 71.190 189.220 ;
        RECT 70.470 182.615 70.730 182.760 ;
        RECT 70.460 182.245 70.740 182.615 ;
        RECT 70.070 181.680 70.670 181.820 ;
        RECT 70.990 181.740 71.130 188.900 ;
        RECT 71.450 186.160 71.590 204.005 ;
        RECT 72.370 202.390 72.510 208.280 ;
        RECT 72.830 208.200 73.430 208.340 ;
        RECT 72.830 204.860 72.970 208.200 ;
        RECT 73.230 207.600 73.490 207.920 ;
        RECT 72.770 204.540 73.030 204.860 ;
        RECT 73.290 203.695 73.430 207.600 ;
        RECT 73.690 207.260 73.950 207.580 ;
        RECT 73.220 203.325 73.500 203.695 ;
        RECT 73.230 202.390 73.490 202.480 ;
        RECT 72.370 202.250 73.490 202.390 ;
        RECT 73.230 202.160 73.490 202.250 ;
        RECT 73.220 201.285 73.500 201.655 ;
        RECT 73.290 198.255 73.430 201.285 ;
        RECT 73.220 197.885 73.500 198.255 ;
        RECT 73.750 198.060 73.890 207.260 ;
        RECT 74.150 204.200 74.410 204.520 ;
        RECT 73.290 197.460 73.430 197.885 ;
        RECT 73.690 197.740 73.950 198.060 ;
        RECT 73.290 197.320 73.890 197.460 ;
        RECT 72.770 196.720 73.030 197.040 ;
        RECT 73.230 196.720 73.490 197.040 ;
        RECT 72.310 195.020 72.570 195.340 ;
        RECT 71.850 194.340 72.110 194.660 ;
        RECT 71.910 193.640 72.050 194.340 ;
        RECT 72.370 193.980 72.510 195.020 ;
        RECT 72.310 193.660 72.570 193.980 ;
        RECT 71.850 193.320 72.110 193.640 ;
        RECT 72.300 193.125 72.580 193.495 ;
        RECT 71.850 190.940 72.110 191.260 ;
        RECT 71.910 189.900 72.050 190.940 ;
        RECT 71.850 189.580 72.110 189.900 ;
        RECT 71.850 187.880 72.110 188.200 ;
        RECT 71.390 185.840 71.650 186.160 ;
        RECT 71.910 183.440 72.050 187.880 ;
        RECT 71.850 183.120 72.110 183.440 ;
        RECT 70.010 180.400 70.270 180.720 ;
        RECT 70.070 177.660 70.210 180.400 ;
        RECT 70.530 180.040 70.670 181.680 ;
        RECT 70.930 181.420 71.190 181.740 ;
        RECT 70.930 180.400 71.190 180.720 ;
        RECT 70.470 179.720 70.730 180.040 ;
        RECT 70.010 177.340 70.270 177.660 ;
        RECT 70.070 175.280 70.210 177.340 ;
        RECT 70.990 175.280 71.130 180.400 ;
        RECT 71.910 180.040 72.050 183.120 ;
        RECT 72.370 180.380 72.510 193.125 ;
        RECT 72.830 192.620 72.970 196.720 ;
        RECT 73.290 194.660 73.430 196.720 ;
        RECT 73.750 194.660 73.890 197.320 ;
        RECT 73.230 194.340 73.490 194.660 ;
        RECT 73.690 194.340 73.950 194.660 ;
        RECT 73.690 193.660 73.950 193.980 ;
        RECT 72.770 192.300 73.030 192.620 ;
        RECT 73.750 192.135 73.890 193.660 ;
        RECT 73.680 191.765 73.960 192.135 ;
        RECT 73.690 191.280 73.950 191.600 ;
        RECT 74.210 191.340 74.350 204.200 ;
        RECT 74.670 202.480 74.810 212.360 ;
        RECT 75.130 204.520 75.270 213.040 ;
        RECT 75.520 210.125 75.800 210.495 ;
        RECT 75.070 204.200 75.330 204.520 ;
        RECT 75.130 202.480 75.270 204.200 ;
        RECT 75.590 203.160 75.730 210.125 ;
        RECT 76.050 207.580 76.190 216.100 ;
        RECT 76.510 214.380 76.650 218.480 ;
        RECT 78.740 218.285 79.020 218.655 ;
        RECT 78.810 217.100 78.950 218.285 ;
        RECT 78.750 216.780 79.010 217.100 ;
        RECT 79.270 216.420 79.410 220.520 ;
        RECT 99.155 219.985 100.695 220.355 ;
        RECT 82.890 219.500 83.150 219.820 ;
        RECT 102.210 219.500 102.470 219.820 ;
        RECT 103.590 219.500 103.850 219.820 ;
        RECT 110.030 219.500 110.290 219.820 ;
        RECT 79.720 217.265 81.260 217.635 ;
        RECT 80.130 216.440 80.390 216.760 ;
        RECT 76.910 216.100 77.170 216.420 ;
        RECT 78.290 216.100 78.550 216.420 ;
        RECT 79.210 216.100 79.470 216.420 ;
        RECT 76.450 214.060 76.710 214.380 ;
        RECT 76.970 213.780 77.110 216.100 ;
        RECT 76.970 213.640 77.570 213.780 ;
        RECT 76.910 212.700 77.170 213.020 ;
        RECT 76.970 208.940 77.110 212.700 ;
        RECT 76.450 208.620 76.710 208.940 ;
        RECT 76.910 208.620 77.170 208.940 ;
        RECT 76.510 207.920 76.650 208.620 ;
        RECT 77.430 207.920 77.570 213.640 ;
        RECT 78.350 213.360 78.490 216.100 ;
        RECT 80.190 214.380 80.330 216.440 ;
        RECT 81.510 216.100 81.770 216.420 ;
        RECT 82.430 216.100 82.690 216.420 ;
        RECT 81.570 214.380 81.710 216.100 ;
        RECT 81.970 215.760 82.230 216.080 ;
        RECT 82.490 215.935 82.630 216.100 ;
        RECT 80.130 214.060 80.390 214.380 ;
        RECT 81.510 214.060 81.770 214.380 ;
        RECT 78.750 213.380 79.010 213.700 ;
        RECT 79.660 213.525 79.940 213.895 ;
        RECT 77.830 213.040 78.090 213.360 ;
        RECT 78.290 213.040 78.550 213.360 ;
        RECT 77.890 210.980 78.030 213.040 ;
        RECT 77.830 210.660 78.090 210.980 ;
        RECT 76.450 207.600 76.710 207.920 ;
        RECT 77.370 207.600 77.630 207.920 ;
        RECT 77.830 207.600 78.090 207.920 ;
        RECT 75.990 207.260 76.250 207.580 ;
        RECT 76.050 206.415 76.190 207.260 ;
        RECT 76.440 206.725 76.720 207.095 ;
        RECT 75.980 206.045 76.260 206.415 ;
        RECT 75.990 204.540 76.250 204.860 ;
        RECT 76.050 203.160 76.190 204.540 ;
        RECT 75.530 202.840 75.790 203.160 ;
        RECT 75.990 202.840 76.250 203.160 ;
        RECT 74.610 202.160 74.870 202.480 ;
        RECT 75.070 202.160 75.330 202.480 ;
        RECT 74.670 196.610 74.810 202.160 ;
        RECT 76.050 199.080 76.190 202.840 ;
        RECT 76.510 201.710 76.650 206.725 ;
        RECT 77.430 202.900 77.570 207.600 ;
        RECT 77.890 205.200 78.030 207.600 ;
        RECT 77.830 204.880 78.090 205.200 ;
        RECT 76.970 202.760 77.570 202.900 ;
        RECT 76.970 202.480 77.110 202.760 ;
        RECT 76.910 202.160 77.170 202.480 ;
        RECT 77.370 202.160 77.630 202.480 ;
        RECT 77.430 201.710 77.570 202.160 ;
        RECT 76.510 201.570 77.570 201.710 ;
        RECT 75.990 198.760 76.250 199.080 ;
        RECT 77.430 198.820 77.570 201.570 ;
        RECT 76.050 197.040 76.190 198.760 ;
        RECT 76.970 198.680 77.570 198.820 ;
        RECT 76.440 197.885 76.720 198.255 ;
        RECT 76.510 197.040 76.650 197.885 ;
        RECT 75.990 196.720 76.250 197.040 ;
        RECT 76.450 196.720 76.710 197.040 ;
        RECT 75.070 196.610 75.330 196.700 ;
        RECT 74.670 196.470 75.330 196.610 ;
        RECT 74.670 194.660 74.810 196.470 ;
        RECT 75.070 196.380 75.330 196.470 ;
        RECT 74.610 194.340 74.870 194.660 ;
        RECT 74.610 193.660 74.870 193.980 ;
        RECT 74.670 192.620 74.810 193.660 ;
        RECT 74.610 192.300 74.870 192.620 ;
        RECT 76.970 192.280 77.110 198.680 ;
        RECT 77.370 197.740 77.630 198.060 ;
        RECT 76.910 191.960 77.170 192.280 ;
        RECT 74.600 191.340 74.880 191.455 ;
        RECT 73.230 188.900 73.490 189.220 ;
        RECT 72.770 183.800 73.030 184.120 ;
        RECT 72.310 180.060 72.570 180.380 ;
        RECT 71.850 179.720 72.110 180.040 ;
        RECT 71.910 178.340 72.050 179.720 ;
        RECT 71.850 178.020 72.110 178.340 ;
        RECT 70.010 174.960 70.270 175.280 ;
        RECT 70.930 174.960 71.190 175.280 ;
        RECT 70.070 172.560 70.210 174.960 ;
        RECT 70.470 172.580 70.730 172.900 ;
        RECT 70.010 172.240 70.270 172.560 ;
        RECT 68.620 167.965 68.900 168.080 ;
        RECT 67.240 165.925 67.520 166.295 ;
        RECT 67.710 166.120 67.970 166.440 ;
        RECT 67.770 165.420 67.910 166.120 ;
        RECT 65.870 165.100 66.130 165.420 ;
        RECT 67.710 165.100 67.970 165.420 ;
        RECT 68.630 165.100 68.890 165.420 ;
        RECT 66.330 164.420 66.590 164.740 ;
        RECT 66.780 164.565 67.060 164.935 ;
        RECT 65.860 163.205 66.140 163.575 ;
        RECT 65.410 159.320 65.670 159.640 ;
        RECT 64.950 157.960 65.210 158.280 ;
        RECT 65.470 156.580 65.610 159.320 ;
        RECT 65.930 158.620 66.070 163.205 ;
        RECT 66.390 158.870 66.530 164.420 ;
        RECT 66.850 159.210 66.990 164.565 ;
        RECT 67.710 163.740 67.970 164.060 ;
        RECT 67.770 162.215 67.910 163.740 ;
        RECT 68.160 163.205 68.440 163.575 ;
        RECT 67.700 161.845 67.980 162.215 ;
        RECT 68.230 159.980 68.370 163.205 ;
        RECT 68.690 161.680 68.830 165.100 ;
        RECT 69.150 162.360 69.290 168.080 ;
        RECT 69.550 167.820 69.810 168.140 ;
        RECT 70.530 167.800 70.670 172.580 ;
        RECT 70.990 171.880 71.130 174.960 ;
        RECT 72.310 174.620 72.570 174.940 ;
        RECT 71.390 174.280 71.650 174.600 ;
        RECT 70.930 171.560 71.190 171.880 ;
        RECT 70.990 170.180 71.130 171.560 ;
        RECT 70.930 169.860 71.190 170.180 ;
        RECT 71.450 167.800 71.590 174.280 ;
        RECT 72.370 173.095 72.510 174.620 ;
        RECT 72.300 172.725 72.580 173.095 ;
        RECT 70.470 167.480 70.730 167.800 ;
        RECT 71.390 167.480 71.650 167.800 ;
        RECT 72.310 166.800 72.570 167.120 ;
        RECT 72.370 165.080 72.510 166.800 ;
        RECT 72.310 164.760 72.570 165.080 ;
        RECT 69.090 162.100 69.350 162.360 ;
        RECT 69.090 162.040 70.670 162.100 ;
        RECT 69.150 162.020 70.670 162.040 ;
        RECT 69.150 161.960 70.730 162.020 ;
        RECT 70.470 161.700 70.730 161.960 ;
        RECT 68.630 161.360 68.890 161.680 ;
        RECT 68.690 159.980 68.830 161.360 ;
        RECT 68.170 159.660 68.430 159.980 ;
        RECT 68.630 159.660 68.890 159.980 ;
        RECT 70.010 159.210 70.270 159.300 ;
        RECT 66.850 159.070 70.270 159.210 ;
        RECT 70.010 158.980 70.270 159.070 ;
        RECT 66.390 158.730 67.910 158.870 ;
        RECT 65.870 158.300 66.130 158.620 ;
        RECT 64.950 156.260 65.210 156.580 ;
        RECT 65.410 156.260 65.670 156.580 ;
        RECT 64.490 155.920 64.750 156.240 ;
        RECT 64.090 155.330 64.690 155.470 ;
        RECT 57.590 154.220 57.850 154.540 ;
        RECT 58.570 154.480 59.630 154.620 ;
        RECT 57.580 152.325 57.860 152.695 ;
        RECT 57.130 148.100 57.390 148.420 ;
        RECT 57.130 147.080 57.390 147.400 ;
        RECT 57.190 146.380 57.330 147.080 ;
        RECT 57.130 146.060 57.390 146.380 ;
        RECT 56.670 145.040 56.930 145.360 ;
        RECT 57.650 145.100 57.790 152.325 ;
        RECT 59.490 150.800 59.630 154.480 ;
        RECT 61.730 154.220 61.990 154.540 ;
        RECT 63.170 154.480 64.230 154.620 ;
        RECT 59.890 153.540 60.150 153.860 ;
        RECT 60.350 153.540 60.610 153.860 ;
        RECT 58.970 150.480 59.230 150.800 ;
        RECT 59.430 150.480 59.690 150.800 ;
        RECT 58.050 148.780 58.310 149.100 ;
        RECT 58.110 147.935 58.250 148.780 ;
        RECT 58.510 148.440 58.770 148.760 ;
        RECT 58.040 147.565 58.320 147.935 ;
        RECT 58.110 146.380 58.250 147.565 ;
        RECT 58.050 146.060 58.310 146.380 ;
        RECT 58.570 145.360 58.710 148.440 ;
        RECT 59.030 146.380 59.170 150.480 ;
        RECT 59.950 150.120 60.090 153.540 ;
        RECT 60.410 151.820 60.550 153.540 ;
        RECT 61.790 153.090 61.930 154.220 ;
        RECT 63.570 153.090 63.830 153.180 ;
        RECT 61.790 152.950 63.830 153.090 ;
        RECT 63.570 152.860 63.830 152.950 ;
        RECT 60.350 151.500 60.610 151.820 ;
        RECT 63.110 150.480 63.370 150.800 ;
        RECT 59.890 149.800 60.150 150.120 ;
        RECT 60.285 149.265 61.825 149.635 ;
        RECT 62.190 148.100 62.450 148.420 ;
        RECT 62.250 146.380 62.390 148.100 ;
        RECT 58.970 146.060 59.230 146.380 ;
        RECT 59.890 146.060 60.150 146.380 ;
        RECT 62.190 146.060 62.450 146.380 ;
        RECT 58.960 145.525 59.240 145.895 ;
        RECT 57.650 144.960 58.250 145.100 ;
        RECT 58.510 145.040 58.770 145.360 ;
        RECT 57.130 144.360 57.390 144.680 ;
        RECT 57.590 144.360 57.850 144.680 ;
        RECT 56.200 143.485 56.480 143.855 ;
        RECT 56.270 142.980 56.410 143.485 ;
        RECT 56.210 142.660 56.470 142.980 ;
        RECT 56.670 141.980 56.930 142.300 ;
        RECT 56.730 139.920 56.870 141.980 ;
        RECT 56.670 139.600 56.930 139.920 ;
        RECT 56.730 139.095 56.870 139.600 ;
        RECT 56.660 138.725 56.940 139.095 ;
        RECT 55.750 136.200 56.010 136.520 ;
        RECT 54.830 135.180 55.090 135.500 ;
        RECT 53.910 134.500 54.170 134.820 ;
        RECT 54.830 134.500 55.090 134.820 ;
        RECT 56.210 134.500 56.470 134.820 ;
        RECT 54.890 132.780 55.030 134.500 ;
        RECT 54.830 132.460 55.090 132.780 ;
        RECT 52.990 131.780 53.250 132.100 ;
        RECT 52.530 131.100 52.790 131.420 ;
        RECT 52.070 130.760 52.330 131.080 ;
        RECT 52.130 129.040 52.270 130.760 ;
        RECT 52.070 128.720 52.330 129.040 ;
        RECT 52.130 125.980 52.270 128.720 ;
        RECT 52.070 125.660 52.330 125.980 ;
        RECT 51.610 125.320 51.870 125.640 ;
        RECT 53.050 125.550 53.190 131.780 ;
        RECT 56.270 129.380 56.410 134.500 ;
        RECT 57.190 130.060 57.330 144.360 ;
        RECT 57.650 143.660 57.790 144.360 ;
        RECT 57.590 143.340 57.850 143.660 ;
        RECT 57.650 137.540 57.790 143.340 ;
        RECT 58.110 140.455 58.250 144.960 ;
        RECT 58.040 140.085 58.320 140.455 ;
        RECT 57.590 137.220 57.850 137.540 ;
        RECT 57.650 132.100 57.790 137.220 ;
        RECT 59.030 136.860 59.170 145.525 ;
        RECT 59.950 143.660 60.090 146.060 ;
        RECT 62.650 145.380 62.910 145.700 ;
        RECT 62.190 145.040 62.450 145.360 ;
        RECT 60.285 143.825 61.825 144.195 ;
        RECT 62.250 143.855 62.390 145.040 ;
        RECT 59.890 143.340 60.150 143.660 ;
        RECT 62.180 143.485 62.460 143.855 ;
        RECT 59.430 143.000 59.690 143.320 ;
        RECT 58.970 136.540 59.230 136.860 ;
        RECT 57.590 131.780 57.850 132.100 ;
        RECT 57.130 129.740 57.390 130.060 ;
        RECT 55.750 129.060 56.010 129.380 ;
        RECT 56.210 129.060 56.470 129.380 ;
        RECT 55.810 127.340 55.950 129.060 ;
        RECT 57.130 128.040 57.390 128.360 ;
        RECT 55.750 127.020 56.010 127.340 ;
        RECT 57.190 127.000 57.330 128.040 ;
        RECT 57.130 126.680 57.390 127.000 ;
        RECT 57.650 126.660 57.790 131.780 ;
        RECT 58.050 131.100 58.310 131.420 ;
        RECT 58.110 129.040 58.250 131.100 ;
        RECT 58.050 128.720 58.310 129.040 ;
        RECT 59.030 127.000 59.170 136.540 ;
        RECT 59.490 135.500 59.630 143.000 ;
        RECT 60.285 138.385 61.825 138.755 ;
        RECT 62.710 137.540 62.850 145.380 ;
        RECT 63.170 144.680 63.310 150.480 ;
        RECT 63.110 144.360 63.370 144.680 ;
        RECT 63.110 142.210 63.370 142.300 ;
        RECT 63.630 142.210 63.770 152.860 ;
        RECT 64.090 152.840 64.230 154.480 ;
        RECT 64.550 153.180 64.690 155.330 ;
        RECT 65.010 153.860 65.150 156.260 ;
        RECT 67.770 156.240 67.910 158.730 ;
        RECT 69.090 158.300 69.350 158.620 ;
        RECT 67.250 155.920 67.510 156.240 ;
        RECT 67.710 155.920 67.970 156.240 ;
        RECT 65.410 155.580 65.670 155.900 ;
        RECT 65.470 153.860 65.610 155.580 ;
        RECT 66.330 154.220 66.590 154.540 ;
        RECT 64.950 153.540 65.210 153.860 ;
        RECT 65.410 153.540 65.670 153.860 ;
        RECT 64.490 152.860 64.750 153.180 ;
        RECT 64.030 152.520 64.290 152.840 ;
        RECT 64.090 151.480 64.230 152.520 ;
        RECT 64.030 151.160 64.290 151.480 ;
        RECT 64.550 148.330 64.690 152.860 ;
        RECT 65.010 151.820 65.150 153.540 ;
        RECT 66.390 153.090 66.530 154.220 ;
        RECT 67.310 154.200 67.450 155.920 ;
        RECT 67.250 153.880 67.510 154.200 ;
        RECT 66.790 153.200 67.050 153.520 ;
        RECT 65.470 152.950 66.530 153.090 ;
        RECT 64.950 151.500 65.210 151.820 ;
        RECT 64.950 150.820 65.210 151.140 ;
        RECT 64.090 148.190 64.690 148.330 ;
        RECT 64.090 145.895 64.230 148.190 ;
        RECT 64.490 147.420 64.750 147.740 ;
        RECT 64.020 145.525 64.300 145.895 ;
        RECT 64.550 145.360 64.690 147.420 ;
        RECT 64.030 145.040 64.290 145.360 ;
        RECT 64.490 145.040 64.750 145.360 ;
        RECT 63.110 142.070 63.770 142.210 ;
        RECT 63.110 141.980 63.370 142.070 ;
        RECT 62.650 137.220 62.910 137.540 ;
        RECT 59.430 135.180 59.690 135.500 ;
        RECT 63.170 134.820 63.310 141.980 ;
        RECT 64.090 139.580 64.230 145.040 ;
        RECT 64.550 140.600 64.690 145.040 ;
        RECT 65.010 144.535 65.150 150.820 ;
        RECT 64.940 144.165 65.220 144.535 ;
        RECT 64.950 143.570 65.210 143.660 ;
        RECT 65.470 143.570 65.610 152.950 ;
        RECT 65.870 151.500 66.130 151.820 ;
        RECT 64.950 143.430 65.610 143.570 ;
        RECT 64.950 143.340 65.210 143.430 ;
        RECT 64.490 140.280 64.750 140.600 ;
        RECT 64.030 139.260 64.290 139.580 ;
        RECT 64.550 137.200 64.690 140.280 ;
        RECT 65.010 140.260 65.150 143.340 ;
        RECT 65.410 142.320 65.670 142.640 ;
        RECT 64.950 139.940 65.210 140.260 ;
        RECT 64.490 136.880 64.750 137.200 ;
        RECT 64.550 136.375 64.690 136.880 ;
        RECT 64.940 136.685 65.220 137.055 ;
        RECT 64.480 136.005 64.760 136.375 ;
        RECT 63.110 134.500 63.370 134.820 ;
        RECT 60.285 132.945 61.825 133.315 ;
        RECT 59.890 129.740 60.150 130.060 ;
        RECT 58.970 126.680 59.230 127.000 ;
        RECT 57.590 126.340 57.850 126.660 ;
        RECT 59.950 126.320 60.090 129.740 ;
        RECT 63.170 129.720 63.310 134.500 ;
        RECT 65.010 134.140 65.150 136.685 ;
        RECT 65.470 134.140 65.610 142.320 ;
        RECT 65.930 134.140 66.070 151.500 ;
        RECT 66.850 151.140 66.990 153.200 ;
        RECT 68.170 152.520 68.430 152.840 ;
        RECT 68.230 151.220 68.370 152.520 ;
        RECT 66.790 150.820 67.050 151.140 ;
        RECT 68.230 151.080 68.830 151.220 ;
        RECT 67.250 149.800 67.510 150.120 ;
        RECT 66.790 148.440 67.050 148.760 ;
        RECT 66.850 147.740 66.990 148.440 ;
        RECT 67.310 148.420 67.450 149.800 ;
        RECT 67.250 148.100 67.510 148.420 ;
        RECT 66.790 147.420 67.050 147.740 ;
        RECT 67.310 146.380 67.450 148.100 ;
        RECT 67.250 146.060 67.510 146.380 ;
        RECT 68.170 146.060 68.430 146.380 ;
        RECT 67.310 145.100 67.450 146.060 ;
        RECT 68.230 145.215 68.370 146.060 ;
        RECT 66.850 144.960 67.450 145.100 ;
        RECT 66.850 142.980 66.990 144.960 ;
        RECT 68.160 144.845 68.440 145.215 ;
        RECT 67.250 144.360 67.510 144.680 ;
        RECT 66.790 142.660 67.050 142.980 ;
        RECT 67.310 141.135 67.450 144.360 ;
        RECT 67.700 143.060 67.980 143.175 ;
        RECT 68.690 143.060 68.830 151.080 ;
        RECT 69.150 148.420 69.290 158.300 ;
        RECT 70.530 156.920 70.670 161.700 ;
        RECT 72.370 161.680 72.510 164.760 ;
        RECT 72.310 161.360 72.570 161.680 ;
        RECT 72.830 159.495 72.970 183.800 ;
        RECT 73.290 183.780 73.430 188.900 ;
        RECT 73.750 188.735 73.890 191.280 ;
        RECT 74.210 191.200 74.880 191.340 ;
        RECT 76.450 191.280 76.710 191.600 ;
        RECT 74.600 191.085 74.880 191.200 ;
        RECT 74.150 188.900 74.410 189.220 ;
        RECT 73.680 188.365 73.960 188.735 ;
        RECT 73.690 185.160 73.950 185.480 ;
        RECT 73.230 183.460 73.490 183.780 ;
        RECT 73.290 181.740 73.430 183.460 ;
        RECT 73.230 181.420 73.490 181.740 ;
        RECT 73.750 181.140 73.890 185.160 ;
        RECT 74.210 184.120 74.350 188.900 ;
        RECT 74.150 183.800 74.410 184.120 ;
        RECT 73.290 181.000 73.890 181.140 ;
        RECT 73.290 173.580 73.430 181.000 ;
        RECT 73.680 177.485 73.960 177.855 ;
        RECT 74.670 177.660 74.810 191.085 ;
        RECT 76.510 186.500 76.650 191.280 ;
        RECT 76.450 186.180 76.710 186.500 ;
        RECT 77.430 185.480 77.570 197.740 ;
        RECT 77.890 195.340 78.030 204.880 ;
        RECT 78.290 202.160 78.550 202.480 ;
        RECT 78.350 200.295 78.490 202.160 ;
        RECT 78.280 199.925 78.560 200.295 ;
        RECT 77.830 195.020 78.090 195.340 ;
        RECT 78.350 189.300 78.490 199.925 ;
        RECT 78.810 197.460 78.950 213.380 ;
        RECT 79.730 213.360 79.870 213.525 ;
        RECT 79.670 213.040 79.930 213.360 ;
        RECT 82.030 212.420 82.170 215.760 ;
        RECT 82.420 215.565 82.700 215.935 ;
        RECT 82.950 214.040 83.090 219.500 ;
        RECT 101.290 219.160 101.550 219.480 ;
        RECT 95.310 218.480 95.570 218.800 ;
        RECT 95.770 218.655 96.030 218.800 ;
        RECT 83.350 217.800 83.610 218.120 ;
        RECT 83.410 216.760 83.550 217.800 ;
        RECT 92.540 217.605 92.820 217.975 ;
        RECT 92.610 217.100 92.750 217.605 ;
        RECT 95.370 217.100 95.510 218.480 ;
        RECT 95.760 218.285 96.040 218.655 ;
        RECT 97.610 218.480 97.870 218.800 ;
        RECT 92.550 216.780 92.810 217.100 ;
        RECT 95.310 217.010 95.570 217.100 ;
        RECT 94.910 216.870 95.570 217.010 ;
        RECT 83.350 216.440 83.610 216.760 ;
        RECT 89.790 216.440 90.050 216.760 ;
        RECT 86.570 215.080 86.830 215.400 ;
        RECT 82.890 213.780 83.150 214.040 ;
        RECT 82.890 213.720 84.010 213.780 ;
        RECT 82.950 213.640 84.010 213.720 ;
        RECT 82.430 213.040 82.690 213.360 ;
        RECT 81.570 212.280 82.170 212.420 ;
        RECT 79.720 211.825 81.260 212.195 ;
        RECT 79.720 206.385 81.260 206.755 ;
        RECT 79.210 203.180 79.470 203.500 ;
        RECT 79.270 202.900 79.410 203.180 ;
        RECT 79.270 202.820 80.790 202.900 ;
        RECT 79.270 202.760 80.850 202.820 ;
        RECT 79.270 198.060 79.410 202.760 ;
        RECT 80.590 202.500 80.850 202.760 ;
        RECT 80.130 202.160 80.390 202.480 ;
        RECT 80.190 201.800 80.330 202.160 ;
        RECT 80.130 201.480 80.390 201.800 ;
        RECT 79.720 200.945 81.260 201.315 ;
        RECT 81.050 199.440 81.310 199.760 ;
        RECT 79.210 197.740 79.470 198.060 ;
        RECT 78.810 197.320 79.410 197.460 ;
        RECT 78.750 196.720 79.010 197.040 ;
        RECT 78.810 191.940 78.950 196.720 ;
        RECT 78.750 191.620 79.010 191.940 ;
        RECT 78.740 189.300 79.020 189.415 ;
        RECT 78.350 189.160 79.020 189.300 ;
        RECT 78.740 189.045 79.020 189.160 ;
        RECT 78.750 187.880 79.010 188.200 ;
        RECT 78.810 186.160 78.950 187.880 ;
        RECT 78.290 185.840 78.550 186.160 ;
        RECT 78.750 185.840 79.010 186.160 ;
        RECT 77.370 185.160 77.630 185.480 ;
        RECT 77.370 184.140 77.630 184.460 ;
        RECT 78.350 184.370 78.490 185.840 ;
        RECT 78.350 184.230 78.950 184.370 ;
        RECT 76.910 183.800 77.170 184.120 ;
        RECT 75.070 183.460 75.330 183.780 ;
        RECT 75.130 180.720 75.270 183.460 ;
        RECT 76.970 181.060 77.110 183.800 ;
        RECT 77.430 183.780 77.570 184.140 ;
        RECT 77.370 183.460 77.630 183.780 ;
        RECT 78.290 183.460 78.550 183.780 ;
        RECT 78.350 181.740 78.490 183.460 ;
        RECT 78.290 181.420 78.550 181.740 ;
        RECT 76.910 180.740 77.170 181.060 ;
        RECT 75.070 180.400 75.330 180.720 ;
        RECT 75.130 178.340 75.270 180.400 ;
        RECT 75.990 180.060 76.250 180.380 ;
        RECT 75.070 178.020 75.330 178.340 ;
        RECT 75.530 178.020 75.790 178.340 ;
        RECT 73.230 173.260 73.490 173.580 ;
        RECT 73.750 172.220 73.890 177.485 ;
        RECT 74.610 177.340 74.870 177.660 ;
        RECT 75.590 176.300 75.730 178.020 ;
        RECT 76.050 176.300 76.190 180.060 ;
        RECT 76.970 178.340 77.110 180.740 ;
        RECT 78.350 180.720 78.490 181.420 ;
        RECT 78.290 180.400 78.550 180.720 ;
        RECT 77.370 180.060 77.630 180.380 ;
        RECT 77.430 178.340 77.570 180.060 ;
        RECT 78.290 179.720 78.550 180.040 ;
        RECT 77.830 178.360 78.090 178.680 ;
        RECT 76.910 178.020 77.170 178.340 ;
        RECT 77.370 178.020 77.630 178.340 ;
        RECT 75.530 175.980 75.790 176.300 ;
        RECT 75.990 175.980 76.250 176.300 ;
        RECT 75.990 175.190 76.250 175.280 ;
        RECT 75.590 175.050 76.250 175.190 ;
        RECT 74.610 174.620 74.870 174.940 ;
        RECT 73.690 171.900 73.950 172.220 ;
        RECT 74.670 170.860 74.810 174.620 ;
        RECT 75.070 172.920 75.330 173.240 ;
        RECT 75.130 171.735 75.270 172.920 ;
        RECT 75.060 171.365 75.340 171.735 ;
        RECT 74.610 170.540 74.870 170.860 ;
        RECT 75.060 170.685 75.340 171.055 ;
        RECT 74.150 167.140 74.410 167.460 ;
        RECT 73.230 166.460 73.490 166.780 ;
        RECT 73.290 162.700 73.430 166.460 ;
        RECT 73.690 164.420 73.950 164.740 ;
        RECT 73.230 162.380 73.490 162.700 ;
        RECT 73.750 161.680 73.890 164.420 ;
        RECT 74.210 164.400 74.350 167.140 ;
        RECT 74.610 166.975 74.870 167.120 ;
        RECT 74.600 166.605 74.880 166.975 ;
        RECT 75.130 166.780 75.270 170.685 ;
        RECT 75.070 166.460 75.330 166.780 ;
        RECT 75.590 165.420 75.730 175.050 ;
        RECT 75.990 174.960 76.250 175.050 ;
        RECT 77.370 174.850 77.630 174.940 ;
        RECT 76.510 174.710 77.630 174.850 ;
        RECT 75.990 174.280 76.250 174.600 ;
        RECT 76.050 173.775 76.190 174.280 ;
        RECT 75.980 173.405 76.260 173.775 ;
        RECT 76.510 172.900 76.650 174.710 ;
        RECT 77.370 174.620 77.630 174.710 ;
        RECT 77.370 173.260 77.630 173.580 ;
        RECT 76.450 172.580 76.710 172.900 ;
        RECT 76.510 169.840 76.650 172.580 ;
        RECT 76.450 169.520 76.710 169.840 ;
        RECT 76.910 168.840 77.170 169.160 ;
        RECT 75.990 166.460 76.250 166.780 ;
        RECT 75.530 165.100 75.790 165.420 ;
        RECT 74.150 164.080 74.410 164.400 ;
        RECT 74.210 162.700 74.350 164.080 ;
        RECT 74.610 163.400 74.870 163.720 ;
        RECT 74.670 162.895 74.810 163.400 ;
        RECT 74.150 162.380 74.410 162.700 ;
        RECT 74.600 162.525 74.880 162.895 ;
        RECT 76.050 162.700 76.190 166.460 ;
        RECT 76.970 165.615 77.110 168.840 ;
        RECT 77.430 168.140 77.570 173.260 ;
        RECT 77.890 170.860 78.030 178.360 ;
        RECT 77.830 170.540 78.090 170.860 ;
        RECT 77.830 169.180 78.090 169.500 ;
        RECT 77.890 168.140 78.030 169.180 ;
        RECT 77.370 167.820 77.630 168.140 ;
        RECT 77.830 167.820 78.090 168.140 ;
        RECT 78.350 167.655 78.490 179.720 ;
        RECT 78.810 177.660 78.950 184.230 ;
        RECT 79.270 178.340 79.410 197.320 ;
        RECT 81.110 196.780 81.250 199.440 ;
        RECT 81.570 197.380 81.710 212.280 ;
        RECT 82.490 211.660 82.630 213.040 ;
        RECT 82.890 212.360 83.150 212.680 ;
        RECT 82.430 211.570 82.690 211.660 ;
        RECT 82.030 211.430 82.690 211.570 ;
        RECT 82.030 209.960 82.170 211.430 ;
        RECT 82.430 211.340 82.690 211.430 ;
        RECT 82.430 210.320 82.690 210.640 ;
        RECT 81.970 209.640 82.230 209.960 ;
        RECT 82.490 208.940 82.630 210.320 ;
        RECT 82.430 208.620 82.690 208.940 ;
        RECT 82.950 208.455 83.090 212.360 ;
        RECT 81.970 208.170 82.230 208.260 ;
        RECT 81.970 208.030 82.630 208.170 ;
        RECT 82.880 208.085 83.160 208.455 ;
        RECT 81.970 207.940 82.230 208.030 ;
        RECT 81.970 207.260 82.230 207.580 ;
        RECT 82.030 203.015 82.170 207.260 ;
        RECT 81.960 202.645 82.240 203.015 ;
        RECT 82.490 202.900 82.630 208.030 ;
        RECT 82.890 207.830 83.150 207.920 ;
        RECT 82.890 207.690 83.550 207.830 ;
        RECT 82.890 207.600 83.150 207.690 ;
        RECT 82.890 206.920 83.150 207.240 ;
        RECT 82.950 205.200 83.090 206.920 ;
        RECT 83.410 206.415 83.550 207.690 ;
        RECT 83.870 207.095 84.010 213.640 ;
        RECT 86.630 213.360 86.770 215.080 ;
        RECT 89.850 214.380 89.990 216.440 ;
        RECT 91.170 216.100 91.430 216.420 ;
        RECT 91.630 216.100 91.890 216.420 ;
        RECT 91.230 214.380 91.370 216.100 ;
        RECT 89.790 214.290 90.050 214.380 ;
        RECT 89.790 214.150 90.450 214.290 ;
        RECT 89.790 214.060 90.050 214.150 ;
        RECT 84.730 213.215 84.990 213.360 ;
        RECT 84.720 212.845 85.000 213.215 ;
        RECT 85.190 213.040 85.450 213.360 ;
        RECT 86.570 213.040 86.830 213.360 ;
        RECT 87.950 213.040 88.210 213.360 ;
        RECT 84.730 212.360 84.990 212.680 ;
        RECT 84.790 207.920 84.930 212.360 ;
        RECT 85.250 210.980 85.390 213.040 ;
        RECT 86.630 211.320 86.770 213.040 ;
        RECT 87.490 212.360 87.750 212.680 ;
        RECT 86.570 211.000 86.830 211.320 ;
        RECT 85.190 210.660 85.450 210.980 ;
        RECT 84.270 207.600 84.530 207.920 ;
        RECT 84.730 207.600 84.990 207.920 ;
        RECT 83.800 206.725 84.080 207.095 ;
        RECT 83.340 206.045 83.620 206.415 ;
        RECT 83.350 205.560 83.610 205.880 ;
        RECT 82.890 204.880 83.150 205.200 ;
        RECT 83.410 203.695 83.550 205.560 ;
        RECT 83.870 204.260 84.010 206.725 ;
        RECT 84.330 204.860 84.470 207.600 ;
        RECT 85.250 205.620 85.390 210.660 ;
        RECT 86.100 208.765 86.380 209.135 ;
        RECT 85.650 207.940 85.910 208.260 ;
        RECT 85.710 206.220 85.850 207.940 ;
        RECT 86.170 207.920 86.310 208.765 ;
        RECT 86.110 207.775 86.370 207.920 ;
        RECT 86.100 207.405 86.380 207.775 ;
        RECT 85.650 205.900 85.910 206.220 ;
        RECT 86.100 206.045 86.380 206.415 ;
        RECT 86.110 205.900 86.370 206.045 ;
        RECT 84.730 205.220 84.990 205.540 ;
        RECT 85.250 205.480 85.850 205.620 ;
        RECT 84.270 204.540 84.530 204.860 ;
        RECT 84.260 204.260 84.540 204.375 ;
        RECT 84.790 204.260 84.930 205.220 ;
        RECT 83.870 204.120 84.930 204.260 ;
        RECT 84.260 204.005 84.540 204.120 ;
        RECT 83.340 203.325 83.620 203.695 ;
        RECT 85.190 203.180 85.450 203.500 ;
        RECT 82.490 202.760 83.550 202.900 ;
        RECT 82.030 199.670 82.170 202.645 ;
        RECT 82.430 201.480 82.690 201.800 ;
        RECT 82.890 201.655 83.150 201.800 ;
        RECT 82.490 200.180 82.630 201.480 ;
        RECT 82.880 201.285 83.160 201.655 ;
        RECT 82.880 200.605 83.160 200.975 ;
        RECT 82.890 200.460 83.150 200.605 ;
        RECT 82.490 200.040 83.090 200.180 ;
        RECT 83.410 200.100 83.550 202.760 ;
        RECT 84.270 202.160 84.530 202.480 ;
        RECT 84.730 202.160 84.990 202.480 ;
        RECT 83.810 201.820 84.070 202.140 ;
        RECT 83.870 200.295 84.010 201.820 ;
        RECT 82.030 199.530 82.630 199.670 ;
        RECT 81.510 197.060 81.770 197.380 ;
        RECT 81.110 196.640 81.710 196.780 ;
        RECT 81.970 196.720 82.230 197.040 ;
        RECT 79.720 195.505 81.260 195.875 ;
        RECT 81.570 193.980 81.710 196.640 ;
        RECT 82.030 194.660 82.170 196.720 ;
        RECT 82.490 196.700 82.630 199.530 ;
        RECT 82.430 196.380 82.690 196.700 ;
        RECT 82.420 195.165 82.700 195.535 ;
        RECT 81.970 194.340 82.230 194.660 ;
        RECT 82.490 194.060 82.630 195.165 ;
        RECT 82.950 195.000 83.090 200.040 ;
        RECT 83.350 199.780 83.610 200.100 ;
        RECT 83.800 199.925 84.080 200.295 ;
        RECT 84.330 199.670 84.470 202.160 ;
        RECT 84.790 200.780 84.930 202.160 ;
        RECT 84.730 200.460 84.990 200.780 ;
        RECT 84.330 199.530 84.930 199.670 ;
        RECT 84.790 198.060 84.930 199.530 ;
        RECT 84.730 197.740 84.990 198.060 ;
        RECT 85.250 197.290 85.390 203.180 ;
        RECT 85.710 202.390 85.850 205.480 ;
        RECT 86.110 205.220 86.370 205.540 ;
        RECT 86.170 203.500 86.310 205.220 ;
        RECT 86.110 203.180 86.370 203.500 ;
        RECT 86.110 202.390 86.370 202.480 ;
        RECT 85.710 202.250 86.370 202.390 ;
        RECT 86.110 202.160 86.370 202.250 ;
        RECT 86.110 201.710 86.370 201.800 ;
        RECT 85.710 201.570 86.370 201.710 ;
        RECT 85.710 198.255 85.850 201.570 ;
        RECT 86.110 201.480 86.370 201.570 ;
        RECT 86.630 200.100 86.770 211.000 ;
        RECT 87.550 210.980 87.690 212.360 ;
        RECT 87.490 210.660 87.750 210.980 ;
        RECT 87.490 209.980 87.750 210.300 ;
        RECT 87.030 209.640 87.290 209.960 ;
        RECT 86.570 199.780 86.830 200.100 ;
        RECT 85.640 197.885 85.920 198.255 ;
        RECT 84.790 197.150 85.390 197.290 ;
        RECT 86.100 197.205 86.380 197.575 ;
        RECT 84.790 195.420 84.930 197.150 ;
        RECT 85.650 196.720 85.910 197.040 ;
        RECT 84.790 195.280 85.390 195.420 ;
        RECT 82.890 194.855 83.150 195.000 ;
        RECT 82.880 194.485 83.160 194.855 ;
        RECT 81.510 193.660 81.770 193.980 ;
        RECT 82.030 193.920 82.630 194.060 ;
        RECT 83.350 194.000 83.610 194.320 ;
        RECT 84.270 194.000 84.530 194.320 ;
        RECT 81.510 192.300 81.770 192.620 ;
        RECT 79.720 190.065 81.260 190.435 ;
        RECT 81.570 189.900 81.710 192.300 ;
        RECT 82.030 192.280 82.170 193.920 ;
        RECT 83.410 193.495 83.550 194.000 ;
        RECT 83.340 193.125 83.620 193.495 ;
        RECT 83.810 193.320 84.070 193.640 ;
        RECT 81.970 191.960 82.230 192.280 ;
        RECT 81.510 189.580 81.770 189.900 ;
        RECT 81.050 189.240 81.310 189.560 ;
        RECT 80.130 188.900 80.390 189.220 ;
        RECT 80.190 186.160 80.330 188.900 ;
        RECT 81.110 187.180 81.250 189.240 ;
        RECT 81.050 186.860 81.310 187.180 ;
        RECT 80.130 185.840 80.390 186.160 ;
        RECT 81.510 185.840 81.770 186.160 ;
        RECT 79.720 184.625 81.260 184.995 ;
        RECT 81.570 184.460 81.710 185.840 ;
        RECT 81.510 184.140 81.770 184.460 ;
        RECT 82.030 182.760 82.170 191.960 ;
        RECT 82.430 189.580 82.690 189.900 ;
        RECT 82.490 189.220 82.630 189.580 ;
        RECT 82.430 188.900 82.690 189.220 ;
        RECT 82.890 188.900 83.150 189.220 ;
        RECT 82.950 184.460 83.090 188.900 ;
        RECT 82.890 184.140 83.150 184.460 ;
        RECT 83.410 183.440 83.550 193.125 ;
        RECT 83.870 192.280 84.010 193.320 ;
        RECT 83.810 191.960 84.070 192.280 ;
        RECT 83.810 188.220 84.070 188.540 ;
        RECT 83.870 187.180 84.010 188.220 ;
        RECT 83.810 186.860 84.070 187.180 ;
        RECT 83.810 185.840 84.070 186.160 ;
        RECT 83.870 183.440 84.010 185.840 ;
        RECT 82.890 183.120 83.150 183.440 ;
        RECT 83.350 183.120 83.610 183.440 ;
        RECT 83.810 183.120 84.070 183.440 ;
        RECT 82.430 182.780 82.690 183.100 ;
        RECT 81.970 182.440 82.230 182.760 ;
        RECT 82.490 180.575 82.630 182.780 ;
        RECT 82.420 180.205 82.700 180.575 ;
        RECT 79.720 179.185 81.260 179.555 ;
        RECT 82.950 178.340 83.090 183.120 ;
        RECT 83.410 181.740 83.550 183.120 ;
        RECT 83.350 181.420 83.610 181.740 ;
        RECT 84.330 179.950 84.470 194.000 ;
        RECT 84.720 193.805 85.000 194.175 ;
        RECT 84.790 193.640 84.930 193.805 ;
        RECT 84.730 193.320 84.990 193.640 ;
        RECT 84.730 189.240 84.990 189.560 ;
        RECT 84.790 188.055 84.930 189.240 ;
        RECT 84.720 187.685 85.000 188.055 ;
        RECT 85.250 186.840 85.390 195.280 ;
        RECT 85.710 193.640 85.850 196.720 ;
        RECT 86.170 196.360 86.310 197.205 ;
        RECT 86.110 196.040 86.370 196.360 ;
        RECT 86.110 194.340 86.370 194.660 ;
        RECT 85.650 193.320 85.910 193.640 ;
        RECT 85.640 189.725 85.920 190.095 ;
        RECT 85.190 186.520 85.450 186.840 ;
        RECT 84.720 185.645 85.000 186.015 ;
        RECT 84.790 180.720 84.930 185.645 ;
        RECT 85.190 183.800 85.450 184.120 ;
        RECT 85.250 182.670 85.390 183.800 ;
        RECT 85.710 183.440 85.850 189.725 ;
        RECT 86.170 186.160 86.310 194.340 ;
        RECT 86.630 192.620 86.770 199.780 ;
        RECT 87.090 197.380 87.230 209.640 ;
        RECT 87.550 208.600 87.690 209.980 ;
        RECT 87.490 208.280 87.750 208.600 ;
        RECT 87.490 207.600 87.750 207.920 ;
        RECT 87.550 203.500 87.690 207.600 ;
        RECT 87.490 203.180 87.750 203.500 ;
        RECT 87.550 200.100 87.690 203.180 ;
        RECT 88.010 201.800 88.150 213.040 ;
        RECT 89.330 212.700 89.590 213.020 ;
        RECT 89.390 212.535 89.530 212.700 ;
        RECT 89.320 212.165 89.600 212.535 ;
        RECT 88.410 211.340 88.670 211.660 ;
        RECT 88.470 207.920 88.610 211.340 ;
        RECT 89.390 210.640 89.530 212.165 ;
        RECT 89.790 210.660 90.050 210.980 ;
        RECT 89.330 210.550 89.590 210.640 ;
        RECT 88.930 210.410 89.590 210.550 ;
        RECT 88.930 209.815 89.070 210.410 ;
        RECT 89.330 210.320 89.590 210.410 ;
        RECT 88.860 209.445 89.140 209.815 ;
        RECT 89.330 209.640 89.590 209.960 ;
        RECT 88.410 207.600 88.670 207.920 ;
        RECT 88.870 207.260 89.130 207.580 ;
        RECT 88.410 206.920 88.670 207.240 ;
        RECT 88.470 206.220 88.610 206.920 ;
        RECT 88.930 206.220 89.070 207.260 ;
        RECT 89.390 207.240 89.530 209.640 ;
        RECT 89.330 206.920 89.590 207.240 ;
        RECT 88.410 205.900 88.670 206.220 ;
        RECT 88.870 205.900 89.130 206.220 ;
        RECT 88.410 204.540 88.670 204.860 ;
        RECT 88.470 202.140 88.610 204.540 ;
        RECT 88.870 204.430 89.130 204.520 ;
        RECT 89.390 204.430 89.530 206.920 ;
        RECT 89.850 205.540 89.990 210.660 ;
        RECT 89.790 205.220 90.050 205.540 ;
        RECT 88.870 204.290 89.530 204.430 ;
        RECT 88.870 204.200 89.130 204.290 ;
        RECT 88.410 201.820 88.670 202.140 ;
        RECT 87.950 201.480 88.210 201.800 ;
        RECT 87.490 199.780 87.750 200.100 ;
        RECT 87.490 199.100 87.750 199.420 ;
        RECT 87.030 197.060 87.290 197.380 ;
        RECT 87.030 196.380 87.290 196.700 ;
        RECT 87.090 194.060 87.230 196.380 ;
        RECT 87.550 195.535 87.690 199.100 ;
        RECT 88.470 198.820 88.610 201.820 ;
        RECT 88.930 200.780 89.070 204.200 ;
        RECT 89.330 202.335 89.590 202.480 ;
        RECT 89.320 201.965 89.600 202.335 ;
        RECT 88.870 200.460 89.130 200.780 ;
        RECT 88.860 199.925 89.140 200.295 ;
        RECT 89.390 200.100 89.530 201.965 ;
        RECT 88.930 199.330 89.070 199.925 ;
        RECT 89.330 199.780 89.590 200.100 ;
        RECT 88.930 199.190 89.530 199.330 ;
        RECT 88.470 198.680 89.070 198.820 ;
        RECT 88.410 197.970 88.670 198.060 ;
        RECT 88.010 197.830 88.670 197.970 ;
        RECT 87.480 195.165 87.760 195.535 ;
        RECT 87.550 194.660 87.690 195.165 ;
        RECT 87.490 194.340 87.750 194.660 ;
        RECT 87.090 193.920 87.690 194.060 ;
        RECT 87.030 193.320 87.290 193.640 ;
        RECT 86.570 192.300 86.830 192.620 ;
        RECT 87.090 192.280 87.230 193.320 ;
        RECT 87.030 191.960 87.290 192.280 ;
        RECT 87.550 192.020 87.690 193.920 ;
        RECT 88.010 193.890 88.150 197.830 ;
        RECT 88.410 197.740 88.670 197.830 ;
        RECT 88.010 193.750 88.610 193.890 ;
        RECT 87.550 191.880 88.150 192.020 ;
        RECT 86.570 191.280 86.830 191.600 ;
        RECT 87.030 191.280 87.290 191.600 ;
        RECT 87.490 191.280 87.750 191.600 ;
        RECT 86.110 185.840 86.370 186.160 ;
        RECT 86.630 185.480 86.770 191.280 ;
        RECT 87.090 190.775 87.230 191.280 ;
        RECT 87.020 190.405 87.300 190.775 ;
        RECT 87.020 189.725 87.300 190.095 ;
        RECT 87.550 189.900 87.690 191.280 ;
        RECT 88.010 190.920 88.150 191.880 ;
        RECT 87.950 190.600 88.210 190.920 ;
        RECT 88.010 189.900 88.150 190.600 ;
        RECT 87.090 189.560 87.230 189.725 ;
        RECT 87.490 189.580 87.750 189.900 ;
        RECT 87.950 189.580 88.210 189.900 ;
        RECT 87.030 189.240 87.290 189.560 ;
        RECT 87.950 187.880 88.210 188.200 ;
        RECT 88.010 187.180 88.150 187.880 ;
        RECT 87.950 186.860 88.210 187.180 ;
        RECT 87.030 185.500 87.290 185.820 ;
        RECT 86.110 185.160 86.370 185.480 ;
        RECT 86.570 185.160 86.830 185.480 ;
        RECT 86.170 184.460 86.310 185.160 ;
        RECT 87.090 184.460 87.230 185.500 ;
        RECT 86.110 184.140 86.370 184.460 ;
        RECT 87.030 184.140 87.290 184.460 ;
        RECT 86.170 183.975 86.310 184.140 ;
        RECT 86.100 183.605 86.380 183.975 ;
        RECT 85.650 183.350 85.910 183.440 ;
        RECT 86.570 183.350 86.830 183.440 ;
        RECT 85.650 183.210 86.830 183.350 ;
        RECT 85.650 183.120 85.910 183.210 ;
        RECT 86.570 183.120 86.830 183.210 ;
        RECT 85.650 182.670 85.910 182.760 ;
        RECT 85.250 182.530 85.910 182.670 ;
        RECT 84.730 180.400 84.990 180.720 ;
        RECT 84.330 179.810 84.930 179.950 ;
        RECT 84.270 178.360 84.530 178.680 ;
        RECT 79.210 178.020 79.470 178.340 ;
        RECT 82.890 178.020 83.150 178.340 ;
        RECT 81.050 177.740 81.310 178.000 ;
        RECT 81.050 177.680 83.090 177.740 ;
        RECT 83.810 177.680 84.070 178.000 ;
        RECT 78.750 177.340 79.010 177.660 ;
        RECT 81.110 177.600 83.090 177.680 ;
        RECT 78.810 175.960 78.950 177.340 ;
        RECT 81.970 175.980 82.230 176.300 ;
        RECT 78.750 175.640 79.010 175.960 ;
        RECT 79.210 174.280 79.470 174.600 ;
        RECT 82.030 174.340 82.170 175.980 ;
        RECT 82.420 174.340 82.700 174.455 ;
        RECT 78.740 173.405 79.020 173.775 ;
        RECT 79.270 173.490 79.410 174.280 ;
        RECT 81.570 174.200 82.700 174.340 ;
        RECT 79.720 173.745 81.260 174.115 ;
        RECT 81.050 173.490 81.310 173.580 ;
        RECT 78.810 173.240 78.950 173.405 ;
        RECT 79.270 173.350 81.310 173.490 ;
        RECT 78.750 172.920 79.010 173.240 ;
        RECT 78.740 172.045 79.020 172.415 ;
        RECT 78.810 171.880 78.950 172.045 ;
        RECT 78.750 171.560 79.010 171.880 ;
        RECT 79.270 169.160 79.410 173.350 ;
        RECT 81.050 173.260 81.310 173.350 ;
        RECT 79.670 172.580 79.930 172.900 ;
        RECT 81.050 172.580 81.310 172.900 ;
        RECT 79.730 169.160 79.870 172.580 ;
        RECT 80.590 171.900 80.850 172.220 ;
        RECT 80.650 169.840 80.790 171.900 ;
        RECT 81.110 170.520 81.250 172.580 ;
        RECT 81.050 170.200 81.310 170.520 ;
        RECT 80.590 169.520 80.850 169.840 ;
        RECT 78.740 168.645 79.020 169.015 ;
        RECT 79.210 168.840 79.470 169.160 ;
        RECT 79.670 168.840 79.930 169.160 ;
        RECT 77.360 167.540 77.640 167.655 ;
        RECT 77.360 167.460 78.030 167.540 ;
        RECT 77.360 167.400 78.090 167.460 ;
        RECT 77.360 167.285 77.640 167.400 ;
        RECT 77.830 167.140 78.090 167.400 ;
        RECT 78.280 167.285 78.560 167.655 ;
        RECT 76.900 165.245 77.180 165.615 ;
        RECT 78.350 164.060 78.490 167.285 ;
        RECT 78.810 164.820 78.950 168.645 ;
        RECT 79.270 166.440 79.410 168.840 ;
        RECT 79.720 168.305 81.260 168.675 ;
        RECT 80.590 166.460 80.850 166.780 ;
        RECT 79.210 166.120 79.470 166.440 ;
        RECT 80.650 164.935 80.790 166.460 ;
        RECT 78.810 164.680 79.410 164.820 ;
        RECT 78.290 163.740 78.550 164.060 ;
        RECT 78.750 163.740 79.010 164.060 ;
        RECT 75.990 162.380 76.250 162.700 ;
        RECT 77.830 161.700 78.090 162.020 ;
        RECT 73.690 161.535 73.950 161.680 ;
        RECT 73.680 161.165 73.960 161.535 ;
        RECT 77.890 161.000 78.030 161.700 ;
        RECT 77.830 160.680 78.090 161.000 ;
        RECT 72.760 159.125 73.040 159.495 ;
        RECT 77.830 159.320 78.090 159.640 ;
        RECT 70.920 157.765 71.200 158.135 ;
        RECT 70.470 156.600 70.730 156.920 ;
        RECT 69.550 155.920 69.810 156.240 ;
        RECT 69.610 152.840 69.750 155.920 ;
        RECT 70.990 153.180 71.130 157.765 ;
        RECT 71.850 153.200 72.110 153.520 ;
        RECT 70.930 152.860 71.190 153.180 ;
        RECT 69.550 152.520 69.810 152.840 ;
        RECT 70.010 152.520 70.270 152.840 ;
        RECT 70.070 150.540 70.210 152.520 ;
        RECT 71.910 151.820 72.050 153.200 ;
        RECT 71.850 151.500 72.110 151.820 ;
        RECT 69.610 150.400 70.210 150.540 ;
        RECT 69.090 148.100 69.350 148.420 ;
        RECT 67.700 142.920 68.830 143.060 ;
        RECT 67.700 142.805 67.980 142.920 ;
        RECT 67.710 142.320 67.970 142.640 ;
        RECT 67.240 140.765 67.520 141.135 ;
        RECT 67.310 139.920 67.450 140.765 ;
        RECT 67.250 139.600 67.510 139.920 ;
        RECT 66.790 137.735 67.050 137.880 ;
        RECT 66.780 137.365 67.060 137.735 ;
        RECT 64.950 133.820 65.210 134.140 ;
        RECT 65.410 133.820 65.670 134.140 ;
        RECT 65.870 133.820 66.130 134.140 ;
        RECT 65.010 132.100 65.150 133.820 ;
        RECT 67.770 132.100 67.910 142.320 ;
        RECT 68.170 141.640 68.430 141.960 ;
        RECT 69.610 141.700 69.750 150.400 ;
        RECT 70.010 149.800 70.270 150.120 ;
        RECT 70.070 142.640 70.210 149.800 ;
        RECT 72.310 148.100 72.570 148.420 ;
        RECT 70.470 147.420 70.730 147.740 ;
        RECT 70.530 143.660 70.670 147.420 ;
        RECT 70.930 145.720 71.190 146.040 ;
        RECT 70.990 144.680 71.130 145.720 ;
        RECT 70.930 144.360 71.190 144.680 ;
        RECT 71.390 144.535 71.650 144.680 ;
        RECT 71.380 144.165 71.660 144.535 ;
        RECT 70.470 143.340 70.730 143.660 ;
        RECT 71.850 143.340 72.110 143.660 ;
        RECT 70.930 142.660 71.190 142.980 ;
        RECT 70.010 142.320 70.270 142.640 ;
        RECT 68.230 140.940 68.370 141.640 ;
        RECT 69.150 141.560 69.750 141.700 ;
        RECT 68.170 140.620 68.430 140.940 ;
        RECT 64.950 131.780 65.210 132.100 ;
        RECT 67.710 131.780 67.970 132.100 ;
        RECT 67.770 131.080 67.910 131.780 ;
        RECT 69.150 131.420 69.290 141.560 ;
        RECT 70.990 137.880 71.130 142.660 ;
        RECT 71.390 142.320 71.650 142.640 ;
        RECT 71.450 139.240 71.590 142.320 ;
        RECT 71.910 140.260 72.050 143.340 ;
        RECT 72.370 141.815 72.510 148.100 ;
        RECT 72.830 145.360 72.970 159.125 ;
        RECT 76.910 158.980 77.170 159.300 ;
        RECT 76.970 158.280 77.110 158.980 ;
        RECT 77.370 158.640 77.630 158.960 ;
        RECT 76.910 157.960 77.170 158.280 ;
        RECT 76.970 157.455 77.110 157.960 ;
        RECT 76.900 157.085 77.180 157.455 ;
        RECT 76.910 155.920 77.170 156.240 ;
        RECT 75.530 154.220 75.790 154.540 ;
        RECT 75.590 153.940 75.730 154.220 ;
        RECT 74.210 153.800 75.730 153.940 ;
        RECT 75.990 153.880 76.250 154.200 ;
        RECT 74.210 153.520 74.350 153.800 ;
        RECT 74.150 153.200 74.410 153.520 ;
        RECT 76.050 153.260 76.190 153.880 ;
        RECT 76.450 153.540 76.710 153.860 ;
        RECT 75.590 153.120 76.190 153.260 ;
        RECT 75.590 147.400 75.730 153.120 ;
        RECT 75.990 152.520 76.250 152.840 ;
        RECT 76.050 148.080 76.190 152.520 ;
        RECT 76.510 150.800 76.650 153.540 ;
        RECT 76.450 150.480 76.710 150.800 ;
        RECT 75.990 147.760 76.250 148.080 ;
        RECT 75.530 147.080 75.790 147.400 ;
        RECT 75.530 145.720 75.790 146.040 ;
        RECT 72.770 145.040 73.030 145.360 ;
        RECT 74.610 145.270 74.870 145.360 ;
        RECT 73.680 144.845 73.960 145.215 ;
        RECT 74.210 145.130 74.870 145.270 ;
        RECT 73.750 143.660 73.890 144.845 ;
        RECT 73.690 143.340 73.950 143.660 ;
        RECT 72.770 142.660 73.030 142.980 ;
        RECT 72.300 141.445 72.580 141.815 ;
        RECT 71.850 139.940 72.110 140.260 ;
        RECT 72.310 139.940 72.570 140.260 ;
        RECT 71.390 138.920 71.650 139.240 ;
        RECT 70.930 137.560 71.190 137.880 ;
        RECT 70.470 136.880 70.730 137.200 ;
        RECT 70.010 136.200 70.270 136.520 ;
        RECT 69.550 135.015 69.810 135.160 ;
        RECT 69.540 134.645 69.820 135.015 ;
        RECT 69.090 131.100 69.350 131.420 ;
        RECT 67.710 130.760 67.970 131.080 ;
        RECT 69.150 129.720 69.290 131.100 ;
        RECT 63.110 129.400 63.370 129.720 ;
        RECT 69.090 129.400 69.350 129.720 ;
        RECT 60.285 127.505 61.825 127.875 ;
        RECT 69.610 126.660 69.750 134.645 ;
        RECT 70.070 134.480 70.210 136.200 ;
        RECT 70.530 135.500 70.670 136.880 ;
        RECT 70.990 136.375 71.130 137.560 ;
        RECT 71.390 136.880 71.650 137.200 ;
        RECT 70.920 136.005 71.200 136.375 ;
        RECT 70.470 135.180 70.730 135.500 ;
        RECT 70.010 134.160 70.270 134.480 ;
        RECT 70.070 132.440 70.210 134.160 ;
        RECT 71.450 132.780 71.590 136.880 ;
        RECT 72.370 134.820 72.510 139.940 ;
        RECT 72.830 139.240 72.970 142.660 ;
        RECT 73.690 139.940 73.950 140.260 ;
        RECT 72.770 138.920 73.030 139.240 ;
        RECT 73.230 137.560 73.490 137.880 ;
        RECT 73.290 134.820 73.430 137.560 ;
        RECT 73.750 135.500 73.890 139.940 ;
        RECT 73.690 135.180 73.950 135.500 ;
        RECT 72.310 134.500 72.570 134.820 ;
        RECT 73.230 134.500 73.490 134.820 ;
        RECT 71.390 132.460 71.650 132.780 ;
        RECT 70.010 132.120 70.270 132.440 ;
        RECT 70.070 129.720 70.210 132.120 ;
        RECT 72.310 130.760 72.570 131.080 ;
        RECT 70.010 129.400 70.270 129.720 ;
        RECT 69.550 126.340 69.810 126.660 ;
        RECT 70.070 126.320 70.210 129.400 ;
        RECT 72.370 129.380 72.510 130.760 ;
        RECT 74.210 130.060 74.350 145.130 ;
        RECT 74.610 145.040 74.870 145.130 ;
        RECT 75.070 144.700 75.330 145.020 ;
        RECT 75.130 142.980 75.270 144.700 ;
        RECT 75.070 142.660 75.330 142.980 ;
        RECT 75.590 142.640 75.730 145.720 ;
        RECT 76.050 144.680 76.190 147.760 ;
        RECT 75.990 144.360 76.250 144.680 ;
        RECT 75.530 142.320 75.790 142.640 ;
        RECT 76.970 142.300 77.110 155.920 ;
        RECT 77.430 153.180 77.570 158.640 ;
        RECT 77.890 156.920 78.030 159.320 ;
        RECT 77.830 156.600 78.090 156.920 ;
        RECT 77.370 152.860 77.630 153.180 ;
        RECT 77.830 152.520 78.090 152.840 ;
        RECT 77.890 151.820 78.030 152.520 ;
        RECT 77.830 151.500 78.090 151.820 ;
        RECT 77.890 148.760 78.030 151.500 ;
        RECT 78.350 151.480 78.490 163.740 ;
        RECT 78.810 162.360 78.950 163.740 ;
        RECT 78.750 162.040 79.010 162.360 ;
        RECT 79.270 159.890 79.410 164.680 ;
        RECT 80.580 164.565 80.860 164.935 ;
        RECT 79.720 162.865 81.260 163.235 ;
        RECT 81.570 162.360 81.710 174.200 ;
        RECT 82.420 174.085 82.700 174.200 ;
        RECT 81.970 172.580 82.230 172.900 ;
        RECT 82.030 172.220 82.170 172.580 ;
        RECT 81.970 171.900 82.230 172.220 ;
        RECT 82.430 168.840 82.690 169.160 ;
        RECT 81.960 167.965 82.240 168.335 ;
        RECT 82.030 167.460 82.170 167.965 ;
        RECT 81.970 167.140 82.230 167.460 ;
        RECT 81.970 163.400 82.230 163.720 ;
        RECT 82.030 162.360 82.170 163.400 ;
        RECT 81.510 162.040 81.770 162.360 ;
        RECT 81.970 162.040 82.230 162.360 ;
        RECT 81.970 161.360 82.230 161.680 ;
        RECT 78.810 159.750 79.410 159.890 ;
        RECT 78.810 155.300 78.950 159.750 ;
        RECT 82.030 159.640 82.170 161.360 ;
        RECT 79.200 159.125 79.480 159.495 ;
        RECT 81.970 159.320 82.230 159.640 ;
        RECT 79.210 158.980 79.470 159.125 ;
        RECT 81.510 158.300 81.770 158.620 ;
        RECT 81.970 158.300 82.230 158.620 ;
        RECT 79.720 157.425 81.260 157.795 ;
        RECT 81.570 156.580 81.710 158.300 ;
        RECT 82.030 157.260 82.170 158.300 ;
        RECT 81.970 156.940 82.230 157.260 ;
        RECT 81.510 156.260 81.770 156.580 ;
        RECT 78.810 155.160 79.410 155.300 ;
        RECT 78.750 154.220 79.010 154.540 ;
        RECT 78.290 151.160 78.550 151.480 ;
        RECT 77.830 148.440 78.090 148.760 ;
        RECT 78.810 143.660 78.950 154.220 ;
        RECT 79.270 151.220 79.410 155.160 ;
        RECT 79.720 151.985 81.260 152.355 ;
        RECT 79.270 151.080 79.870 151.220 ;
        RECT 79.730 148.420 79.870 151.080 ;
        RECT 81.570 148.420 81.710 156.260 ;
        RECT 81.970 155.240 82.230 155.560 ;
        RECT 82.030 154.735 82.170 155.240 ;
        RECT 81.960 154.365 82.240 154.735 ;
        RECT 82.490 154.540 82.630 168.840 ;
        RECT 82.950 167.800 83.090 177.600 ;
        RECT 83.350 177.340 83.610 177.660 ;
        RECT 83.410 175.700 83.550 177.340 ;
        RECT 83.870 176.300 84.010 177.680 ;
        RECT 84.330 176.495 84.470 178.360 ;
        RECT 84.790 177.855 84.930 179.810 ;
        RECT 85.250 178.680 85.390 182.530 ;
        RECT 85.650 182.440 85.910 182.530 ;
        RECT 85.650 180.740 85.910 181.060 ;
        RECT 85.190 178.360 85.450 178.680 ;
        RECT 84.720 177.485 85.000 177.855 ;
        RECT 83.810 175.980 84.070 176.300 ;
        RECT 84.260 176.125 84.540 176.495 ;
        RECT 83.410 175.560 84.010 175.700 ;
        RECT 83.870 174.600 84.010 175.560 ;
        RECT 83.810 174.280 84.070 174.600 ;
        RECT 83.870 173.580 84.010 174.280 ;
        RECT 83.810 173.260 84.070 173.580 ;
        RECT 84.730 173.260 84.990 173.580 ;
        RECT 84.270 172.810 84.530 172.900 ;
        RECT 84.790 172.810 84.930 173.260 ;
        RECT 85.250 173.240 85.390 178.360 ;
        RECT 85.190 172.920 85.450 173.240 ;
        RECT 84.270 172.670 84.930 172.810 ;
        RECT 84.270 172.580 84.530 172.670 ;
        RECT 84.270 171.900 84.530 172.220 ;
        RECT 83.340 171.365 83.620 171.735 ;
        RECT 83.410 170.180 83.550 171.365 ;
        RECT 84.330 170.180 84.470 171.900 ;
        RECT 83.350 169.860 83.610 170.180 ;
        RECT 84.270 169.860 84.530 170.180 ;
        RECT 82.890 167.480 83.150 167.800 ;
        RECT 82.890 167.030 83.150 167.120 ;
        RECT 83.410 167.030 83.550 169.860 ;
        RECT 83.810 169.520 84.070 169.840 ;
        RECT 82.890 166.975 83.550 167.030 ;
        RECT 82.890 166.890 83.620 166.975 ;
        RECT 82.890 166.800 83.150 166.890 ;
        RECT 83.340 166.605 83.620 166.890 ;
        RECT 82.890 163.400 83.150 163.720 ;
        RECT 82.950 158.960 83.090 163.400 ;
        RECT 83.870 159.640 84.010 169.520 ;
        RECT 84.270 169.180 84.530 169.500 ;
        RECT 84.330 162.700 84.470 169.180 ;
        RECT 84.790 169.160 84.930 172.670 ;
        RECT 85.710 170.375 85.850 180.740 ;
        RECT 87.090 178.340 87.230 184.140 ;
        RECT 87.950 181.420 88.210 181.740 ;
        RECT 87.030 178.020 87.290 178.340 ;
        RECT 87.090 177.175 87.230 178.020 ;
        RECT 88.010 178.000 88.150 181.420 ;
        RECT 88.470 180.720 88.610 193.750 ;
        RECT 88.930 191.600 89.070 198.680 ;
        RECT 89.390 198.060 89.530 199.190 ;
        RECT 89.330 197.740 89.590 198.060 ;
        RECT 89.850 197.040 89.990 205.220 ;
        RECT 90.310 197.460 90.450 214.150 ;
        RECT 91.170 214.060 91.430 214.380 ;
        RECT 91.690 212.680 91.830 216.100 ;
        RECT 94.390 215.990 94.650 216.080 ;
        RECT 94.910 215.990 95.050 216.870 ;
        RECT 95.310 216.780 95.570 216.870 ;
        RECT 96.230 216.780 96.490 217.100 ;
        RECT 96.290 216.615 96.430 216.780 ;
        RECT 96.220 216.245 96.500 216.615 ;
        RECT 97.150 216.440 97.410 216.760 ;
        RECT 94.390 215.850 95.050 215.990 ;
        RECT 94.390 215.760 94.650 215.850 ;
        RECT 95.310 215.760 95.570 216.080 ;
        RECT 92.080 214.885 92.360 215.255 ;
        RECT 93.930 215.080 94.190 215.400 ;
        RECT 92.150 214.040 92.290 214.885 ;
        RECT 92.090 213.720 92.350 214.040 ;
        RECT 93.010 213.720 93.270 214.040 ;
        RECT 92.550 213.380 92.810 213.700 ;
        RECT 91.630 212.360 91.890 212.680 ;
        RECT 92.610 211.660 92.750 213.380 ;
        RECT 92.550 211.340 92.810 211.660 ;
        RECT 92.090 211.000 92.350 211.320 ;
        RECT 93.070 211.060 93.210 213.720 ;
        RECT 90.710 210.320 90.970 210.640 ;
        RECT 90.770 205.880 90.910 210.320 ;
        RECT 92.150 208.260 92.290 211.000 ;
        RECT 92.610 210.920 93.210 211.060 ;
        RECT 92.610 209.960 92.750 210.920 ;
        RECT 93.460 210.805 93.740 211.175 ;
        RECT 92.550 209.640 92.810 209.960 ;
        RECT 93.000 209.445 93.280 209.815 ;
        RECT 93.070 208.600 93.210 209.445 ;
        RECT 93.010 208.280 93.270 208.600 ;
        RECT 92.090 207.940 92.350 208.260 ;
        RECT 93.010 207.260 93.270 207.580 ;
        RECT 91.630 205.900 91.890 206.220 ;
        RECT 92.090 205.900 92.350 206.220 ;
        RECT 90.710 205.560 90.970 205.880 ;
        RECT 90.770 198.255 90.910 205.560 ;
        RECT 91.170 199.100 91.430 199.420 ;
        RECT 90.700 197.885 90.980 198.255 ;
        RECT 90.310 197.320 90.910 197.460 ;
        RECT 89.790 196.720 90.050 197.040 ;
        RECT 90.250 196.720 90.510 197.040 ;
        RECT 89.790 196.040 90.050 196.360 ;
        RECT 89.330 194.680 89.590 195.000 ;
        RECT 89.390 193.495 89.530 194.680 ;
        RECT 89.850 193.640 89.990 196.040 ;
        RECT 90.310 193.980 90.450 196.720 ;
        RECT 90.250 193.660 90.510 193.980 ;
        RECT 89.320 193.125 89.600 193.495 ;
        RECT 89.790 193.320 90.050 193.640 ;
        RECT 90.770 192.280 90.910 197.320 ;
        RECT 89.790 192.190 90.050 192.280 ;
        RECT 89.390 192.050 90.050 192.190 ;
        RECT 89.390 192.020 89.530 192.050 ;
        RECT 89.310 191.880 89.530 192.020 ;
        RECT 89.790 191.960 90.050 192.050 ;
        RECT 90.710 191.960 90.970 192.280 ;
        RECT 88.870 191.280 89.130 191.600 ;
        RECT 89.310 191.170 89.450 191.880 ;
        RECT 89.790 191.280 90.050 191.600 ;
        RECT 89.310 191.030 89.530 191.170 ;
        RECT 88.860 189.725 89.140 190.095 ;
        RECT 88.930 188.540 89.070 189.725 ;
        RECT 88.870 188.220 89.130 188.540 ;
        RECT 89.390 188.200 89.530 191.030 ;
        RECT 89.330 187.880 89.590 188.200 ;
        RECT 89.850 187.340 89.990 191.280 ;
        RECT 90.250 188.560 90.510 188.880 ;
        RECT 88.930 187.200 89.990 187.340 ;
        RECT 88.930 182.615 89.070 187.200 ;
        RECT 89.330 186.520 89.590 186.840 ;
        RECT 88.860 182.245 89.140 182.615 ;
        RECT 88.860 181.565 89.140 181.935 ;
        RECT 88.870 181.420 89.130 181.565 ;
        RECT 89.390 181.400 89.530 186.520 ;
        RECT 90.310 185.480 90.450 188.560 ;
        RECT 90.250 185.160 90.510 185.480 ;
        RECT 90.310 184.460 90.450 185.160 ;
        RECT 90.250 184.140 90.510 184.460 ;
        RECT 90.250 183.460 90.510 183.780 ;
        RECT 89.790 182.780 90.050 183.100 ;
        RECT 89.330 181.080 89.590 181.400 ;
        RECT 88.410 180.400 88.670 180.720 ;
        RECT 88.860 179.780 89.140 179.895 ;
        RECT 88.860 179.640 89.530 179.780 ;
        RECT 88.860 179.525 89.140 179.640 ;
        RECT 87.950 177.680 88.210 178.000 ;
        RECT 89.390 177.320 89.530 179.640 ;
        RECT 89.850 178.340 89.990 182.780 ;
        RECT 90.310 178.680 90.450 183.460 ;
        RECT 91.230 183.440 91.370 199.100 ;
        RECT 91.690 198.060 91.830 205.900 ;
        RECT 92.150 205.200 92.290 205.900 ;
        RECT 92.540 205.365 92.820 205.735 ;
        RECT 92.090 204.880 92.350 205.200 ;
        RECT 91.630 197.740 91.890 198.060 ;
        RECT 92.150 197.460 92.290 204.880 ;
        RECT 92.610 201.800 92.750 205.365 ;
        RECT 92.550 201.480 92.810 201.800 ;
        RECT 92.550 200.460 92.810 200.780 ;
        RECT 92.610 199.615 92.750 200.460 ;
        RECT 92.540 199.245 92.820 199.615 ;
        RECT 91.690 197.320 92.290 197.460 ;
        RECT 91.690 191.260 91.830 197.320 ;
        RECT 92.080 195.845 92.360 196.215 ;
        RECT 92.550 196.040 92.810 196.360 ;
        RECT 92.150 195.340 92.290 195.845 ;
        RECT 92.090 195.020 92.350 195.340 ;
        RECT 91.630 190.940 91.890 191.260 ;
        RECT 91.630 189.580 91.890 189.900 ;
        RECT 91.690 188.200 91.830 189.580 ;
        RECT 91.630 187.880 91.890 188.200 ;
        RECT 92.150 187.180 92.290 195.020 ;
        RECT 92.610 189.900 92.750 196.040 ;
        RECT 93.070 194.320 93.210 207.260 ;
        RECT 93.530 202.480 93.670 210.805 ;
        RECT 93.470 202.160 93.730 202.480 ;
        RECT 93.530 200.780 93.670 202.160 ;
        RECT 93.470 200.460 93.730 200.780 ;
        RECT 93.990 196.700 94.130 215.080 ;
        RECT 94.390 211.340 94.650 211.660 ;
        RECT 94.450 210.980 94.590 211.340 ;
        RECT 94.390 210.660 94.650 210.980 ;
        RECT 94.450 209.815 94.590 210.660 ;
        RECT 94.380 209.445 94.660 209.815 ;
        RECT 95.370 208.940 95.510 215.760 ;
        RECT 96.690 215.420 96.950 215.740 ;
        RECT 95.770 213.380 96.030 213.700 ;
        RECT 95.830 211.320 95.970 213.380 ;
        RECT 96.750 212.680 96.890 215.420 ;
        RECT 96.690 212.360 96.950 212.680 ;
        RECT 96.220 211.485 96.500 211.855 ;
        RECT 95.770 211.000 96.030 211.320 ;
        RECT 96.290 210.550 96.430 211.485 ;
        RECT 96.750 210.980 96.890 212.360 ;
        RECT 97.210 210.980 97.350 216.440 ;
        RECT 97.670 215.255 97.810 218.480 ;
        RECT 98.070 217.800 98.330 218.120 ;
        RECT 97.600 214.885 97.880 215.255 ;
        RECT 96.690 210.660 96.950 210.980 ;
        RECT 97.150 210.660 97.410 210.980 ;
        RECT 97.610 210.660 97.870 210.980 ;
        RECT 95.830 210.410 96.430 210.550 ;
        RECT 94.390 208.620 94.650 208.940 ;
        RECT 95.310 208.620 95.570 208.940 ;
        RECT 94.450 200.100 94.590 208.620 ;
        RECT 95.370 207.920 95.510 208.620 ;
        RECT 94.850 207.600 95.110 207.920 ;
        RECT 95.310 207.600 95.570 207.920 ;
        RECT 94.910 205.450 95.050 207.600 ;
        RECT 95.830 205.540 95.970 210.410 ;
        RECT 96.750 209.020 96.890 210.660 ;
        RECT 96.290 208.880 96.890 209.020 ;
        RECT 95.310 205.450 95.570 205.540 ;
        RECT 94.910 205.310 95.570 205.450 ;
        RECT 95.310 205.220 95.570 205.310 ;
        RECT 95.770 205.220 96.030 205.540 ;
        RECT 95.370 202.900 95.510 205.220 ;
        RECT 95.760 202.900 96.040 203.015 ;
        RECT 94.850 202.500 95.110 202.820 ;
        RECT 95.370 202.760 96.040 202.900 ;
        RECT 95.760 202.645 96.040 202.760 ;
        RECT 94.910 201.655 95.050 202.500 ;
        RECT 95.310 202.160 95.570 202.480 ;
        RECT 94.840 201.285 95.120 201.655 ;
        RECT 94.840 200.605 95.120 200.975 ;
        RECT 94.910 200.440 95.050 200.605 ;
        RECT 94.850 200.120 95.110 200.440 ;
        RECT 94.390 199.780 94.650 200.100 ;
        RECT 93.470 196.380 93.730 196.700 ;
        RECT 93.930 196.380 94.190 196.700 ;
        RECT 93.010 194.000 93.270 194.320 ;
        RECT 93.010 193.320 93.270 193.640 ;
        RECT 93.070 191.600 93.210 193.320 ;
        RECT 93.530 192.280 93.670 196.380 ;
        RECT 93.470 191.960 93.730 192.280 ;
        RECT 93.010 191.280 93.270 191.600 ;
        RECT 92.550 189.580 92.810 189.900 ;
        RECT 92.610 188.790 92.750 189.580 ;
        RECT 93.010 188.790 93.270 188.880 ;
        RECT 92.610 188.650 93.270 188.790 ;
        RECT 93.010 188.560 93.270 188.650 ;
        RECT 93.530 187.340 93.670 191.960 ;
        RECT 93.990 188.790 94.130 196.380 ;
        RECT 94.450 196.215 94.590 199.780 ;
        RECT 94.380 195.845 94.660 196.215 ;
        RECT 94.910 192.620 95.050 200.120 ;
        RECT 95.370 197.040 95.510 202.160 ;
        RECT 95.770 201.480 96.030 201.800 ;
        RECT 95.830 200.100 95.970 201.480 ;
        RECT 96.290 200.860 96.430 208.880 ;
        RECT 97.150 208.280 97.410 208.600 ;
        RECT 97.210 207.240 97.350 208.280 ;
        RECT 97.150 206.920 97.410 207.240 ;
        RECT 97.670 206.220 97.810 210.660 ;
        RECT 98.130 208.600 98.270 217.800 ;
        RECT 101.350 216.420 101.490 219.160 ;
        RECT 101.290 216.100 101.550 216.420 ;
        RECT 99.155 214.545 100.695 214.915 ;
        RECT 101.350 214.040 101.490 216.100 ;
        RECT 98.990 213.720 99.250 214.040 ;
        RECT 101.290 213.720 101.550 214.040 ;
        RECT 98.530 213.040 98.790 213.360 ;
        RECT 98.590 211.175 98.730 213.040 ;
        RECT 98.520 210.805 98.800 211.175 ;
        RECT 99.050 210.300 99.190 213.720 ;
        RECT 101.290 213.040 101.550 213.360 ;
        RECT 101.350 212.680 101.490 213.040 ;
        RECT 99.910 212.590 100.170 212.680 ;
        RECT 99.910 212.450 100.570 212.590 ;
        RECT 99.910 212.360 100.170 212.450 ;
        RECT 100.430 210.980 100.570 212.450 ;
        RECT 101.290 212.360 101.550 212.680 ;
        RECT 100.370 210.660 100.630 210.980 ;
        RECT 98.990 209.980 99.250 210.300 ;
        RECT 99.155 209.105 100.695 209.475 ;
        RECT 98.070 208.280 98.330 208.600 ;
        RECT 97.610 205.900 97.870 206.220 ;
        RECT 96.690 205.220 96.950 205.540 ;
        RECT 97.140 205.365 97.420 205.735 ;
        RECT 97.150 205.220 97.410 205.365 ;
        RECT 96.750 204.940 96.890 205.220 ;
        RECT 96.750 204.800 97.810 204.940 ;
        RECT 96.690 204.430 96.950 204.520 ;
        RECT 96.690 204.290 97.350 204.430 ;
        RECT 96.690 204.200 96.950 204.290 ;
        RECT 96.680 203.325 96.960 203.695 ;
        RECT 96.750 202.140 96.890 203.325 ;
        RECT 96.690 201.820 96.950 202.140 ;
        RECT 97.210 201.655 97.350 204.290 ;
        RECT 97.670 203.500 97.810 204.800 ;
        RECT 98.130 203.500 98.270 208.280 ;
        RECT 102.270 207.920 102.410 219.500 ;
        RECT 102.670 218.480 102.930 218.800 ;
        RECT 102.730 217.100 102.870 218.480 ;
        RECT 103.130 217.800 103.390 218.120 ;
        RECT 102.670 216.780 102.930 217.100 ;
        RECT 102.670 212.360 102.930 212.680 ;
        RECT 98.530 207.260 98.790 207.580 ;
        RECT 100.430 207.520 101.490 207.660 ;
        RECT 101.750 207.600 102.010 207.920 ;
        RECT 102.210 207.600 102.470 207.920 ;
        RECT 97.610 203.180 97.870 203.500 ;
        RECT 98.070 203.180 98.330 203.500 ;
        RECT 98.590 202.900 98.730 207.260 ;
        RECT 100.430 207.240 100.570 207.520 ;
        RECT 98.990 206.920 99.250 207.240 ;
        RECT 100.370 206.920 100.630 207.240 ;
        RECT 100.830 206.920 101.090 207.240 ;
        RECT 99.050 206.130 99.190 206.920 ;
        RECT 99.050 205.990 100.570 206.130 ;
        RECT 99.050 205.540 99.190 205.990 ;
        RECT 98.990 205.220 99.250 205.540 ;
        RECT 99.910 205.220 100.170 205.540 ;
        RECT 99.970 204.520 100.110 205.220 ;
        RECT 99.910 204.200 100.170 204.520 ;
        RECT 100.430 204.430 100.570 205.990 ;
        RECT 100.890 205.450 101.030 206.920 ;
        RECT 101.350 206.415 101.490 207.520 ;
        RECT 101.810 207.240 101.950 207.600 ;
        RECT 101.750 206.920 102.010 207.240 ;
        RECT 101.280 206.045 101.560 206.415 ;
        RECT 102.730 206.300 102.870 212.360 ;
        RECT 103.190 207.920 103.330 217.800 ;
        RECT 103.650 216.420 103.790 219.500 ;
        RECT 107.270 219.160 107.530 219.480 ;
        RECT 107.330 218.800 107.470 219.160 ;
        RECT 107.270 218.480 107.530 218.800 ;
        RECT 104.970 218.140 105.230 218.460 ;
        RECT 103.590 216.100 103.850 216.420 ;
        RECT 103.580 215.565 103.860 215.935 ;
        RECT 103.650 214.380 103.790 215.565 ;
        RECT 103.590 214.060 103.850 214.380 ;
        RECT 103.650 213.360 103.790 214.060 ;
        RECT 103.590 213.040 103.850 213.360 ;
        RECT 104.510 212.700 104.770 213.020 ;
        RECT 103.590 210.660 103.850 210.980 ;
        RECT 103.650 208.260 103.790 210.660 ;
        RECT 104.570 210.640 104.710 212.700 ;
        RECT 104.510 210.320 104.770 210.640 ;
        RECT 104.050 209.640 104.310 209.960 ;
        RECT 104.510 209.640 104.770 209.960 ;
        RECT 103.590 207.940 103.850 208.260 ;
        RECT 104.110 207.920 104.250 209.640 ;
        RECT 104.570 208.940 104.710 209.640 ;
        RECT 104.510 208.620 104.770 208.940 ;
        RECT 105.030 207.920 105.170 218.140 ;
        RECT 107.270 216.670 107.530 216.760 ;
        RECT 107.270 216.530 108.390 216.670 ;
        RECT 107.270 216.440 107.530 216.530 ;
        RECT 106.350 215.080 106.610 215.400 ;
        RECT 106.410 213.360 106.550 215.080 ;
        RECT 107.720 214.885 108.000 215.255 ;
        RECT 107.790 213.360 107.930 214.885 ;
        RECT 106.350 213.040 106.610 213.360 ;
        RECT 107.730 213.040 107.990 213.360 ;
        RECT 106.800 212.420 107.080 212.535 ;
        RECT 107.270 212.420 107.530 212.680 ;
        RECT 106.800 212.360 107.530 212.420 ;
        RECT 106.800 212.280 107.470 212.360 ;
        RECT 106.800 212.165 107.080 212.280 ;
        RECT 105.420 211.740 105.700 211.855 ;
        RECT 105.420 211.600 106.550 211.740 ;
        RECT 105.420 211.485 105.700 211.600 ;
        RECT 105.890 210.660 106.150 210.980 ;
        RECT 103.130 207.600 103.390 207.920 ;
        RECT 104.050 207.600 104.310 207.920 ;
        RECT 104.970 207.600 105.230 207.920 ;
        RECT 103.590 207.260 103.850 207.580 ;
        RECT 103.650 206.980 103.790 207.260 ;
        RECT 104.040 206.980 104.320 207.095 ;
        RECT 103.650 206.840 104.320 206.980 ;
        RECT 104.040 206.725 104.320 206.840 ;
        RECT 103.120 206.300 103.400 206.415 ;
        RECT 102.730 206.160 103.400 206.300 ;
        RECT 105.030 206.220 105.170 207.600 ;
        RECT 103.120 206.045 103.400 206.160 ;
        RECT 104.510 205.900 104.770 206.220 ;
        RECT 104.970 205.900 105.230 206.220 ;
        RECT 100.890 205.310 102.410 205.450 ;
        RECT 101.290 204.430 101.550 204.520 ;
        RECT 100.430 204.290 101.030 204.430 ;
        RECT 99.155 203.665 100.695 204.035 ;
        RECT 100.890 203.410 101.030 204.290 ;
        RECT 101.290 204.290 101.950 204.430 ;
        RECT 101.290 204.200 101.550 204.290 ;
        RECT 97.670 202.760 98.730 202.900 ;
        RECT 100.430 203.270 101.030 203.410 ;
        RECT 101.280 203.325 101.560 203.695 ;
        RECT 97.140 201.285 97.420 201.655 ;
        RECT 97.140 200.860 97.420 200.975 ;
        RECT 96.290 200.720 97.420 200.860 ;
        RECT 97.140 200.605 97.420 200.720 ;
        RECT 97.210 200.440 97.350 200.605 ;
        RECT 97.150 200.120 97.410 200.440 ;
        RECT 95.770 200.010 96.030 200.100 ;
        RECT 95.770 199.870 96.430 200.010 ;
        RECT 95.770 199.780 96.030 199.870 ;
        RECT 95.770 198.760 96.030 199.080 ;
        RECT 95.310 196.720 95.570 197.040 ;
        RECT 95.830 193.980 95.970 198.760 ;
        RECT 96.290 198.060 96.430 199.870 ;
        RECT 96.680 199.245 96.960 199.615 ;
        RECT 97.150 199.440 97.410 199.760 ;
        RECT 96.690 199.100 96.950 199.245 ;
        RECT 96.230 197.740 96.490 198.060 ;
        RECT 96.230 196.380 96.490 196.700 ;
        RECT 95.770 193.660 96.030 193.980 ;
        RECT 94.850 192.300 95.110 192.620 ;
        RECT 94.850 191.280 95.110 191.600 ;
        RECT 95.310 191.280 95.570 191.600 ;
        RECT 94.390 190.600 94.650 190.920 ;
        RECT 94.450 189.560 94.590 190.600 ;
        RECT 94.910 189.900 95.050 191.280 ;
        RECT 94.850 189.580 95.110 189.900 ;
        RECT 94.390 189.240 94.650 189.560 ;
        RECT 95.370 189.300 95.510 191.280 ;
        RECT 94.910 189.160 95.510 189.300 ;
        RECT 94.910 188.880 95.050 189.160 ;
        RECT 93.990 188.650 94.590 188.790 ;
        RECT 94.450 188.110 94.590 188.650 ;
        RECT 94.850 188.560 95.110 188.880 ;
        RECT 93.070 187.200 93.670 187.340 ;
        RECT 93.990 187.970 94.590 188.110 ;
        RECT 92.090 186.860 92.350 187.180 ;
        RECT 93.070 183.780 93.210 187.200 ;
        RECT 93.460 186.325 93.740 186.695 ;
        RECT 93.010 183.460 93.270 183.780 ;
        RECT 91.170 183.120 91.430 183.440 ;
        RECT 92.090 183.295 92.350 183.440 ;
        RECT 92.080 182.925 92.360 183.295 ;
        RECT 91.160 180.885 91.440 181.255 ;
        RECT 93.530 181.060 93.670 186.325 ;
        RECT 93.990 183.440 94.130 187.970 ;
        RECT 94.840 187.685 95.120 188.055 ;
        RECT 94.910 187.340 95.050 187.685 ;
        RECT 94.450 187.200 95.050 187.340 ;
        RECT 93.930 183.120 94.190 183.440 ;
        RECT 91.230 180.720 91.370 180.885 ;
        RECT 93.470 180.740 93.730 181.060 ;
        RECT 91.170 180.400 91.430 180.720 ;
        RECT 90.250 178.360 90.510 178.680 ;
        RECT 89.790 178.020 90.050 178.340 ;
        RECT 89.790 177.340 90.050 177.660 ;
        RECT 87.020 176.805 87.300 177.175 ;
        RECT 89.330 177.000 89.590 177.320 ;
        RECT 89.850 177.175 89.990 177.340 ;
        RECT 89.780 176.805 90.060 177.175 ;
        RECT 88.870 175.980 89.130 176.300 ;
        RECT 86.570 174.620 86.830 174.940 ;
        RECT 86.630 174.455 86.770 174.620 ;
        RECT 86.560 174.085 86.840 174.455 ;
        RECT 87.950 174.280 88.210 174.600 ;
        RECT 88.010 173.540 88.150 174.280 ;
        RECT 87.090 173.400 88.150 173.540 ;
        RECT 87.090 172.900 87.230 173.400 ;
        RECT 87.030 172.580 87.290 172.900 ;
        RECT 88.410 172.240 88.670 172.560 ;
        RECT 87.950 171.560 88.210 171.880 ;
        RECT 88.010 170.375 88.150 171.560 ;
        RECT 85.640 170.005 85.920 170.375 ;
        RECT 87.940 170.005 88.220 170.375 ;
        RECT 84.730 168.840 84.990 169.160 ;
        RECT 84.730 167.140 84.990 167.460 ;
        RECT 84.790 165.420 84.930 167.140 ;
        RECT 85.710 166.780 85.850 170.005 ;
        RECT 88.470 167.800 88.610 172.240 ;
        RECT 88.930 170.860 89.070 175.980 ;
        RECT 89.330 174.620 89.590 174.940 ;
        RECT 89.390 172.900 89.530 174.620 ;
        RECT 89.850 174.600 89.990 176.805 ;
        RECT 90.310 175.280 90.450 178.360 ;
        RECT 90.250 174.960 90.510 175.280 ;
        RECT 89.790 174.280 90.050 174.600 ;
        RECT 91.230 173.580 91.370 180.400 ;
        RECT 92.550 179.720 92.810 180.040 ;
        RECT 92.610 177.660 92.750 179.720 ;
        RECT 94.450 177.740 94.590 187.200 ;
        RECT 95.830 185.820 95.970 193.660 ;
        RECT 96.290 192.620 96.430 196.380 ;
        RECT 97.210 193.980 97.350 199.440 ;
        RECT 97.150 193.660 97.410 193.980 ;
        RECT 97.670 193.380 97.810 202.760 ;
        RECT 98.530 202.160 98.790 202.480 ;
        RECT 98.070 199.780 98.330 200.100 ;
        RECT 98.130 197.575 98.270 199.780 ;
        RECT 98.060 197.205 98.340 197.575 ;
        RECT 98.590 197.380 98.730 202.160 ;
        RECT 100.430 202.140 100.570 203.270 ;
        RECT 101.350 203.160 101.490 203.325 ;
        RECT 100.820 202.645 101.100 203.015 ;
        RECT 101.290 202.840 101.550 203.160 ;
        RECT 100.370 201.820 100.630 202.140 ;
        RECT 98.990 200.460 99.250 200.780 ;
        RECT 99.050 200.100 99.190 200.460 ;
        RECT 100.890 200.440 101.030 202.645 ;
        RECT 100.830 200.120 101.090 200.440 ;
        RECT 98.990 199.780 99.250 200.100 ;
        RECT 99.155 198.225 100.695 198.595 ;
        RECT 101.280 198.140 101.560 198.255 ;
        RECT 101.810 198.140 101.950 204.290 ;
        RECT 102.270 203.500 102.410 205.310 ;
        RECT 102.670 205.220 102.930 205.540 ;
        RECT 102.210 203.180 102.470 203.500 ;
        RECT 99.450 197.740 99.710 198.060 ;
        RECT 100.890 198.000 101.950 198.140 ;
        RECT 99.510 197.575 99.650 197.740 ;
        RECT 98.530 197.060 98.790 197.380 ;
        RECT 99.440 197.205 99.720 197.575 ;
        RECT 99.510 194.660 99.650 197.205 ;
        RECT 100.890 194.660 101.030 198.000 ;
        RECT 101.280 197.885 101.560 198.000 ;
        RECT 101.290 197.060 101.550 197.380 ;
        RECT 98.530 194.570 98.790 194.660 ;
        RECT 98.530 194.430 99.190 194.570 ;
        RECT 98.530 194.340 98.790 194.430 ;
        RECT 99.050 194.060 99.190 194.430 ;
        RECT 99.450 194.340 99.710 194.660 ;
        RECT 100.830 194.340 101.090 194.660 ;
        RECT 99.910 194.060 100.170 194.320 ;
        RECT 99.050 194.000 100.170 194.060 ;
        RECT 98.530 193.660 98.790 193.980 ;
        RECT 99.050 193.920 100.110 194.000 ;
        RECT 100.830 193.660 101.090 193.980 ;
        RECT 96.750 193.240 97.810 193.380 ;
        RECT 98.070 193.320 98.330 193.640 ;
        RECT 96.230 192.300 96.490 192.620 ;
        RECT 96.230 191.620 96.490 191.940 ;
        RECT 96.290 188.200 96.430 191.620 ;
        RECT 96.230 187.880 96.490 188.200 ;
        RECT 95.770 185.500 96.030 185.820 ;
        RECT 95.300 184.285 95.580 184.655 ;
        RECT 95.370 183.440 95.510 184.285 ;
        RECT 94.850 183.120 95.110 183.440 ;
        RECT 95.310 183.120 95.570 183.440 ;
        RECT 94.910 181.060 95.050 183.120 ;
        RECT 95.830 182.760 95.970 185.500 ;
        RECT 96.750 184.460 96.890 193.240 ;
        RECT 98.130 192.815 98.270 193.320 ;
        RECT 98.060 192.445 98.340 192.815 ;
        RECT 97.150 190.940 97.410 191.260 ;
        RECT 98.070 190.940 98.330 191.260 ;
        RECT 97.210 189.900 97.350 190.940 ;
        RECT 97.150 189.580 97.410 189.900 ;
        RECT 97.600 189.045 97.880 189.415 ;
        RECT 97.610 188.900 97.870 189.045 ;
        RECT 97.610 186.860 97.870 187.180 ;
        RECT 97.150 185.160 97.410 185.480 ;
        RECT 96.690 184.140 96.950 184.460 ;
        RECT 97.210 183.780 97.350 185.160 ;
        RECT 97.670 184.655 97.810 186.860 ;
        RECT 98.130 185.820 98.270 190.940 ;
        RECT 98.590 189.560 98.730 193.660 ;
        RECT 99.155 192.785 100.695 193.155 ;
        RECT 100.370 191.850 100.630 191.940 ;
        RECT 99.050 191.710 100.630 191.850 ;
        RECT 98.530 189.240 98.790 189.560 ;
        RECT 99.050 188.790 99.190 191.710 ;
        RECT 100.370 191.620 100.630 191.710 ;
        RECT 100.890 191.260 101.030 193.660 ;
        RECT 100.830 190.940 101.090 191.260 ;
        RECT 100.360 189.725 100.640 190.095 ;
        RECT 98.590 188.650 99.190 188.790 ;
        RECT 98.070 185.500 98.330 185.820 ;
        RECT 97.600 184.285 97.880 184.655 ;
        RECT 98.590 184.370 98.730 188.650 ;
        RECT 100.430 188.200 100.570 189.725 ;
        RECT 100.370 187.880 100.630 188.200 ;
        RECT 99.155 187.345 100.695 187.715 ;
        RECT 100.890 187.180 101.030 190.940 ;
        RECT 100.830 186.860 101.090 187.180 ;
        RECT 99.910 186.580 100.170 186.840 ;
        RECT 99.910 186.520 100.570 186.580 ;
        RECT 99.970 186.440 100.570 186.520 ;
        RECT 99.450 185.335 99.710 185.480 ;
        RECT 99.440 184.965 99.720 185.335 ;
        RECT 99.910 185.160 100.170 185.480 ;
        RECT 97.610 184.140 97.870 184.285 ;
        RECT 98.590 184.230 99.190 184.370 ;
        RECT 96.230 183.460 96.490 183.780 ;
        RECT 97.150 183.460 97.410 183.780 ;
        RECT 97.600 183.605 97.880 183.975 ;
        RECT 98.520 183.605 98.800 183.975 ;
        RECT 99.050 183.780 99.190 184.230 ;
        RECT 99.970 184.120 100.110 185.160 ;
        RECT 99.910 183.800 100.170 184.120 ;
        RECT 96.290 182.760 96.430 183.460 ;
        RECT 96.690 183.120 96.950 183.440 ;
        RECT 95.770 182.440 96.030 182.760 ;
        RECT 96.230 182.440 96.490 182.760 ;
        RECT 96.750 181.740 96.890 183.120 ;
        RECT 96.690 181.420 96.950 181.740 ;
        RECT 94.850 180.740 95.110 181.060 ;
        RECT 94.910 179.020 95.050 180.740 ;
        RECT 97.210 180.720 97.350 183.460 ;
        RECT 96.690 180.400 96.950 180.720 ;
        RECT 97.150 180.400 97.410 180.720 ;
        RECT 94.850 178.700 95.110 179.020 ;
        RECT 91.630 177.340 91.890 177.660 ;
        RECT 92.550 177.340 92.810 177.660 ;
        RECT 94.450 177.600 95.970 177.740 ;
        RECT 96.230 177.680 96.490 178.000 ;
        RECT 91.690 176.300 91.830 177.340 ;
        RECT 95.310 177.000 95.570 177.320 ;
        RECT 91.630 175.980 91.890 176.300 ;
        RECT 92.080 176.125 92.360 176.495 ;
        RECT 92.090 175.980 92.350 176.125 ;
        RECT 92.090 174.620 92.350 174.940 ;
        RECT 90.710 173.260 90.970 173.580 ;
        RECT 91.170 173.260 91.430 173.580 ;
        RECT 89.330 172.580 89.590 172.900 ;
        RECT 89.790 172.580 90.050 172.900 ;
        RECT 89.390 170.860 89.530 172.580 ;
        RECT 89.850 172.415 89.990 172.580 ;
        RECT 89.780 172.045 90.060 172.415 ;
        RECT 90.250 171.900 90.510 172.220 ;
        RECT 88.870 170.540 89.130 170.860 ;
        RECT 89.330 170.540 89.590 170.860 ;
        RECT 88.870 167.820 89.130 168.140 ;
        RECT 88.410 167.480 88.670 167.800 ;
        RECT 88.930 167.460 89.070 167.820 ;
        RECT 88.870 167.140 89.130 167.460 ;
        RECT 86.110 166.800 86.370 167.120 ;
        RECT 85.650 166.460 85.910 166.780 ;
        RECT 84.730 165.100 84.990 165.420 ;
        RECT 84.270 162.380 84.530 162.700 ;
        RECT 86.170 162.020 86.310 166.800 ;
        RECT 87.030 164.080 87.290 164.400 ;
        RECT 86.570 163.400 86.830 163.720 ;
        RECT 86.630 162.020 86.770 163.400 ;
        RECT 86.110 161.700 86.370 162.020 ;
        RECT 86.570 161.700 86.830 162.020 ;
        RECT 83.810 159.320 84.070 159.640 ;
        RECT 82.890 158.640 83.150 158.960 ;
        RECT 86.630 158.280 86.770 161.700 ;
        RECT 87.090 159.980 87.230 164.080 ;
        RECT 89.390 162.700 89.530 170.540 ;
        RECT 90.310 170.180 90.450 171.900 ;
        RECT 90.770 170.860 90.910 173.260 ;
        RECT 92.150 172.900 92.290 174.620 ;
        RECT 95.370 174.600 95.510 177.000 ;
        RECT 95.830 175.960 95.970 177.600 ;
        RECT 96.290 176.300 96.430 177.680 ;
        RECT 96.230 175.980 96.490 176.300 ;
        RECT 95.770 175.640 96.030 175.960 ;
        RECT 96.220 175.445 96.500 175.815 ;
        RECT 95.310 174.280 95.570 174.600 ;
        RECT 95.370 173.580 95.510 174.280 ;
        RECT 92.550 173.260 92.810 173.580 ;
        RECT 95.310 173.260 95.570 173.580 ;
        RECT 95.770 173.260 96.030 173.580 ;
        RECT 91.170 172.580 91.430 172.900 ;
        RECT 92.090 172.580 92.350 172.900 ;
        RECT 90.710 170.540 90.970 170.860 ;
        RECT 90.250 169.860 90.510 170.180 ;
        RECT 91.230 167.460 91.370 172.580 ;
        RECT 92.610 170.260 92.750 173.260 ;
        RECT 93.930 172.580 94.190 172.900 ;
        RECT 94.390 172.580 94.650 172.900 ;
        RECT 93.010 172.240 93.270 172.560 ;
        RECT 92.150 170.120 92.750 170.260 ;
        RECT 91.630 169.520 91.890 169.840 ;
        RECT 91.170 167.140 91.430 167.460 ;
        RECT 90.250 167.030 90.510 167.120 ;
        RECT 89.850 166.890 90.510 167.030 ;
        RECT 89.850 164.740 89.990 166.890 ;
        RECT 90.250 166.800 90.510 166.890 ;
        RECT 90.250 166.120 90.510 166.440 ;
        RECT 89.790 164.420 90.050 164.740 ;
        RECT 89.330 162.380 89.590 162.700 ;
        RECT 89.850 161.930 89.990 164.420 ;
        RECT 90.310 164.400 90.450 166.120 ;
        RECT 91.230 165.420 91.370 167.140 ;
        RECT 91.690 166.975 91.830 169.520 ;
        RECT 92.150 169.160 92.290 170.120 ;
        RECT 92.550 169.520 92.810 169.840 ;
        RECT 92.090 168.840 92.350 169.160 ;
        RECT 92.610 168.140 92.750 169.520 ;
        RECT 92.550 167.820 92.810 168.140 ;
        RECT 93.070 167.460 93.210 172.240 ;
        RECT 93.470 171.900 93.730 172.220 ;
        RECT 93.530 169.500 93.670 171.900 ;
        RECT 93.990 170.180 94.130 172.580 ;
        RECT 94.450 171.055 94.590 172.580 ;
        RECT 95.830 172.560 95.970 173.260 ;
        RECT 94.850 172.240 95.110 172.560 ;
        RECT 95.770 172.470 96.030 172.560 ;
        RECT 95.370 172.330 96.030 172.470 ;
        RECT 94.380 170.685 94.660 171.055 ;
        RECT 94.910 170.430 95.050 172.240 ;
        RECT 94.450 170.290 95.050 170.430 ;
        RECT 93.930 169.860 94.190 170.180 ;
        RECT 94.450 169.840 94.590 170.290 ;
        RECT 94.390 169.520 94.650 169.840 ;
        RECT 93.470 169.180 93.730 169.500 ;
        RECT 94.840 169.325 95.120 169.695 ;
        RECT 94.910 167.460 95.050 169.325 ;
        RECT 93.010 167.140 93.270 167.460 ;
        RECT 94.850 167.140 95.110 167.460 ;
        RECT 91.620 166.605 91.900 166.975 ;
        RECT 92.090 166.800 92.350 167.120 ;
        RECT 91.630 166.460 91.890 166.605 ;
        RECT 91.170 165.100 91.430 165.420 ;
        RECT 90.250 164.080 90.510 164.400 ;
        RECT 91.630 164.080 91.890 164.400 ;
        RECT 91.690 162.100 91.830 164.080 ;
        RECT 92.150 162.700 92.290 166.800 ;
        RECT 92.540 165.925 92.820 166.295 ;
        RECT 92.610 162.700 92.750 165.925 ;
        RECT 93.070 162.700 93.210 167.140 ;
        RECT 93.470 166.800 93.730 167.120 ;
        RECT 93.530 165.420 93.670 166.800 ;
        RECT 93.470 165.100 93.730 165.420 ;
        RECT 95.370 164.400 95.510 172.330 ;
        RECT 95.770 172.240 96.030 172.330 ;
        RECT 95.770 166.120 96.030 166.440 ;
        RECT 95.830 165.420 95.970 166.120 ;
        RECT 95.770 165.100 96.030 165.420 ;
        RECT 95.310 164.080 95.570 164.400 ;
        RECT 94.850 163.575 95.110 163.720 ;
        RECT 94.840 163.205 95.120 163.575 ;
        RECT 92.090 162.380 92.350 162.700 ;
        RECT 92.550 162.380 92.810 162.700 ;
        RECT 93.010 162.380 93.270 162.700 ;
        RECT 95.770 162.380 96.030 162.700 ;
        RECT 93.070 162.100 93.210 162.380 ;
        RECT 90.250 161.930 90.510 162.020 ;
        RECT 89.850 161.790 90.510 161.930 ;
        RECT 88.410 161.020 88.670 161.340 ;
        RECT 88.470 159.980 88.610 161.020 ;
        RECT 87.030 159.660 87.290 159.980 ;
        RECT 88.410 159.890 88.670 159.980 ;
        RECT 88.010 159.750 88.670 159.890 ;
        RECT 88.010 159.300 88.150 159.750 ;
        RECT 88.410 159.660 88.670 159.750 ;
        RECT 89.850 159.740 89.990 161.790 ;
        RECT 90.250 161.700 90.510 161.790 ;
        RECT 91.170 161.700 91.430 162.020 ;
        RECT 91.690 161.960 93.210 162.100 ;
        RECT 94.380 161.845 94.660 162.215 ;
        RECT 94.390 161.700 94.650 161.845 ;
        RECT 90.710 160.680 90.970 161.000 ;
        RECT 89.390 159.600 89.990 159.740 ;
        RECT 87.950 158.980 88.210 159.300 ;
        RECT 87.030 158.640 87.290 158.960 ;
        RECT 88.410 158.640 88.670 158.960 ;
        RECT 82.890 157.960 83.150 158.280 ;
        RECT 86.570 157.960 86.830 158.280 ;
        RECT 82.950 154.540 83.090 157.960 ;
        RECT 85.190 156.600 85.450 156.920 ;
        RECT 84.720 155.725 85.000 156.095 ;
        RECT 83.810 155.240 84.070 155.560 ;
        RECT 84.270 155.240 84.530 155.560 ;
        RECT 82.430 154.220 82.690 154.540 ;
        RECT 82.890 154.220 83.150 154.540 ;
        RECT 83.350 153.880 83.610 154.200 ;
        RECT 82.890 152.860 83.150 153.180 ;
        RECT 81.970 152.520 82.230 152.840 ;
        RECT 79.670 148.100 79.930 148.420 ;
        RECT 81.510 148.100 81.770 148.420 ;
        RECT 79.720 146.545 81.260 146.915 ;
        RECT 79.210 144.360 79.470 144.680 ;
        RECT 78.750 143.340 79.010 143.660 ;
        RECT 76.910 141.980 77.170 142.300 ;
        RECT 77.830 141.980 78.090 142.300 ;
        RECT 74.610 141.640 74.870 141.960 ;
        RECT 74.670 140.940 74.810 141.640 ;
        RECT 74.610 140.620 74.870 140.940 ;
        RECT 75.070 138.920 75.330 139.240 ;
        RECT 74.610 136.880 74.870 137.200 ;
        RECT 74.150 129.740 74.410 130.060 ;
        RECT 72.310 129.060 72.570 129.380 ;
        RECT 72.770 128.720 73.030 129.040 ;
        RECT 59.890 126.000 60.150 126.320 ;
        RECT 70.010 126.000 70.270 126.320 ;
        RECT 70.930 126.175 71.190 126.320 ;
        RECT 67.710 125.660 67.970 125.980 ;
        RECT 53.910 125.550 54.170 125.640 ;
        RECT 53.050 125.410 54.170 125.550 ;
        RECT 53.910 125.320 54.170 125.410 ;
        RECT 48.450 125.100 49.970 125.240 ;
        RECT 46.090 124.300 46.350 124.620 ;
        RECT 48.450 123.940 48.590 125.100 ;
        RECT 67.770 124.280 67.910 125.660 ;
        RECT 67.710 123.960 67.970 124.280 ;
        RECT 70.070 123.940 70.210 126.000 ;
        RECT 70.920 125.805 71.200 126.175 ;
        RECT 70.990 125.240 71.130 125.805 ;
        RECT 70.990 125.100 71.590 125.240 ;
        RECT 71.450 123.940 71.590 125.100 ;
        RECT 43.330 123.620 43.590 123.940 ;
        RECT 48.390 123.620 48.650 123.940 ;
        RECT 70.010 123.620 70.270 123.940 ;
        RECT 70.930 123.620 71.190 123.940 ;
        RECT 71.390 123.620 71.650 123.940 ;
        RECT 70.990 123.340 71.130 123.620 ;
        RECT 72.830 123.340 72.970 128.720 ;
        RECT 74.670 127.340 74.810 136.880 ;
        RECT 75.130 132.440 75.270 138.920 ;
        RECT 76.450 137.220 76.710 137.540 ;
        RECT 76.510 135.500 76.650 137.220 ;
        RECT 77.890 137.055 78.030 141.980 ;
        RECT 79.270 140.600 79.410 144.360 ;
        RECT 81.510 141.640 81.770 141.960 ;
        RECT 79.720 141.105 81.260 141.475 ;
        RECT 79.210 140.280 79.470 140.600 ;
        RECT 81.570 139.920 81.710 141.640 ;
        RECT 80.590 139.600 80.850 139.920 ;
        RECT 81.510 139.600 81.770 139.920 ;
        RECT 80.650 137.880 80.790 139.600 ;
        RECT 81.040 138.045 81.320 138.415 ;
        RECT 80.590 137.560 80.850 137.880 ;
        RECT 81.110 137.200 81.250 138.045 ;
        RECT 78.750 137.055 79.010 137.200 ;
        RECT 81.050 137.110 81.310 137.200 ;
        RECT 77.820 136.685 78.100 137.055 ;
        RECT 78.740 136.685 79.020 137.055 ;
        RECT 79.270 136.970 81.310 137.110 ;
        RECT 76.910 136.200 77.170 136.520 ;
        RECT 76.970 135.500 77.110 136.200 ;
        RECT 77.360 136.005 77.640 136.375 ;
        RECT 77.430 135.500 77.570 136.005 ;
        RECT 75.990 135.180 76.250 135.500 ;
        RECT 76.450 135.180 76.710 135.500 ;
        RECT 76.910 135.180 77.170 135.500 ;
        RECT 77.370 135.180 77.630 135.500 ;
        RECT 78.740 135.325 79.020 135.695 ;
        RECT 78.750 135.180 79.010 135.325 ;
        RECT 75.530 134.160 75.790 134.480 ;
        RECT 75.070 132.120 75.330 132.440 ;
        RECT 75.130 131.760 75.270 132.120 ;
        RECT 75.590 131.760 75.730 134.160 ;
        RECT 76.050 132.180 76.190 135.180 ;
        RECT 79.270 134.900 79.410 136.970 ;
        RECT 81.050 136.880 81.310 136.970 ;
        RECT 79.720 135.665 81.260 136.035 ;
        RECT 76.970 134.820 79.410 134.900 ;
        RECT 76.910 134.760 79.410 134.820 ;
        RECT 76.910 134.500 77.170 134.760 ;
        RECT 76.050 132.040 76.650 132.180 ;
        RECT 75.070 131.440 75.330 131.760 ;
        RECT 75.530 131.440 75.790 131.760 ;
        RECT 75.990 131.100 76.250 131.420 ;
        RECT 75.530 130.760 75.790 131.080 ;
        RECT 75.590 129.460 75.730 130.760 ;
        RECT 76.050 130.060 76.190 131.100 ;
        RECT 76.510 130.060 76.650 132.040 ;
        RECT 76.970 131.760 77.110 134.500 ;
        RECT 81.050 134.160 81.310 134.480 ;
        RECT 77.830 133.820 78.090 134.140 ;
        RECT 78.290 133.820 78.550 134.140 ;
        RECT 76.910 131.440 77.170 131.760 ;
        RECT 75.990 129.740 76.250 130.060 ;
        RECT 76.450 129.740 76.710 130.060 ;
        RECT 75.590 129.320 76.190 129.460 ;
        RECT 74.610 127.020 74.870 127.340 ;
        RECT 76.050 123.940 76.190 129.320 ;
        RECT 76.510 126.660 76.650 129.740 ;
        RECT 76.910 129.060 77.170 129.380 ;
        RECT 76.970 127.340 77.110 129.060 ;
        RECT 77.370 128.040 77.630 128.360 ;
        RECT 77.430 127.340 77.570 128.040 ;
        RECT 76.910 127.020 77.170 127.340 ;
        RECT 77.370 127.020 77.630 127.340 ;
        RECT 76.450 126.340 76.710 126.660 ;
        RECT 76.970 123.940 77.110 127.020 ;
        RECT 77.890 126.660 78.030 133.820 ;
        RECT 78.350 132.780 78.490 133.820 ;
        RECT 78.290 132.460 78.550 132.780 ;
        RECT 80.130 132.460 80.390 132.780 ;
        RECT 80.190 131.760 80.330 132.460 ;
        RECT 80.130 131.440 80.390 131.760 ;
        RECT 81.110 131.420 81.250 134.160 ;
        RECT 81.570 132.100 81.710 139.600 ;
        RECT 81.510 131.780 81.770 132.100 ;
        RECT 81.050 131.100 81.310 131.420 ;
        RECT 79.720 130.225 81.260 130.595 ;
        RECT 77.830 126.340 78.090 126.660 ;
        RECT 78.290 126.000 78.550 126.320 ;
        RECT 79.210 126.000 79.470 126.320 ;
        RECT 78.350 124.620 78.490 126.000 ;
        RECT 78.290 124.300 78.550 124.620 ;
        RECT 79.270 124.280 79.410 126.000 ;
        RECT 82.030 125.980 82.170 152.520 ;
        RECT 82.950 151.820 83.090 152.860 ;
        RECT 82.890 151.500 83.150 151.820 ;
        RECT 83.410 151.480 83.550 153.880 ;
        RECT 83.870 153.520 84.010 155.240 ;
        RECT 84.330 153.860 84.470 155.240 ;
        RECT 84.790 153.860 84.930 155.725 ;
        RECT 84.270 153.540 84.530 153.860 ;
        RECT 84.730 153.540 84.990 153.860 ;
        RECT 83.810 153.200 84.070 153.520 ;
        RECT 83.810 151.500 84.070 151.820 ;
        RECT 83.350 151.160 83.610 151.480 ;
        RECT 82.430 149.800 82.690 150.120 ;
        RECT 82.490 148.760 82.630 149.800 ;
        RECT 82.430 148.440 82.690 148.760 ;
        RECT 82.490 145.360 82.630 148.440 ;
        RECT 83.870 147.400 84.010 151.500 ;
        RECT 84.330 148.420 84.470 153.540 ;
        RECT 85.250 151.480 85.390 156.600 ;
        RECT 87.090 154.540 87.230 158.640 ;
        RECT 88.470 154.540 88.610 158.640 ;
        RECT 89.390 158.280 89.530 159.600 ;
        RECT 88.870 157.960 89.130 158.280 ;
        RECT 89.330 157.960 89.590 158.280 ;
        RECT 88.930 157.260 89.070 157.960 ;
        RECT 88.870 156.940 89.130 157.260 ;
        RECT 87.030 154.220 87.290 154.540 ;
        RECT 88.410 154.220 88.670 154.540 ;
        RECT 90.770 153.940 90.910 160.680 ;
        RECT 91.230 159.980 91.370 161.700 ;
        RECT 94.850 160.680 95.110 161.000 ;
        RECT 91.170 159.660 91.430 159.980 ;
        RECT 93.010 158.640 93.270 158.960 ;
        RECT 92.550 157.960 92.810 158.280 ;
        RECT 92.090 156.260 92.350 156.580 ;
        RECT 92.150 155.900 92.290 156.260 ;
        RECT 92.090 155.580 92.350 155.900 ;
        RECT 89.850 153.800 90.910 153.940 ;
        RECT 89.850 153.520 89.990 153.800 ;
        RECT 89.790 153.200 90.050 153.520 ;
        RECT 90.250 153.200 90.510 153.520 ;
        RECT 89.790 152.520 90.050 152.840 ;
        RECT 85.190 151.160 85.450 151.480 ;
        RECT 85.250 150.800 85.390 151.160 ;
        RECT 85.190 150.480 85.450 150.800 ;
        RECT 87.950 150.480 88.210 150.800 ;
        RECT 88.410 150.480 88.670 150.800 ;
        RECT 84.270 148.100 84.530 148.420 ;
        RECT 83.810 147.080 84.070 147.400 ;
        RECT 84.730 147.080 84.990 147.400 ;
        RECT 82.880 145.525 83.160 145.895 ;
        RECT 82.430 145.040 82.690 145.360 ;
        RECT 82.950 144.535 83.090 145.525 ;
        RECT 82.880 144.165 83.160 144.535 ;
        RECT 84.270 144.360 84.530 144.680 ;
        RECT 83.350 142.660 83.610 142.980 ;
        RECT 82.430 141.640 82.690 141.960 ;
        RECT 82.490 136.520 82.630 141.640 ;
        RECT 82.430 136.200 82.690 136.520 ;
        RECT 82.880 135.325 83.160 135.695 ;
        RECT 82.950 133.800 83.090 135.325 ;
        RECT 83.410 134.220 83.550 142.660 ;
        RECT 83.810 137.900 84.070 138.220 ;
        RECT 83.870 135.500 84.010 137.900 ;
        RECT 84.330 137.880 84.470 144.360 ;
        RECT 84.790 143.855 84.930 147.080 ;
        RECT 87.490 145.950 87.750 146.040 ;
        RECT 88.010 145.950 88.150 150.480 ;
        RECT 88.470 148.080 88.610 150.480 ;
        RECT 89.330 148.100 89.590 148.420 ;
        RECT 88.410 147.760 88.670 148.080 ;
        RECT 87.490 145.810 88.150 145.950 ;
        RECT 87.490 145.720 87.750 145.810 ;
        RECT 88.410 145.380 88.670 145.700 ;
        RECT 84.720 143.485 85.000 143.855 ;
        RECT 88.470 143.660 88.610 145.380 ;
        RECT 88.870 144.360 89.130 144.680 ;
        RECT 88.930 143.660 89.070 144.360 ;
        RECT 89.390 143.660 89.530 148.100 ;
        RECT 89.850 146.290 89.990 152.520 ;
        RECT 90.310 149.100 90.450 153.200 ;
        RECT 90.250 148.780 90.510 149.100 ;
        RECT 90.770 148.080 90.910 153.800 ;
        RECT 92.090 152.860 92.350 153.180 ;
        RECT 91.170 150.820 91.430 151.140 ;
        RECT 91.230 149.295 91.370 150.820 ;
        RECT 91.160 148.925 91.440 149.295 ;
        RECT 90.710 147.760 90.970 148.080 ;
        RECT 91.630 147.760 91.890 148.080 ;
        RECT 89.850 146.150 91.370 146.290 ;
        RECT 90.250 145.380 90.510 145.700 ;
        RECT 89.790 144.700 90.050 145.020 ;
        RECT 88.410 143.340 88.670 143.660 ;
        RECT 88.870 143.340 89.130 143.660 ;
        RECT 89.330 143.340 89.590 143.660 ;
        RECT 85.190 141.980 85.450 142.300 ;
        RECT 85.250 140.260 85.390 141.980 ;
        RECT 89.850 140.260 89.990 144.700 ;
        RECT 90.310 143.660 90.450 145.380 ;
        RECT 91.230 145.360 91.370 146.150 ;
        RECT 91.690 146.040 91.830 147.760 ;
        RECT 91.630 145.720 91.890 146.040 ;
        RECT 92.150 145.360 92.290 152.860 ;
        RECT 92.610 148.080 92.750 157.960 ;
        RECT 93.070 156.240 93.210 158.640 ;
        RECT 93.010 155.920 93.270 156.240 ;
        RECT 93.070 151.140 93.210 155.920 ;
        RECT 93.470 155.580 93.730 155.900 ;
        RECT 93.010 150.820 93.270 151.140 ;
        RECT 93.530 148.420 93.670 155.580 ;
        RECT 94.910 151.480 95.050 160.680 ;
        RECT 95.830 158.960 95.970 162.380 ;
        RECT 96.290 161.000 96.430 175.445 ;
        RECT 96.750 173.540 96.890 180.400 ;
        RECT 97.150 177.000 97.410 177.320 ;
        RECT 97.210 174.940 97.350 177.000 ;
        RECT 97.670 175.960 97.810 183.605 ;
        RECT 98.590 182.615 98.730 183.605 ;
        RECT 98.990 183.460 99.250 183.780 ;
        RECT 100.430 182.670 100.570 186.440 ;
        RECT 100.830 185.840 101.090 186.160 ;
        RECT 100.890 183.440 101.030 185.840 ;
        RECT 100.830 183.120 101.090 183.440 ;
        RECT 98.520 182.245 98.800 182.615 ;
        RECT 100.430 182.530 101.030 182.670 ;
        RECT 99.155 181.905 100.695 182.275 ;
        RECT 100.890 180.380 101.030 182.530 ;
        RECT 100.830 180.060 101.090 180.380 ;
        RECT 98.070 178.020 98.330 178.340 ;
        RECT 98.520 178.165 98.800 178.535 ;
        RECT 101.350 178.340 101.490 197.060 ;
        RECT 102.270 192.815 102.410 203.180 ;
        RECT 102.730 199.760 102.870 205.220 ;
        RECT 103.130 204.880 103.390 205.200 ;
        RECT 103.190 203.160 103.330 204.880 ;
        RECT 103.590 203.180 103.850 203.500 ;
        RECT 103.130 202.840 103.390 203.160 ;
        RECT 102.670 199.440 102.930 199.760 ;
        RECT 102.660 198.565 102.940 198.935 ;
        RECT 102.730 197.040 102.870 198.565 ;
        RECT 103.190 197.720 103.330 202.840 ;
        RECT 103.650 200.100 103.790 203.180 ;
        RECT 104.050 202.840 104.310 203.160 ;
        RECT 104.110 200.440 104.250 202.840 ;
        RECT 104.050 200.120 104.310 200.440 ;
        RECT 103.590 199.780 103.850 200.100 ;
        RECT 103.130 197.400 103.390 197.720 ;
        RECT 102.670 196.720 102.930 197.040 ;
        RECT 102.730 194.660 102.870 196.720 ;
        RECT 103.120 196.525 103.400 196.895 ;
        RECT 103.190 195.340 103.330 196.525 ;
        RECT 103.130 195.020 103.390 195.340 ;
        RECT 102.670 194.340 102.930 194.660 ;
        RECT 103.650 193.980 103.790 199.780 ;
        RECT 104.050 199.440 104.310 199.760 ;
        RECT 104.110 197.040 104.250 199.440 ;
        RECT 104.050 196.720 104.310 197.040 ;
        RECT 103.590 193.660 103.850 193.980 ;
        RECT 102.200 192.445 102.480 192.815 ;
        RECT 101.750 190.940 102.010 191.260 ;
        RECT 101.810 190.095 101.950 190.940 ;
        RECT 101.740 189.725 102.020 190.095 ;
        RECT 102.270 188.880 102.410 192.445 ;
        RECT 104.110 191.940 104.250 196.720 ;
        RECT 104.570 194.660 104.710 205.900 ;
        RECT 105.950 205.540 106.090 210.660 ;
        RECT 105.890 205.220 106.150 205.540 ;
        RECT 105.890 204.540 106.150 204.860 ;
        RECT 104.970 204.200 105.230 204.520 ;
        RECT 105.030 201.800 105.170 204.200 ;
        RECT 104.970 201.480 105.230 201.800 ;
        RECT 104.970 199.440 105.230 199.760 ;
        RECT 105.030 198.060 105.170 199.440 ;
        RECT 104.970 197.740 105.230 198.060 ;
        RECT 105.430 196.380 105.690 196.700 ;
        RECT 104.960 195.845 105.240 196.215 ;
        RECT 104.510 194.340 104.770 194.660 ;
        RECT 104.510 192.300 104.770 192.620 ;
        RECT 104.050 191.620 104.310 191.940 ;
        RECT 103.130 191.510 103.390 191.600 ;
        RECT 102.730 191.370 103.390 191.510 ;
        RECT 102.730 188.880 102.870 191.370 ;
        RECT 103.130 191.280 103.390 191.370 ;
        RECT 103.580 191.085 103.860 191.455 ;
        RECT 104.570 191.340 104.710 192.300 ;
        RECT 105.030 191.940 105.170 195.845 ;
        RECT 104.970 191.620 105.230 191.940 ;
        RECT 104.110 191.200 104.710 191.340 ;
        RECT 103.130 188.900 103.390 189.220 ;
        RECT 102.210 188.560 102.470 188.880 ;
        RECT 102.670 188.560 102.930 188.880 ;
        RECT 103.190 188.055 103.330 188.900 ;
        RECT 103.120 187.685 103.400 188.055 ;
        RECT 102.660 187.005 102.940 187.375 ;
        RECT 102.210 186.520 102.470 186.840 ;
        RECT 101.750 185.160 102.010 185.480 ;
        RECT 101.810 183.440 101.950 185.160 ;
        RECT 102.270 183.780 102.410 186.520 ;
        RECT 102.210 183.460 102.470 183.780 ;
        RECT 101.750 183.120 102.010 183.440 ;
        RECT 101.810 181.740 101.950 183.120 ;
        RECT 102.210 182.780 102.470 183.100 ;
        RECT 102.270 181.740 102.410 182.780 ;
        RECT 101.750 181.420 102.010 181.740 ;
        RECT 102.210 181.420 102.470 181.740 ;
        RECT 102.730 181.140 102.870 187.005 ;
        RECT 103.190 185.820 103.330 187.685 ;
        RECT 103.650 186.015 103.790 191.085 ;
        RECT 104.110 188.540 104.250 191.200 ;
        RECT 104.970 190.600 105.230 190.920 ;
        RECT 105.030 189.220 105.170 190.600 ;
        RECT 104.970 189.130 105.230 189.220 ;
        RECT 104.570 188.990 105.230 189.130 ;
        RECT 104.050 188.220 104.310 188.540 ;
        RECT 104.570 186.500 104.710 188.990 ;
        RECT 104.970 188.900 105.230 188.990 ;
        RECT 104.510 186.180 104.770 186.500 ;
        RECT 103.130 185.500 103.390 185.820 ;
        RECT 103.580 185.645 103.860 186.015 ;
        RECT 104.970 185.840 105.230 186.160 ;
        RECT 104.510 185.160 104.770 185.480 ;
        RECT 103.130 182.440 103.390 182.760 ;
        RECT 103.190 181.740 103.330 182.440 ;
        RECT 103.130 181.420 103.390 181.740 ;
        RECT 103.590 181.420 103.850 181.740 ;
        RECT 102.270 181.000 102.870 181.140 ;
        RECT 102.270 178.340 102.410 181.000 ;
        RECT 102.670 178.700 102.930 179.020 ;
        RECT 97.610 175.640 97.870 175.960 ;
        RECT 97.150 174.620 97.410 174.940 ;
        RECT 98.130 174.600 98.270 178.020 ;
        RECT 98.070 174.280 98.330 174.600 ;
        RECT 98.590 173.540 98.730 178.165 ;
        RECT 101.290 178.020 101.550 178.340 ;
        RECT 102.210 178.020 102.470 178.340 ;
        RECT 100.830 177.340 101.090 177.660 ;
        RECT 99.155 176.465 100.695 176.835 ;
        RECT 100.890 176.300 101.030 177.340 ;
        RECT 101.350 177.175 101.490 178.020 ;
        RECT 101.280 176.805 101.560 177.175 ;
        RECT 101.750 177.000 102.010 177.320 ;
        RECT 100.830 175.980 101.090 176.300 ;
        RECT 100.370 175.815 100.630 175.960 ;
        RECT 100.360 175.445 100.640 175.815 ;
        RECT 101.810 175.620 101.950 177.000 ;
        RECT 102.730 176.300 102.870 178.700 ;
        RECT 103.650 178.340 103.790 181.420 ;
        RECT 104.570 180.040 104.710 185.160 ;
        RECT 105.030 184.460 105.170 185.840 ;
        RECT 104.970 184.140 105.230 184.460 ;
        RECT 104.970 180.060 105.230 180.380 ;
        RECT 104.510 179.720 104.770 180.040 ;
        RECT 104.050 178.360 104.310 178.680 ;
        RECT 103.590 178.020 103.850 178.340 ;
        RECT 102.670 175.980 102.930 176.300 ;
        RECT 101.750 175.300 102.010 175.620 ;
        RECT 102.200 174.765 102.480 175.135 ;
        RECT 103.130 174.960 103.390 175.280 ;
        RECT 96.750 173.400 97.350 173.540 ;
        RECT 96.690 169.180 96.950 169.500 ;
        RECT 96.750 166.440 96.890 169.180 ;
        RECT 96.690 166.120 96.950 166.440 ;
        RECT 96.750 165.080 96.890 166.120 ;
        RECT 96.690 164.760 96.950 165.080 ;
        RECT 96.680 163.460 96.960 163.575 ;
        RECT 97.210 163.460 97.350 173.400 ;
        RECT 98.130 173.400 98.730 173.540 ;
        RECT 100.830 173.490 101.090 173.580 ;
        RECT 97.610 169.860 97.870 170.180 ;
        RECT 97.670 163.720 97.810 169.860 ;
        RECT 96.680 163.320 97.350 163.460 ;
        RECT 97.610 163.400 97.870 163.720 ;
        RECT 96.680 163.205 96.960 163.320 ;
        RECT 97.150 162.380 97.410 162.700 ;
        RECT 96.690 161.360 96.950 161.680 ;
        RECT 96.230 160.680 96.490 161.000 ;
        RECT 95.770 158.640 96.030 158.960 ;
        RECT 96.230 158.640 96.490 158.960 ;
        RECT 95.760 156.405 96.040 156.775 ;
        RECT 95.830 154.540 95.970 156.405 ;
        RECT 96.290 156.240 96.430 158.640 ;
        RECT 96.750 158.280 96.890 161.360 ;
        RECT 96.690 157.960 96.950 158.280 ;
        RECT 96.230 155.920 96.490 156.240 ;
        RECT 95.770 154.220 96.030 154.540 ;
        RECT 96.290 154.200 96.430 155.920 ;
        RECT 95.760 153.685 96.040 154.055 ;
        RECT 96.230 153.880 96.490 154.200 ;
        RECT 94.850 151.160 95.110 151.480 ;
        RECT 95.830 150.800 95.970 153.685 ;
        RECT 96.680 150.965 96.960 151.335 ;
        RECT 96.690 150.820 96.950 150.965 ;
        RECT 95.310 150.480 95.570 150.800 ;
        RECT 95.770 150.480 96.030 150.800 ;
        RECT 93.470 148.100 93.730 148.420 ;
        RECT 94.850 148.100 95.110 148.420 ;
        RECT 92.550 147.760 92.810 148.080 ;
        RECT 90.710 145.040 90.970 145.360 ;
        RECT 91.170 145.040 91.430 145.360 ;
        RECT 92.090 145.040 92.350 145.360 ;
        RECT 90.250 143.340 90.510 143.660 ;
        RECT 90.770 143.320 90.910 145.040 ;
        RECT 90.710 143.000 90.970 143.320 ;
        RECT 92.150 143.060 92.290 145.040 ;
        RECT 94.910 145.020 95.050 148.100 ;
        RECT 94.390 144.700 94.650 145.020 ;
        RECT 94.850 144.700 95.110 145.020 ;
        RECT 93.010 144.360 93.270 144.680 ;
        RECT 93.070 143.660 93.210 144.360 ;
        RECT 93.010 143.340 93.270 143.660 ;
        RECT 85.190 139.940 85.450 140.260 ;
        RECT 88.870 139.940 89.130 140.260 ;
        RECT 89.790 139.940 90.050 140.260 ;
        RECT 90.770 140.170 90.910 143.000 ;
        RECT 92.150 142.920 92.750 143.060 ;
        RECT 92.610 142.640 92.750 142.920 ;
        RECT 92.090 142.320 92.350 142.640 ;
        RECT 92.550 142.320 92.810 142.640 ;
        RECT 91.170 141.980 91.430 142.300 ;
        RECT 91.630 141.980 91.890 142.300 ;
        RECT 91.230 140.940 91.370 141.980 ;
        RECT 91.170 140.620 91.430 140.940 ;
        RECT 91.170 140.170 91.430 140.260 ;
        RECT 90.770 140.030 91.430 140.170 ;
        RECT 91.170 139.940 91.430 140.030 ;
        RECT 84.270 137.560 84.530 137.880 ;
        RECT 84.330 135.500 84.470 137.560 ;
        RECT 85.250 137.200 85.390 139.940 ;
        RECT 85.650 137.220 85.910 137.540 ;
        RECT 85.190 136.880 85.450 137.200 ;
        RECT 83.810 135.180 84.070 135.500 ;
        RECT 84.270 135.180 84.530 135.500 ;
        RECT 83.410 134.080 84.010 134.220 ;
        RECT 82.890 133.480 83.150 133.800 ;
        RECT 83.350 133.480 83.610 133.800 ;
        RECT 83.410 132.100 83.550 133.480 ;
        RECT 83.350 131.780 83.610 132.100 ;
        RECT 83.350 130.760 83.610 131.080 ;
        RECT 83.410 128.360 83.550 130.760 ;
        RECT 83.350 128.040 83.610 128.360 ;
        RECT 83.410 127.340 83.550 128.040 ;
        RECT 83.350 127.020 83.610 127.340 ;
        RECT 83.870 126.320 84.010 134.080 ;
        RECT 85.250 133.800 85.390 136.880 ;
        RECT 85.710 135.500 85.850 137.220 ;
        RECT 86.110 136.200 86.370 136.520 ;
        RECT 85.650 135.180 85.910 135.500 ;
        RECT 86.170 135.160 86.310 136.200 ;
        RECT 88.930 135.500 89.070 139.940 ;
        RECT 90.250 139.600 90.510 139.920 ;
        RECT 90.310 137.540 90.450 139.600 ;
        RECT 91.690 138.415 91.830 141.980 ;
        RECT 91.620 138.045 91.900 138.415 ;
        RECT 92.150 137.540 92.290 142.320 ;
        RECT 94.450 140.600 94.590 144.700 ;
        RECT 94.390 140.280 94.650 140.600 ;
        RECT 94.850 139.260 95.110 139.580 ;
        RECT 90.250 137.220 90.510 137.540 ;
        RECT 92.090 137.220 92.350 137.540 ;
        RECT 90.310 135.500 90.450 137.220 ;
        RECT 90.710 136.880 90.970 137.200 ;
        RECT 90.770 135.500 90.910 136.880 ;
        RECT 91.620 136.685 91.900 137.055 ;
        RECT 91.690 135.500 91.830 136.685 ;
        RECT 88.870 135.180 89.130 135.500 ;
        RECT 90.250 135.180 90.510 135.500 ;
        RECT 90.710 135.180 90.970 135.500 ;
        RECT 91.630 135.180 91.890 135.500 ;
        RECT 86.110 134.840 86.370 135.160 ;
        RECT 90.710 133.820 90.970 134.140 ;
        RECT 85.190 133.480 85.450 133.800 ;
        RECT 88.870 133.480 89.130 133.800 ;
        RECT 88.930 131.760 89.070 133.480 ;
        RECT 86.570 131.440 86.830 131.760 ;
        RECT 88.870 131.440 89.130 131.760 ;
        RECT 85.650 130.760 85.910 131.080 ;
        RECT 85.710 129.040 85.850 130.760 ;
        RECT 85.650 128.720 85.910 129.040 ;
        RECT 84.270 128.040 84.530 128.360 ;
        RECT 84.330 127.340 84.470 128.040 ;
        RECT 84.270 127.020 84.530 127.340 ;
        RECT 83.810 126.000 84.070 126.320 ;
        RECT 85.650 126.000 85.910 126.320 ;
        RECT 81.970 125.660 82.230 125.980 ;
        RECT 82.890 125.320 83.150 125.640 ;
        RECT 79.720 124.785 81.260 125.155 ;
        RECT 79.210 123.960 79.470 124.280 ;
        RECT 75.990 123.620 76.250 123.940 ;
        RECT 76.910 123.620 77.170 123.940 ;
        RECT 70.990 123.200 72.970 123.340 ;
        RECT 76.450 123.280 76.710 123.600 ;
        RECT 78.750 123.280 79.010 123.600 ;
        RECT 21.415 122.065 22.955 122.435 ;
        RECT 60.285 122.065 61.825 122.435 ;
        RECT 40.850 119.345 42.390 119.715 ;
        RECT 70.990 118.840 71.130 123.200 ;
        RECT 76.510 121.900 76.650 123.280 ;
        RECT 76.450 121.580 76.710 121.900 ;
        RECT 78.810 120.200 78.950 123.280 ;
        RECT 79.270 121.900 79.410 123.960 ;
        RECT 82.950 123.600 83.090 125.320 ;
        RECT 83.870 125.240 84.010 126.000 ;
        RECT 83.410 125.100 84.010 125.240 ;
        RECT 83.410 123.940 83.550 125.100 ;
        RECT 83.350 123.620 83.610 123.940 ;
        RECT 82.890 123.280 83.150 123.600 ;
        RECT 79.210 121.580 79.470 121.900 ;
        RECT 82.950 120.880 83.090 123.280 ;
        RECT 85.710 121.900 85.850 126.000 ;
        RECT 86.630 124.620 86.770 131.440 ;
        RECT 90.770 130.820 90.910 133.820 ;
        RECT 91.170 132.120 91.430 132.440 ;
        RECT 89.390 130.680 90.910 130.820 ;
        RECT 89.390 129.380 89.530 130.680 ;
        RECT 90.770 130.060 90.910 130.680 ;
        RECT 89.790 129.740 90.050 130.060 ;
        RECT 90.710 129.740 90.970 130.060 ;
        RECT 87.030 129.060 87.290 129.380 ;
        RECT 89.330 129.060 89.590 129.380 ;
        RECT 87.090 126.320 87.230 129.060 ;
        RECT 87.490 128.380 87.750 128.700 ;
        RECT 87.550 127.340 87.690 128.380 ;
        RECT 87.490 127.020 87.750 127.340 ;
        RECT 87.030 126.000 87.290 126.320 ;
        RECT 86.570 124.300 86.830 124.620 ;
        RECT 85.650 121.580 85.910 121.900 ;
        RECT 87.550 121.560 87.690 127.020 ;
        RECT 87.950 125.660 88.210 125.980 ;
        RECT 88.010 124.620 88.150 125.660 ;
        RECT 88.410 125.320 88.670 125.640 ;
        RECT 88.470 124.620 88.610 125.320 ;
        RECT 87.950 124.300 88.210 124.620 ;
        RECT 88.410 124.300 88.670 124.620 ;
        RECT 88.470 123.940 88.610 124.300 ;
        RECT 89.850 123.940 89.990 129.740 ;
        RECT 91.230 124.620 91.370 132.120 ;
        RECT 92.150 125.980 92.290 137.220 ;
        RECT 93.930 133.480 94.190 133.800 ;
        RECT 93.990 131.760 94.130 133.480 ;
        RECT 93.930 131.440 94.190 131.760 ;
        RECT 93.010 127.020 93.270 127.340 ;
        RECT 92.090 125.660 92.350 125.980 ;
        RECT 91.170 124.300 91.430 124.620 ;
        RECT 92.550 124.300 92.810 124.620 ;
        RECT 92.610 123.940 92.750 124.300 ;
        RECT 93.070 123.940 93.210 127.020 ;
        RECT 93.470 125.660 93.730 125.980 ;
        RECT 93.530 125.240 93.670 125.660 ;
        RECT 94.390 125.320 94.650 125.640 ;
        RECT 93.530 125.100 94.130 125.240 ;
        RECT 88.410 123.620 88.670 123.940 ;
        RECT 89.790 123.620 90.050 123.940 ;
        RECT 92.550 123.620 92.810 123.940 ;
        RECT 93.010 123.620 93.270 123.940 ;
        RECT 93.990 123.600 94.130 125.100 ;
        RECT 94.450 124.620 94.590 125.320 ;
        RECT 94.390 124.300 94.650 124.620 ;
        RECT 93.930 123.280 94.190 123.600 ;
        RECT 90.710 122.940 90.970 123.260 ;
        RECT 90.770 121.900 90.910 122.940 ;
        RECT 94.450 121.900 94.590 124.300 ;
        RECT 94.910 123.600 95.050 139.260 ;
        RECT 95.370 130.060 95.510 150.480 ;
        RECT 97.210 146.380 97.350 162.380 ;
        RECT 98.130 159.380 98.270 173.400 ;
        RECT 99.050 173.350 101.090 173.490 ;
        RECT 99.050 171.880 99.190 173.350 ;
        RECT 100.830 173.260 101.090 173.350 ;
        RECT 100.820 172.725 101.100 173.095 ;
        RECT 100.830 172.580 101.090 172.725 ;
        RECT 100.830 171.900 101.090 172.220 ;
        RECT 101.290 171.900 101.550 172.220 ;
        RECT 98.990 171.560 99.250 171.880 ;
        RECT 99.155 171.025 100.695 171.395 ;
        RECT 100.890 170.520 101.030 171.900 ;
        RECT 101.350 170.860 101.490 171.900 ;
        RECT 101.290 170.540 101.550 170.860 ;
        RECT 101.740 170.685 102.020 171.055 ;
        RECT 100.830 170.260 101.090 170.520 ;
        RECT 101.810 170.260 101.950 170.685 ;
        RECT 102.270 170.520 102.410 174.765 ;
        RECT 103.190 173.240 103.330 174.960 ;
        RECT 103.130 172.920 103.390 173.240 ;
        RECT 102.670 172.240 102.930 172.560 ;
        RECT 100.830 170.200 101.950 170.260 ;
        RECT 102.210 170.200 102.470 170.520 ;
        RECT 100.890 170.120 101.950 170.200 ;
        RECT 101.810 169.840 101.950 170.120 ;
        RECT 98.980 169.325 99.260 169.695 ;
        RECT 101.750 169.520 102.010 169.840 ;
        RECT 102.210 169.520 102.470 169.840 ;
        RECT 99.050 167.800 99.190 169.325 ;
        RECT 102.270 168.335 102.410 169.520 ;
        RECT 102.200 167.965 102.480 168.335 ;
        RECT 102.730 168.140 102.870 172.240 ;
        RECT 103.130 171.900 103.390 172.220 ;
        RECT 102.670 167.820 102.930 168.140 ;
        RECT 98.990 167.480 99.250 167.800 ;
        RECT 103.190 167.460 103.330 171.900 ;
        RECT 103.650 170.520 103.790 178.020 ;
        RECT 104.110 176.300 104.250 178.360 ;
        RECT 104.050 175.980 104.310 176.300 ;
        RECT 104.110 175.280 104.250 175.980 ;
        RECT 104.570 175.960 104.710 179.720 ;
        RECT 105.030 177.320 105.170 180.060 ;
        RECT 104.970 177.000 105.230 177.320 ;
        RECT 104.510 175.640 104.770 175.960 ;
        RECT 104.050 174.960 104.310 175.280 ;
        RECT 104.510 174.620 104.770 174.940 ;
        RECT 104.040 172.725 104.320 173.095 ;
        RECT 104.110 170.520 104.250 172.725 ;
        RECT 104.570 172.560 104.710 174.620 ;
        RECT 104.970 173.260 105.230 173.580 ;
        RECT 105.490 173.540 105.630 196.380 ;
        RECT 105.950 191.940 106.090 204.540 ;
        RECT 106.410 204.520 106.550 211.600 ;
        RECT 106.800 210.805 107.080 211.175 ;
        RECT 107.330 210.980 107.470 212.280 ;
        RECT 107.720 212.165 108.000 212.535 ;
        RECT 107.790 211.320 107.930 212.165 ;
        RECT 108.250 211.660 108.390 216.530 ;
        RECT 109.110 216.100 109.370 216.420 ;
        RECT 108.190 211.340 108.450 211.660 ;
        RECT 107.730 211.000 107.990 211.320 ;
        RECT 106.870 210.210 107.010 210.805 ;
        RECT 107.270 210.660 107.530 210.980 ;
        RECT 107.270 210.210 107.530 210.300 ;
        RECT 106.870 210.070 107.530 210.210 ;
        RECT 107.270 209.980 107.530 210.070 ;
        RECT 106.800 209.445 107.080 209.815 ;
        RECT 106.350 204.200 106.610 204.520 ;
        RECT 106.340 203.325 106.620 203.695 ;
        RECT 106.410 203.160 106.550 203.325 ;
        RECT 106.350 202.840 106.610 203.160 ;
        RECT 106.870 199.615 107.010 209.445 ;
        RECT 107.330 209.135 107.470 209.980 ;
        RECT 107.260 208.765 107.540 209.135 ;
        RECT 108.250 208.260 108.390 211.340 ;
        RECT 108.190 207.940 108.450 208.260 ;
        RECT 109.170 207.920 109.310 216.100 ;
        RECT 109.570 215.420 109.830 215.740 ;
        RECT 109.630 214.380 109.770 215.420 ;
        RECT 109.570 214.060 109.830 214.380 ;
        RECT 109.570 210.660 109.830 210.980 ;
        RECT 109.630 209.135 109.770 210.660 ;
        RECT 109.560 208.765 109.840 209.135 ;
        RECT 108.650 207.600 108.910 207.920 ;
        RECT 109.110 207.600 109.370 207.920 ;
        RECT 107.260 206.045 107.540 206.415 ;
        RECT 107.330 205.540 107.470 206.045 ;
        RECT 108.190 205.900 108.450 206.220 ;
        RECT 107.270 205.220 107.530 205.540 ;
        RECT 106.800 199.245 107.080 199.615 ;
        RECT 106.350 198.760 106.610 199.080 ;
        RECT 106.410 197.290 106.550 198.760 ;
        RECT 106.410 197.150 107.010 197.290 ;
        RECT 106.350 196.380 106.610 196.700 ;
        RECT 106.410 195.340 106.550 196.380 ;
        RECT 106.870 196.360 107.010 197.150 ;
        RECT 106.810 196.040 107.070 196.360 ;
        RECT 106.350 195.020 106.610 195.340 ;
        RECT 106.340 193.805 106.620 194.175 ;
        RECT 106.810 194.000 107.070 194.320 ;
        RECT 106.410 193.640 106.550 193.805 ;
        RECT 106.350 193.320 106.610 193.640 ;
        RECT 106.410 191.940 106.550 193.320 ;
        RECT 105.890 191.620 106.150 191.940 ;
        RECT 106.350 191.620 106.610 191.940 ;
        RECT 105.890 190.940 106.150 191.260 ;
        RECT 105.950 190.775 106.090 190.940 ;
        RECT 106.410 190.920 106.550 191.620 ;
        RECT 105.880 190.405 106.160 190.775 ;
        RECT 106.350 190.600 106.610 190.920 ;
        RECT 106.870 189.220 107.010 194.000 ;
        RECT 107.330 189.220 107.470 205.220 ;
        RECT 107.730 204.880 107.990 205.200 ;
        RECT 107.790 200.780 107.930 204.880 ;
        RECT 107.730 200.460 107.990 200.780 ;
        RECT 108.250 200.440 108.390 205.900 ;
        RECT 108.190 200.120 108.450 200.440 ;
        RECT 108.180 199.245 108.460 199.615 ;
        RECT 108.250 196.360 108.390 199.245 ;
        RECT 108.190 196.040 108.450 196.360 ;
        RECT 108.190 195.250 108.450 195.340 ;
        RECT 108.710 195.250 108.850 207.600 ;
        RECT 109.570 201.480 109.830 201.800 ;
        RECT 109.110 199.780 109.370 200.100 ;
        RECT 108.190 195.110 108.850 195.250 ;
        RECT 108.190 195.020 108.450 195.110 ;
        RECT 107.730 194.340 107.990 194.660 ;
        RECT 107.790 193.495 107.930 194.340 ;
        RECT 107.720 193.125 108.000 193.495 ;
        RECT 107.790 191.260 107.930 193.125 ;
        RECT 107.730 190.940 107.990 191.260 ;
        RECT 107.720 190.405 108.000 190.775 ;
        RECT 107.790 189.560 107.930 190.405 ;
        RECT 107.730 189.240 107.990 189.560 ;
        RECT 106.810 188.900 107.070 189.220 ;
        RECT 107.270 188.900 107.530 189.220 ;
        RECT 105.890 185.840 106.150 186.160 ;
        RECT 105.950 182.760 106.090 185.840 ;
        RECT 106.350 185.500 106.610 185.820 ;
        RECT 106.410 184.460 106.550 185.500 ;
        RECT 106.350 184.140 106.610 184.460 ;
        RECT 106.870 183.440 107.010 188.900 ;
        RECT 108.250 186.160 108.390 195.020 ;
        RECT 109.170 192.620 109.310 199.780 ;
        RECT 109.630 194.175 109.770 201.480 ;
        RECT 110.090 197.040 110.230 219.500 ;
        RECT 119.690 218.540 119.950 218.800 ;
        RECT 119.690 218.480 121.270 218.540 ;
        RECT 119.750 218.400 121.270 218.480 ;
        RECT 121.130 218.120 121.270 218.400 ;
        RECT 116.920 217.605 117.200 217.975 ;
        RECT 120.610 217.800 120.870 218.120 ;
        RECT 121.070 217.800 121.330 218.120 ;
        RECT 111.870 216.780 112.130 217.100 ;
        RECT 111.930 216.080 112.070 216.780 ;
        RECT 112.330 216.440 112.590 216.760 ;
        RECT 111.870 215.760 112.130 216.080 ;
        RECT 110.950 213.380 111.210 213.700 ;
        RECT 111.010 210.640 111.150 213.380 ;
        RECT 111.400 212.165 111.680 212.535 ;
        RECT 111.470 211.320 111.610 212.165 ;
        RECT 111.410 211.000 111.670 211.320 ;
        RECT 111.930 210.980 112.070 215.760 ;
        RECT 112.390 212.680 112.530 216.440 ;
        RECT 114.160 216.245 114.440 216.615 ;
        RECT 116.990 216.420 117.130 217.605 ;
        RECT 118.590 217.265 120.130 217.635 ;
        RECT 120.670 217.100 120.810 217.800 ;
        RECT 120.610 216.780 120.870 217.100 ;
        RECT 119.230 216.440 119.490 216.760 ;
        RECT 114.170 216.100 114.430 216.245 ;
        RECT 114.630 216.100 114.890 216.420 ;
        RECT 116.470 216.100 116.730 216.420 ;
        RECT 116.930 216.100 117.190 216.420 ;
        RECT 117.850 216.100 118.110 216.420 ;
        RECT 112.790 214.060 113.050 214.380 ;
        RECT 112.330 212.360 112.590 212.680 ;
        RECT 112.850 211.740 112.990 214.060 ;
        RECT 113.250 212.360 113.510 212.680 ;
        RECT 112.390 211.600 112.990 211.740 ;
        RECT 111.870 210.660 112.130 210.980 ;
        RECT 110.490 210.320 110.750 210.640 ;
        RECT 110.950 210.320 111.210 210.640 ;
        RECT 110.550 208.600 110.690 210.320 ;
        RECT 111.410 208.620 111.670 208.940 ;
        RECT 110.490 208.280 110.750 208.600 ;
        RECT 110.950 207.940 111.210 208.260 ;
        RECT 111.010 207.580 111.150 207.940 ;
        RECT 110.950 207.260 111.210 207.580 ;
        RECT 110.490 204.200 110.750 204.520 ;
        RECT 110.030 196.720 110.290 197.040 ;
        RECT 110.550 194.240 110.690 204.200 ;
        RECT 111.470 199.080 111.610 208.620 ;
        RECT 111.870 206.920 112.130 207.240 ;
        RECT 111.930 206.220 112.070 206.920 ;
        RECT 111.870 205.900 112.130 206.220 ;
        RECT 112.390 205.620 112.530 211.600 ;
        RECT 113.310 208.260 113.450 212.360 ;
        RECT 113.700 210.125 113.980 210.495 ;
        RECT 113.250 207.940 113.510 208.260 ;
        RECT 112.790 207.600 113.050 207.920 ;
        RECT 112.850 206.220 112.990 207.600 ;
        RECT 113.250 207.260 113.510 207.580 ;
        RECT 112.790 205.900 113.050 206.220 ;
        RECT 113.310 205.620 113.450 207.260 ;
        RECT 111.930 205.480 112.530 205.620 ;
        RECT 112.850 205.480 113.450 205.620 ;
        RECT 111.930 203.500 112.070 205.480 ;
        RECT 111.870 203.180 112.130 203.500 ;
        RECT 112.330 202.840 112.590 203.160 ;
        RECT 111.410 198.760 111.670 199.080 ;
        RECT 111.410 197.630 111.670 197.720 ;
        RECT 109.560 193.805 109.840 194.175 ;
        RECT 110.090 194.100 110.690 194.240 ;
        RECT 111.010 197.490 111.670 197.630 ;
        RECT 109.110 192.300 109.370 192.620 ;
        RECT 109.570 192.530 109.830 192.620 ;
        RECT 110.090 192.530 110.230 194.100 ;
        RECT 111.010 193.640 111.150 197.490 ;
        RECT 111.410 197.400 111.670 197.490 ;
        RECT 111.870 197.400 112.130 197.720 ;
        RECT 111.410 196.950 111.670 197.040 ;
        RECT 111.930 196.950 112.070 197.400 ;
        RECT 111.410 196.895 112.070 196.950 ;
        RECT 111.400 196.810 112.070 196.895 ;
        RECT 111.400 196.525 111.680 196.810 ;
        RECT 112.390 196.610 112.530 202.840 ;
        RECT 112.850 196.895 112.990 205.480 ;
        RECT 113.250 204.540 113.510 204.860 ;
        RECT 113.310 201.655 113.450 204.540 ;
        RECT 113.770 202.820 113.910 210.125 ;
        RECT 114.690 207.490 114.830 216.100 ;
        RECT 116.530 214.380 116.670 216.100 ;
        RECT 117.910 214.380 118.050 216.100 ;
        RECT 118.310 215.760 118.570 216.080 ;
        RECT 116.470 214.060 116.730 214.380 ;
        RECT 117.850 214.060 118.110 214.380 ;
        RECT 116.460 213.780 116.740 213.895 ;
        RECT 116.460 213.640 117.590 213.780 ;
        RECT 118.370 213.700 118.510 215.760 ;
        RECT 119.290 215.740 119.430 216.440 ;
        RECT 122.450 216.100 122.710 216.420 ;
        RECT 119.230 215.420 119.490 215.740 ;
        RECT 116.460 213.525 116.740 213.640 ;
        RECT 115.540 212.845 115.820 213.215 ;
        RECT 115.090 210.495 115.350 210.640 ;
        RECT 115.080 210.125 115.360 210.495 ;
        RECT 115.610 208.260 115.750 212.845 ;
        RECT 116.930 212.700 117.190 213.020 ;
        RECT 116.470 211.340 116.730 211.660 ;
        RECT 115.550 207.940 115.810 208.260 ;
        RECT 116.010 207.600 116.270 207.920 ;
        RECT 115.550 207.490 115.810 207.580 ;
        RECT 114.690 207.350 115.810 207.490 ;
        RECT 114.170 206.920 114.430 207.240 ;
        RECT 113.710 202.500 113.970 202.820 ;
        RECT 114.230 202.480 114.370 206.920 ;
        RECT 114.690 206.220 114.830 207.350 ;
        RECT 115.550 207.260 115.810 207.350 ;
        RECT 116.070 207.095 116.210 207.600 ;
        RECT 116.530 207.240 116.670 211.340 ;
        RECT 116.990 210.980 117.130 212.700 ;
        RECT 117.450 210.980 117.590 213.640 ;
        RECT 117.850 213.380 118.110 213.700 ;
        RECT 118.310 213.380 118.570 213.700 ;
        RECT 118.760 213.525 119.040 213.895 ;
        RECT 116.930 210.660 117.190 210.980 ;
        RECT 117.390 210.660 117.650 210.980 ;
        RECT 117.450 209.135 117.590 210.660 ;
        RECT 117.910 209.960 118.050 213.380 ;
        RECT 118.830 213.020 118.970 213.525 ;
        RECT 121.530 213.040 121.790 213.360 ;
        RECT 118.770 212.700 119.030 213.020 ;
        RECT 118.590 211.825 120.130 212.195 ;
        RECT 121.590 210.980 121.730 213.040 ;
        RECT 121.990 211.000 122.250 211.320 ;
        RECT 119.690 210.660 119.950 210.980 ;
        RECT 121.530 210.660 121.790 210.980 ;
        RECT 117.850 209.640 118.110 209.960 ;
        RECT 118.770 209.640 119.030 209.960 ;
        RECT 116.930 208.620 117.190 208.940 ;
        RECT 117.380 208.765 117.660 209.135 ;
        RECT 116.000 206.725 116.280 207.095 ;
        RECT 116.470 206.920 116.730 207.240 ;
        RECT 114.630 205.900 114.890 206.220 ;
        RECT 115.090 205.900 115.350 206.220 ;
        RECT 114.630 204.880 114.890 205.200 ;
        RECT 114.690 203.015 114.830 204.880 ;
        RECT 115.150 203.160 115.290 205.900 ;
        RECT 116.070 205.540 116.210 206.725 ;
        RECT 116.010 205.220 116.270 205.540 ;
        RECT 114.620 202.645 114.900 203.015 ;
        RECT 115.090 202.840 115.350 203.160 ;
        RECT 114.170 202.160 114.430 202.480 ;
        RECT 113.240 201.285 113.520 201.655 ;
        RECT 111.930 196.470 112.530 196.610 ;
        RECT 112.780 196.525 113.060 196.895 ;
        RECT 111.400 195.165 111.680 195.535 ;
        RECT 111.470 195.000 111.610 195.165 ;
        RECT 111.410 194.680 111.670 195.000 ;
        RECT 110.950 193.320 111.210 193.640 ;
        RECT 109.570 192.390 110.230 192.530 ;
        RECT 109.570 192.300 109.830 192.390 ;
        RECT 109.630 191.600 109.770 192.300 ;
        RECT 109.570 191.280 109.830 191.600 ;
        RECT 108.650 186.180 108.910 186.500 ;
        RECT 108.190 185.840 108.450 186.160 ;
        RECT 108.710 183.440 108.850 186.180 ;
        RECT 109.630 184.460 109.770 191.280 ;
        RECT 111.010 189.220 111.150 193.320 ;
        RECT 110.950 188.900 111.210 189.220 ;
        RECT 110.020 186.325 110.300 186.695 ;
        RECT 111.010 186.500 111.150 188.900 ;
        RECT 109.570 184.140 109.830 184.460 ;
        RECT 106.810 183.120 107.070 183.440 ;
        RECT 107.730 183.120 107.990 183.440 ;
        RECT 108.650 183.120 108.910 183.440 ;
        RECT 105.890 182.440 106.150 182.760 ;
        RECT 107.790 181.400 107.930 183.120 ;
        RECT 108.710 181.740 108.850 183.120 ;
        RECT 109.100 182.925 109.380 183.295 ;
        RECT 108.650 181.420 108.910 181.740 ;
        RECT 107.730 181.080 107.990 181.400 ;
        RECT 108.190 180.400 108.450 180.720 ;
        RECT 107.730 180.060 107.990 180.380 ;
        RECT 105.890 178.700 106.150 179.020 ;
        RECT 105.950 178.340 106.090 178.700 ;
        RECT 107.790 178.340 107.930 180.060 ;
        RECT 108.250 179.020 108.390 180.400 ;
        RECT 109.170 179.020 109.310 182.925 ;
        RECT 108.190 178.700 108.450 179.020 ;
        RECT 109.110 178.700 109.370 179.020 ;
        RECT 105.890 178.020 106.150 178.340 ;
        RECT 107.730 178.020 107.990 178.340 ;
        RECT 107.270 177.000 107.530 177.320 ;
        RECT 107.730 177.000 107.990 177.320 ;
        RECT 106.350 175.980 106.610 176.300 ;
        RECT 106.410 175.280 106.550 175.980 ;
        RECT 106.350 175.190 106.610 175.280 ;
        RECT 106.350 175.050 107.010 175.190 ;
        RECT 106.350 174.960 106.610 175.050 ;
        RECT 105.490 173.400 106.550 173.540 ;
        RECT 104.510 172.240 104.770 172.560 ;
        RECT 103.590 170.200 103.850 170.520 ;
        RECT 104.050 170.200 104.310 170.520 ;
        RECT 105.030 169.840 105.170 173.260 ;
        RECT 105.430 172.810 105.690 172.900 ;
        RECT 105.430 172.670 106.090 172.810 ;
        RECT 105.430 172.580 105.690 172.670 ;
        RECT 105.430 171.900 105.690 172.220 ;
        RECT 105.490 169.840 105.630 171.900 ;
        RECT 104.970 169.520 105.230 169.840 ;
        RECT 105.430 169.520 105.690 169.840 ;
        RECT 104.510 168.840 104.770 169.160 ;
        RECT 104.050 167.820 104.310 168.140 ;
        RECT 101.750 167.140 102.010 167.460 ;
        RECT 103.130 167.140 103.390 167.460 ;
        RECT 98.530 166.975 98.790 167.120 ;
        RECT 98.520 166.605 98.800 166.975 ;
        RECT 98.590 162.700 98.730 166.605 ;
        RECT 99.155 165.585 100.695 165.955 ;
        RECT 101.810 165.420 101.950 167.140 ;
        RECT 102.670 166.800 102.930 167.120 ;
        RECT 102.210 166.120 102.470 166.440 ;
        RECT 101.750 165.100 102.010 165.420 ;
        RECT 102.270 164.255 102.410 166.120 ;
        RECT 100.830 163.740 101.090 164.060 ;
        RECT 102.200 163.885 102.480 164.255 ;
        RECT 98.530 162.380 98.790 162.700 ;
        RECT 99.155 160.145 100.695 160.515 ;
        RECT 97.670 159.240 98.270 159.380 ;
        RECT 97.670 152.840 97.810 159.240 ;
        RECT 98.070 158.300 98.330 158.620 ;
        RECT 99.910 158.300 100.170 158.620 ;
        RECT 97.610 152.520 97.870 152.840 ;
        RECT 98.130 149.100 98.270 158.300 ;
        RECT 99.970 157.260 100.110 158.300 ;
        RECT 99.910 156.940 100.170 157.260 ;
        RECT 98.530 155.920 98.790 156.240 ;
        RECT 98.590 153.940 98.730 155.920 ;
        RECT 99.155 154.705 100.695 155.075 ;
        RECT 98.980 153.940 99.260 154.055 ;
        RECT 98.590 153.800 99.260 153.940 ;
        RECT 98.980 153.685 99.260 153.800 ;
        RECT 98.990 153.540 99.250 153.685 ;
        RECT 98.530 151.160 98.790 151.480 ;
        RECT 98.070 148.780 98.330 149.100 ;
        RECT 97.150 146.060 97.410 146.380 ;
        RECT 96.690 144.360 96.950 144.680 ;
        RECT 96.230 141.980 96.490 142.300 ;
        RECT 96.290 141.815 96.430 141.980 ;
        RECT 96.220 141.445 96.500 141.815 ;
        RECT 96.750 140.455 96.890 144.360 ;
        RECT 98.590 143.320 98.730 151.160 ;
        RECT 100.890 150.460 101.030 163.740 ;
        RECT 102.730 162.360 102.870 166.800 ;
        RECT 103.590 166.350 103.850 166.440 ;
        RECT 104.110 166.350 104.250 167.820 ;
        RECT 104.570 167.800 104.710 168.840 ;
        RECT 104.510 167.480 104.770 167.800 ;
        RECT 103.590 166.210 104.250 166.350 ;
        RECT 103.590 166.120 103.850 166.210 ;
        RECT 103.130 163.400 103.390 163.720 ;
        RECT 104.510 163.400 104.770 163.720 ;
        RECT 102.670 162.040 102.930 162.360 ;
        RECT 102.730 161.680 102.870 162.040 ;
        RECT 102.670 161.360 102.930 161.680 ;
        RECT 103.190 159.890 103.330 163.400 ;
        RECT 104.570 161.535 104.710 163.400 ;
        RECT 104.970 162.040 105.230 162.360 ;
        RECT 104.500 161.165 104.780 161.535 ;
        RECT 103.190 159.750 103.790 159.890 ;
        RECT 103.120 159.125 103.400 159.495 ;
        RECT 103.190 158.280 103.330 159.125 ;
        RECT 103.650 158.530 103.790 159.750 ;
        RECT 105.030 159.640 105.170 162.040 ;
        RECT 105.950 160.855 106.090 172.670 ;
        RECT 105.880 160.740 106.160 160.855 ;
        RECT 105.490 160.600 106.160 160.740 ;
        RECT 104.970 159.320 105.230 159.640 ;
        RECT 104.970 158.530 105.230 158.620 ;
        RECT 103.650 158.390 105.230 158.530 ;
        RECT 104.970 158.300 105.230 158.390 ;
        RECT 102.670 157.960 102.930 158.280 ;
        RECT 103.130 157.960 103.390 158.280 ;
        RECT 101.290 156.940 101.550 157.260 ;
        RECT 101.350 153.180 101.490 156.940 ;
        RECT 102.730 156.775 102.870 157.960 ;
        RECT 102.660 156.405 102.940 156.775 ;
        RECT 101.750 154.220 102.010 154.540 ;
        RECT 101.290 152.860 101.550 153.180 ;
        RECT 100.830 150.140 101.090 150.460 ;
        RECT 101.280 150.285 101.560 150.655 ;
        RECT 99.155 149.265 100.695 149.635 ;
        RECT 100.370 147.990 100.630 148.080 ;
        RECT 100.890 147.990 101.030 150.140 ;
        RECT 100.370 147.850 101.030 147.990 ;
        RECT 100.370 147.760 100.630 147.850 ;
        RECT 100.820 146.885 101.100 147.255 ;
        RECT 100.890 145.700 101.030 146.885 ;
        RECT 101.350 146.380 101.490 150.285 ;
        RECT 101.290 146.060 101.550 146.380 ;
        RECT 101.350 145.700 101.490 146.060 ;
        RECT 98.990 145.380 99.250 145.700 ;
        RECT 100.830 145.380 101.090 145.700 ;
        RECT 101.290 145.380 101.550 145.700 ;
        RECT 99.050 144.680 99.190 145.380 ;
        RECT 98.990 144.360 99.250 144.680 ;
        RECT 100.830 144.360 101.090 144.680 ;
        RECT 99.155 143.825 100.695 144.195 ;
        RECT 98.530 143.000 98.790 143.320 ;
        RECT 98.990 142.320 99.250 142.640 ;
        RECT 99.910 142.320 100.170 142.640 ;
        RECT 98.070 141.640 98.330 141.960 ;
        RECT 96.680 140.085 96.960 140.455 ;
        RECT 97.610 139.940 97.870 140.260 ;
        RECT 97.150 138.920 97.410 139.240 ;
        RECT 97.210 137.540 97.350 138.920 ;
        RECT 97.150 137.220 97.410 137.540 ;
        RECT 96.690 136.540 96.950 136.860 ;
        RECT 96.230 136.200 96.490 136.520 ;
        RECT 96.290 134.820 96.430 136.200 ;
        RECT 96.750 134.820 96.890 136.540 ;
        RECT 96.230 134.500 96.490 134.820 ;
        RECT 96.690 134.500 96.950 134.820 ;
        RECT 97.670 134.390 97.810 139.940 ;
        RECT 98.130 138.220 98.270 141.640 ;
        RECT 99.050 140.940 99.190 142.320 ;
        RECT 98.990 140.620 99.250 140.940 ;
        RECT 99.970 140.600 100.110 142.320 ;
        RECT 100.370 141.980 100.630 142.300 ;
        RECT 99.910 140.280 100.170 140.600 ;
        RECT 100.430 140.260 100.570 141.980 ;
        RECT 100.370 139.940 100.630 140.260 ;
        RECT 98.530 139.600 98.790 139.920 ;
        RECT 98.070 137.900 98.330 138.220 ;
        RECT 98.590 137.880 98.730 139.600 ;
        RECT 99.155 138.385 100.695 138.755 ;
        RECT 98.530 137.560 98.790 137.880 ;
        RECT 98.530 136.880 98.790 137.200 ;
        RECT 98.070 134.390 98.330 134.480 ;
        RECT 97.670 134.250 98.330 134.390 ;
        RECT 98.070 134.160 98.330 134.250 ;
        RECT 95.770 133.820 96.030 134.140 ;
        RECT 95.830 131.760 95.970 133.820 ;
        RECT 97.150 133.480 97.410 133.800 ;
        RECT 97.210 131.760 97.350 133.480 ;
        RECT 98.130 132.100 98.270 134.160 ;
        RECT 98.590 132.780 98.730 136.880 ;
        RECT 99.155 132.945 100.695 133.315 ;
        RECT 98.530 132.460 98.790 132.780 ;
        RECT 98.070 131.780 98.330 132.100 ;
        RECT 98.590 131.760 98.730 132.460 ;
        RECT 95.770 131.440 96.030 131.760 ;
        RECT 97.150 131.440 97.410 131.760 ;
        RECT 98.530 131.440 98.790 131.760 ;
        RECT 100.370 131.440 100.630 131.760 ;
        RECT 97.150 130.760 97.410 131.080 ;
        RECT 98.530 130.760 98.790 131.080 ;
        RECT 95.310 129.740 95.570 130.060 ;
        RECT 95.370 129.380 95.510 129.740 ;
        RECT 95.310 129.060 95.570 129.380 ;
        RECT 95.310 125.320 95.570 125.640 ;
        RECT 96.690 125.320 96.950 125.640 ;
        RECT 95.370 123.940 95.510 125.320 ;
        RECT 96.750 123.940 96.890 125.320 ;
        RECT 97.210 123.940 97.350 130.760 ;
        RECT 98.070 128.380 98.330 128.700 ;
        RECT 98.130 126.660 98.270 128.380 ;
        RECT 98.590 126.660 98.730 130.760 ;
        RECT 100.430 128.700 100.570 131.440 ;
        RECT 100.890 129.380 101.030 144.360 ;
        RECT 101.290 142.660 101.550 142.980 ;
        RECT 101.810 142.890 101.950 154.220 ;
        RECT 102.210 153.540 102.470 153.860 ;
        RECT 102.270 151.900 102.410 153.540 ;
        RECT 102.660 151.900 102.940 152.015 ;
        RECT 102.270 151.760 102.940 151.900 ;
        RECT 102.270 151.480 102.410 151.760 ;
        RECT 102.660 151.645 102.940 151.760 ;
        RECT 102.210 151.160 102.470 151.480 ;
        RECT 102.670 151.160 102.930 151.480 ;
        RECT 102.270 147.255 102.410 151.160 ;
        RECT 102.200 146.885 102.480 147.255 ;
        RECT 102.730 146.575 102.870 151.160 ;
        RECT 103.190 150.800 103.330 157.960 ;
        RECT 105.490 157.340 105.630 160.600 ;
        RECT 105.880 160.485 106.160 160.600 ;
        RECT 105.890 159.660 106.150 159.980 ;
        RECT 103.650 157.200 105.630 157.340 ;
        RECT 103.650 155.560 103.790 157.200 ;
        RECT 105.950 156.920 106.090 159.660 ;
        RECT 105.890 156.600 106.150 156.920 ;
        RECT 103.590 155.240 103.850 155.560 ;
        RECT 105.890 150.820 106.150 151.140 ;
        RECT 103.130 150.480 103.390 150.800 ;
        RECT 104.970 150.480 105.230 150.800 ;
        RECT 103.590 149.975 103.850 150.120 ;
        RECT 103.580 149.605 103.860 149.975 ;
        RECT 104.050 149.800 104.310 150.120 ;
        RECT 104.110 148.760 104.250 149.800 ;
        RECT 104.050 148.440 104.310 148.760 ;
        RECT 102.660 146.205 102.940 146.575 ;
        RECT 102.670 145.380 102.930 145.700 ;
        RECT 102.210 144.930 102.470 145.020 ;
        RECT 102.730 144.930 102.870 145.380 ;
        RECT 102.210 144.790 102.870 144.930 ;
        RECT 102.210 144.700 102.470 144.790 ;
        RECT 101.810 142.750 102.410 142.890 ;
        RECT 101.350 140.260 101.490 142.660 ;
        RECT 101.290 139.940 101.550 140.260 ;
        RECT 101.290 138.920 101.550 139.240 ;
        RECT 101.350 136.860 101.490 138.920 ;
        RECT 101.290 136.540 101.550 136.860 ;
        RECT 102.270 136.520 102.410 142.750 ;
        RECT 102.670 141.980 102.930 142.300 ;
        RECT 102.730 140.600 102.870 141.980 ;
        RECT 102.670 140.280 102.930 140.600 ;
        RECT 103.130 140.170 103.390 140.260 ;
        RECT 103.130 140.030 104.250 140.170 ;
        RECT 103.130 139.940 103.390 140.030 ;
        RECT 102.670 138.920 102.930 139.240 ;
        RECT 102.730 136.520 102.870 138.920 ;
        RECT 102.210 136.200 102.470 136.520 ;
        RECT 102.670 136.200 102.930 136.520 ;
        RECT 102.270 134.820 102.410 136.200 ;
        RECT 102.210 134.500 102.470 134.820 ;
        RECT 102.730 132.440 102.870 136.200 ;
        RECT 104.110 134.820 104.250 140.030 ;
        RECT 104.510 139.940 104.770 140.260 ;
        RECT 104.570 134.820 104.710 139.940 ;
        RECT 104.050 134.500 104.310 134.820 ;
        RECT 104.510 134.500 104.770 134.820 ;
        RECT 102.200 132.180 102.480 132.295 ;
        RECT 101.350 132.040 102.480 132.180 ;
        RECT 102.670 132.120 102.930 132.440 ;
        RECT 101.350 131.760 101.490 132.040 ;
        RECT 102.200 131.925 102.480 132.040 ;
        RECT 101.290 131.440 101.550 131.760 ;
        RECT 101.750 131.440 102.010 131.760 ;
        RECT 102.210 131.440 102.470 131.760 ;
        RECT 101.290 130.760 101.550 131.080 ;
        RECT 101.350 130.060 101.490 130.760 ;
        RECT 101.810 130.060 101.950 131.440 ;
        RECT 101.290 129.740 101.550 130.060 ;
        RECT 101.750 129.740 102.010 130.060 ;
        RECT 100.830 129.060 101.090 129.380 ;
        RECT 101.290 129.060 101.550 129.380 ;
        RECT 100.370 128.380 100.630 128.700 ;
        RECT 99.155 127.505 100.695 127.875 ;
        RECT 101.350 126.740 101.490 129.060 ;
        RECT 102.270 127.340 102.410 131.440 ;
        RECT 104.570 129.460 104.710 134.500 ;
        RECT 105.030 130.060 105.170 150.480 ;
        RECT 105.950 145.020 106.090 150.820 ;
        RECT 106.410 148.080 106.550 173.400 ;
        RECT 106.870 170.860 107.010 175.050 ;
        RECT 107.330 170.860 107.470 177.000 ;
        RECT 107.790 174.600 107.930 177.000 ;
        RECT 108.250 174.600 108.390 178.700 ;
        RECT 109.630 177.320 109.770 184.140 ;
        RECT 110.090 183.350 110.230 186.325 ;
        RECT 110.950 186.180 111.210 186.500 ;
        RECT 110.490 183.350 110.750 183.440 ;
        RECT 110.090 183.210 110.750 183.350 ;
        RECT 110.090 181.935 110.230 183.210 ;
        RECT 110.490 183.120 110.750 183.210 ;
        RECT 110.020 181.565 110.300 181.935 ;
        RECT 110.020 180.885 110.300 181.255 ;
        RECT 110.030 180.740 110.290 180.885 ;
        RECT 111.010 179.020 111.150 186.180 ;
        RECT 111.470 180.575 111.610 194.680 ;
        RECT 111.930 186.160 112.070 196.470 ;
        RECT 112.790 194.340 113.050 194.660 ;
        RECT 112.850 189.900 112.990 194.340 ;
        RECT 112.790 189.580 113.050 189.900 ;
        RECT 113.310 189.300 113.450 201.285 ;
        RECT 114.690 199.420 114.830 202.645 ;
        RECT 115.550 202.500 115.810 202.820 ;
        RECT 115.090 202.160 115.350 202.480 ;
        RECT 114.630 199.100 114.890 199.420 ;
        RECT 114.690 197.040 114.830 199.100 ;
        RECT 114.630 196.720 114.890 197.040 ;
        RECT 113.710 194.680 113.970 195.000 ;
        RECT 113.770 193.640 113.910 194.680 ;
        RECT 114.630 193.660 114.890 193.980 ;
        RECT 113.710 193.320 113.970 193.640 ;
        RECT 114.170 193.320 114.430 193.640 ;
        RECT 114.230 191.940 114.370 193.320 ;
        RECT 114.170 191.620 114.430 191.940 ;
        RECT 114.690 191.600 114.830 193.660 ;
        RECT 115.150 192.620 115.290 202.160 ;
        RECT 115.610 196.780 115.750 202.500 ;
        RECT 116.070 200.440 116.210 205.220 ;
        RECT 116.470 200.460 116.730 200.780 ;
        RECT 116.010 200.120 116.270 200.440 ;
        RECT 116.530 199.615 116.670 200.460 ;
        RECT 116.460 199.245 116.740 199.615 ;
        RECT 115.610 196.640 116.210 196.780 ;
        RECT 115.550 196.040 115.810 196.360 ;
        RECT 115.610 194.660 115.750 196.040 ;
        RECT 115.550 194.340 115.810 194.660 ;
        RECT 115.090 192.300 115.350 192.620 ;
        RECT 115.550 192.300 115.810 192.620 ;
        RECT 114.630 191.280 114.890 191.600 ;
        RECT 115.090 189.470 115.350 189.560 ;
        RECT 112.390 189.160 113.450 189.300 ;
        RECT 114.690 189.330 115.350 189.470 ;
        RECT 111.870 185.840 112.130 186.160 ;
        RECT 111.930 184.460 112.070 185.840 ;
        RECT 111.870 184.140 112.130 184.460 ;
        RECT 112.390 183.100 112.530 189.160 ;
        RECT 113.710 188.900 113.970 189.220 ;
        RECT 112.790 187.880 113.050 188.200 ;
        RECT 113.770 187.940 113.910 188.900 ;
        RECT 114.160 188.365 114.440 188.735 ;
        RECT 112.850 187.180 112.990 187.880 ;
        RECT 113.310 187.800 113.910 187.940 ;
        RECT 112.790 186.860 113.050 187.180 ;
        RECT 113.310 183.860 113.450 187.800 ;
        RECT 114.230 187.180 114.370 188.365 ;
        RECT 113.710 186.860 113.970 187.180 ;
        RECT 114.170 186.860 114.430 187.180 ;
        RECT 113.770 186.580 113.910 186.860 ;
        RECT 114.160 186.580 114.440 186.695 ;
        RECT 113.770 186.440 114.440 186.580 ;
        RECT 114.160 186.325 114.440 186.440 ;
        RECT 114.170 185.840 114.430 186.160 ;
        RECT 113.710 185.500 113.970 185.820 ;
        RECT 113.770 183.975 113.910 185.500 ;
        RECT 112.850 183.720 113.450 183.860 ;
        RECT 112.330 182.780 112.590 183.100 ;
        RECT 111.400 180.205 111.680 180.575 ;
        RECT 110.950 178.700 111.210 179.020 ;
        RECT 112.850 178.535 112.990 183.720 ;
        RECT 113.700 183.605 113.980 183.975 ;
        RECT 114.230 182.760 114.370 185.840 ;
        RECT 114.690 185.820 114.830 189.330 ;
        RECT 115.090 189.240 115.350 189.330 ;
        RECT 115.090 186.860 115.350 187.180 ;
        RECT 115.150 186.160 115.290 186.860 ;
        RECT 115.090 185.840 115.350 186.160 ;
        RECT 114.630 185.500 114.890 185.820 ;
        RECT 114.630 183.460 114.890 183.780 ;
        RECT 114.170 182.440 114.430 182.760 ;
        RECT 113.710 181.420 113.970 181.740 ;
        RECT 113.250 180.400 113.510 180.720 ;
        RECT 113.310 178.680 113.450 180.400 ;
        RECT 113.770 180.380 113.910 181.420 ;
        RECT 114.690 180.720 114.830 183.460 ;
        RECT 115.090 183.120 115.350 183.440 ;
        RECT 114.630 180.400 114.890 180.720 ;
        RECT 113.710 180.060 113.970 180.380 ;
        RECT 110.490 178.020 110.750 178.340 ;
        RECT 112.780 178.165 113.060 178.535 ;
        RECT 113.250 178.360 113.510 178.680 ;
        RECT 113.770 178.340 113.910 180.060 ;
        RECT 113.710 178.020 113.970 178.340 ;
        RECT 109.570 177.000 109.830 177.320 ;
        RECT 110.020 176.805 110.300 177.175 ;
        RECT 110.090 175.620 110.230 176.805 ;
        RECT 110.550 176.300 110.690 178.020 ;
        RECT 113.770 176.300 113.910 178.020 ;
        RECT 110.490 175.980 110.750 176.300 ;
        RECT 113.710 175.980 113.970 176.300 ;
        RECT 110.030 175.300 110.290 175.620 ;
        RECT 111.410 174.960 111.670 175.280 ;
        RECT 112.330 174.960 112.590 175.280 ;
        RECT 113.770 175.135 113.910 175.980 ;
        RECT 114.630 175.530 114.890 175.620 ;
        RECT 115.150 175.530 115.290 183.120 ;
        RECT 114.630 175.390 115.290 175.530 ;
        RECT 114.630 175.300 114.890 175.390 ;
        RECT 107.730 174.280 107.990 174.600 ;
        RECT 108.190 174.280 108.450 174.600 ;
        RECT 111.470 173.580 111.610 174.960 ;
        RECT 109.570 173.260 109.830 173.580 ;
        RECT 111.410 173.260 111.670 173.580 ;
        RECT 108.640 172.725 108.920 173.095 ;
        RECT 109.630 172.900 109.770 173.260 ;
        RECT 110.950 172.920 111.210 173.240 ;
        RECT 108.710 172.560 108.850 172.725 ;
        RECT 109.570 172.580 109.830 172.900 ;
        RECT 108.650 172.240 108.910 172.560 ;
        RECT 108.650 171.735 108.910 171.880 ;
        RECT 108.640 171.365 108.920 171.735 ;
        RECT 110.490 171.560 110.750 171.880 ;
        RECT 106.810 170.540 107.070 170.860 ;
        RECT 107.270 170.540 107.530 170.860 ;
        RECT 107.270 169.520 107.530 169.840 ;
        RECT 106.800 168.645 107.080 169.015 ;
        RECT 106.870 167.800 107.010 168.645 ;
        RECT 107.330 168.140 107.470 169.520 ;
        RECT 107.270 167.820 107.530 168.140 ;
        RECT 106.810 167.480 107.070 167.800 ;
        RECT 109.560 167.285 109.840 167.655 ;
        RECT 109.570 167.140 109.830 167.285 ;
        RECT 108.650 166.460 108.910 166.780 ;
        RECT 107.270 165.100 107.530 165.420 ;
        RECT 107.330 164.310 107.470 165.100 ;
        RECT 108.190 164.310 108.450 164.400 ;
        RECT 107.330 164.170 108.450 164.310 ;
        RECT 108.190 164.080 108.450 164.170 ;
        RECT 108.250 162.700 108.390 164.080 ;
        RECT 108.190 162.380 108.450 162.700 ;
        RECT 108.190 161.360 108.450 161.680 ;
        RECT 106.800 159.125 107.080 159.495 ;
        RECT 106.870 157.260 107.010 159.125 ;
        RECT 106.810 156.940 107.070 157.260 ;
        RECT 106.870 154.540 107.010 156.940 ;
        RECT 106.810 154.220 107.070 154.540 ;
        RECT 107.730 148.100 107.990 148.420 ;
        RECT 106.350 147.760 106.610 148.080 ;
        RECT 105.890 144.700 106.150 145.020 ;
        RECT 105.890 143.340 106.150 143.660 ;
        RECT 105.430 142.320 105.690 142.640 ;
        RECT 105.490 139.920 105.630 142.320 ;
        RECT 105.950 140.940 106.090 143.340 ;
        RECT 106.350 143.000 106.610 143.320 ;
        RECT 106.810 143.000 107.070 143.320 ;
        RECT 105.890 140.620 106.150 140.940 ;
        RECT 105.430 139.600 105.690 139.920 ;
        RECT 105.490 137.880 105.630 139.600 ;
        RECT 105.430 137.560 105.690 137.880 ;
        RECT 105.950 135.160 106.090 140.620 ;
        RECT 105.890 134.840 106.150 135.160 ;
        RECT 105.950 131.760 106.090 134.840 ;
        RECT 106.410 131.760 106.550 143.000 ;
        RECT 106.870 137.735 107.010 143.000 ;
        RECT 106.800 137.365 107.080 137.735 ;
        RECT 106.810 133.820 107.070 134.140 ;
        RECT 105.890 131.440 106.150 131.760 ;
        RECT 106.350 131.615 106.610 131.760 ;
        RECT 106.340 131.245 106.620 131.615 ;
        RECT 104.970 129.740 105.230 130.060 ;
        RECT 103.650 129.320 104.710 129.460 ;
        RECT 102.670 128.040 102.930 128.360 ;
        RECT 102.730 127.340 102.870 128.040 ;
        RECT 102.210 127.020 102.470 127.340 ;
        RECT 102.670 127.020 102.930 127.340 ;
        RECT 103.650 127.000 103.790 129.320 ;
        RECT 104.960 129.205 105.240 129.575 ;
        RECT 106.870 129.290 107.010 133.820 ;
        RECT 107.790 131.500 107.930 148.100 ;
        RECT 108.250 147.740 108.390 161.360 ;
        RECT 108.710 159.980 108.850 166.460 ;
        RECT 108.650 159.660 108.910 159.980 ;
        RECT 109.110 159.320 109.370 159.640 ;
        RECT 108.650 157.960 108.910 158.280 ;
        RECT 108.710 157.260 108.850 157.960 ;
        RECT 108.650 156.940 108.910 157.260 ;
        RECT 109.170 156.240 109.310 159.320 ;
        RECT 109.630 158.960 109.770 167.140 ;
        RECT 110.550 167.120 110.690 171.560 ;
        RECT 111.010 170.180 111.150 172.920 ;
        RECT 111.410 171.560 111.670 171.880 ;
        RECT 111.470 170.520 111.610 171.560 ;
        RECT 111.410 170.200 111.670 170.520 ;
        RECT 110.950 169.860 111.210 170.180 ;
        RECT 110.490 166.800 110.750 167.120 ;
        RECT 111.010 166.440 111.150 169.860 ;
        RECT 111.470 169.840 111.610 170.200 ;
        RECT 111.410 169.520 111.670 169.840 ;
        RECT 110.950 166.120 111.210 166.440 ;
        RECT 112.390 161.680 112.530 174.960 ;
        RECT 113.700 174.765 113.980 175.135 ;
        RECT 115.610 174.340 115.750 192.300 ;
        RECT 116.070 189.900 116.210 196.640 ;
        RECT 116.530 194.660 116.670 199.245 ;
        RECT 116.470 194.340 116.730 194.660 ;
        RECT 116.990 192.620 117.130 208.620 ;
        RECT 117.910 207.490 118.050 209.640 ;
        RECT 118.830 208.040 118.970 209.640 ;
        RECT 119.750 208.260 119.890 210.660 ;
        RECT 118.370 207.920 118.970 208.040 ;
        RECT 119.690 207.940 119.950 208.260 ;
        RECT 121.070 207.940 121.330 208.260 ;
        RECT 118.310 207.900 118.970 207.920 ;
        RECT 118.310 207.600 118.570 207.900 ;
        RECT 119.230 207.600 119.490 207.920 ;
        RECT 117.450 207.350 118.050 207.490 ;
        RECT 117.450 204.520 117.590 207.350 ;
        RECT 119.290 207.150 119.430 207.600 ;
        RECT 117.910 207.010 119.430 207.150 ;
        RECT 117.390 204.200 117.650 204.520 ;
        RECT 117.390 202.160 117.650 202.480 ;
        RECT 117.450 200.780 117.590 202.160 ;
        RECT 117.910 200.975 118.050 207.010 ;
        RECT 120.610 206.920 120.870 207.240 ;
        RECT 118.590 206.385 120.130 206.755 ;
        RECT 118.770 205.560 119.030 205.880 ;
        RECT 118.830 202.480 118.970 205.560 ;
        RECT 120.670 205.200 120.810 206.920 ;
        RECT 120.610 204.880 120.870 205.200 ;
        RECT 120.150 204.200 120.410 204.520 ;
        RECT 120.210 202.480 120.350 204.200 ;
        RECT 120.610 203.180 120.870 203.500 ;
        RECT 118.770 202.160 119.030 202.480 ;
        RECT 120.150 202.160 120.410 202.480 ;
        RECT 117.390 200.460 117.650 200.780 ;
        RECT 117.840 200.605 118.120 200.975 ;
        RECT 118.590 200.945 120.130 201.315 ;
        RECT 117.910 200.440 118.050 200.605 ;
        RECT 117.850 200.120 118.110 200.440 ;
        RECT 119.690 198.760 119.950 199.080 ;
        RECT 117.390 197.400 117.650 197.720 ;
        RECT 118.770 197.400 119.030 197.720 ;
        RECT 116.930 192.300 117.190 192.620 ;
        RECT 116.470 190.600 116.730 190.920 ;
        RECT 116.010 189.580 116.270 189.900 ;
        RECT 116.010 188.900 116.270 189.220 ;
        RECT 116.070 182.760 116.210 188.900 ;
        RECT 116.530 186.160 116.670 190.600 ;
        RECT 116.920 189.725 117.200 190.095 ;
        RECT 116.930 189.580 117.190 189.725 ;
        RECT 116.920 189.045 117.200 189.415 ;
        RECT 116.470 185.840 116.730 186.160 ;
        RECT 116.460 183.605 116.740 183.975 ;
        RECT 116.990 183.780 117.130 189.045 ;
        RECT 117.450 188.880 117.590 197.400 ;
        RECT 117.850 197.060 118.110 197.380 ;
        RECT 117.910 193.980 118.050 197.060 ;
        RECT 118.830 196.700 118.970 197.400 ;
        RECT 119.750 197.380 119.890 198.760 ;
        RECT 120.670 198.060 120.810 203.180 ;
        RECT 121.130 198.935 121.270 207.940 ;
        RECT 121.590 202.820 121.730 210.660 ;
        RECT 121.530 202.500 121.790 202.820 ;
        RECT 121.590 200.975 121.730 202.500 ;
        RECT 121.520 200.605 121.800 200.975 ;
        RECT 121.530 199.440 121.790 199.760 ;
        RECT 121.060 198.565 121.340 198.935 ;
        RECT 120.610 197.740 120.870 198.060 ;
        RECT 120.140 197.460 120.420 197.575 ;
        RECT 121.070 197.460 121.330 197.720 ;
        RECT 120.140 197.400 121.330 197.460 ;
        RECT 119.690 197.060 119.950 197.380 ;
        RECT 120.140 197.320 121.270 197.400 ;
        RECT 120.140 197.205 120.420 197.320 ;
        RECT 118.770 196.380 119.030 196.700 ;
        RECT 118.590 195.505 120.130 195.875 ;
        RECT 120.600 195.165 120.880 195.535 ;
        RECT 117.850 193.660 118.110 193.980 ;
        RECT 119.680 193.805 119.960 194.175 ;
        RECT 117.850 191.280 118.110 191.600 ;
        RECT 117.910 190.775 118.050 191.280 ;
        RECT 119.750 191.260 119.890 193.805 ;
        RECT 119.690 190.940 119.950 191.260 ;
        RECT 117.840 190.405 118.120 190.775 ;
        RECT 117.390 188.560 117.650 188.880 ;
        RECT 117.910 188.200 118.050 190.405 ;
        RECT 118.590 190.065 120.130 190.435 ;
        RECT 120.150 189.580 120.410 189.900 ;
        RECT 118.770 189.240 119.030 189.560 ;
        RECT 117.850 187.880 118.110 188.200 ;
        RECT 117.390 186.860 117.650 187.180 ;
        RECT 117.450 184.120 117.590 186.860 ;
        RECT 118.830 186.500 118.970 189.240 ;
        RECT 119.690 188.900 119.950 189.220 ;
        RECT 119.750 186.500 119.890 188.900 ;
        RECT 118.770 186.180 119.030 186.500 ;
        RECT 119.690 186.180 119.950 186.500 ;
        RECT 120.210 186.160 120.350 189.580 ;
        RECT 120.150 185.840 120.410 186.160 ;
        RECT 118.590 184.625 120.130 184.995 ;
        RECT 117.390 183.800 117.650 184.120 ;
        RECT 116.010 182.440 116.270 182.760 ;
        RECT 116.010 180.060 116.270 180.380 ;
        RECT 116.070 178.000 116.210 180.060 ;
        RECT 116.010 177.680 116.270 178.000 ;
        RECT 116.070 174.940 116.210 177.680 ;
        RECT 116.530 177.660 116.670 183.605 ;
        RECT 116.930 183.460 117.190 183.780 ;
        RECT 119.230 183.460 119.490 183.780 ;
        RECT 119.290 181.740 119.430 183.460 ;
        RECT 119.690 182.780 119.950 183.100 ;
        RECT 120.150 182.780 120.410 183.100 ;
        RECT 119.750 181.935 119.890 182.780 ;
        RECT 119.230 181.420 119.490 181.740 ;
        RECT 119.680 181.565 119.960 181.935 ;
        RECT 119.290 180.720 119.430 181.420 ;
        RECT 119.230 180.400 119.490 180.720 ;
        RECT 120.210 180.040 120.350 182.780 ;
        RECT 117.850 179.720 118.110 180.040 ;
        RECT 120.150 179.720 120.410 180.040 ;
        RECT 117.910 178.340 118.050 179.720 ;
        RECT 118.590 179.185 120.130 179.555 ;
        RECT 117.850 178.020 118.110 178.340 ;
        RECT 118.310 178.020 118.570 178.340 ;
        RECT 120.150 178.020 120.410 178.340 ;
        RECT 116.470 177.340 116.730 177.660 ;
        RECT 116.010 174.620 116.270 174.940 ;
        RECT 117.910 174.600 118.050 178.020 ;
        RECT 118.370 176.300 118.510 178.020 ;
        RECT 118.310 175.980 118.570 176.300 ;
        RECT 115.610 174.200 116.210 174.340 ;
        RECT 117.850 174.280 118.110 174.600 ;
        RECT 120.210 174.510 120.350 178.020 ;
        RECT 120.670 175.620 120.810 195.165 ;
        RECT 121.130 195.000 121.270 197.320 ;
        RECT 121.590 195.000 121.730 199.440 ;
        RECT 122.050 195.000 122.190 211.000 ;
        RECT 122.510 203.500 122.650 216.100 ;
        RECT 122.970 213.700 123.110 221.200 ;
        RECT 130.260 221.005 130.540 221.375 ;
        RECT 134.410 221.200 134.670 221.520 ;
        RECT 123.360 220.325 123.640 220.695 ;
        RECT 126.590 220.520 126.850 220.840 ;
        RECT 123.430 218.800 123.570 220.325 ;
        RECT 123.370 218.480 123.630 218.800 ;
        RECT 124.290 218.480 124.550 218.800 ;
        RECT 124.350 218.120 124.490 218.480 ;
        RECT 124.290 217.800 124.550 218.120 ;
        RECT 123.360 214.885 123.640 215.255 ;
        RECT 123.430 214.380 123.570 214.885 ;
        RECT 123.370 214.060 123.630 214.380 ;
        RECT 122.910 213.380 123.170 213.700 ;
        RECT 122.450 203.180 122.710 203.500 ;
        RECT 122.450 202.500 122.710 202.820 ;
        RECT 122.510 200.100 122.650 202.500 ;
        RECT 122.450 199.780 122.710 200.100 ;
        RECT 121.070 194.680 121.330 195.000 ;
        RECT 121.530 194.680 121.790 195.000 ;
        RECT 121.990 194.680 122.250 195.000 ;
        RECT 121.070 192.300 121.330 192.620 ;
        RECT 121.130 189.560 121.270 192.300 ;
        RECT 121.590 189.900 121.730 194.680 ;
        RECT 122.050 192.620 122.190 194.680 ;
        RECT 122.970 193.640 123.110 213.380 ;
        RECT 123.430 211.320 123.570 214.060 ;
        RECT 124.350 213.020 124.490 217.800 ;
        RECT 126.650 216.420 126.790 220.520 ;
        RECT 129.350 218.820 129.610 219.140 ;
        RECT 129.410 218.540 129.550 218.820 ;
        RECT 130.330 218.800 130.470 221.005 ;
        RECT 133.020 220.325 133.300 220.695 ;
        RECT 133.090 218.800 133.230 220.325 ;
        RECT 129.410 218.400 130.010 218.540 ;
        RECT 130.270 218.480 130.530 218.800 ;
        RECT 133.030 218.480 133.290 218.800 ;
        RECT 129.350 217.800 129.610 218.120 ;
        RECT 125.670 216.100 125.930 216.420 ;
        RECT 126.590 216.100 126.850 216.420 ;
        RECT 127.040 216.245 127.320 216.615 ;
        RECT 127.050 216.100 127.310 216.245 ;
        RECT 127.510 216.100 127.770 216.420 ;
        RECT 128.430 216.100 128.690 216.420 ;
        RECT 128.890 216.100 129.150 216.420 ;
        RECT 125.730 214.380 125.870 216.100 ;
        RECT 125.670 214.060 125.930 214.380 ;
        RECT 127.570 214.040 127.710 216.100 ;
        RECT 127.970 215.420 128.230 215.740 ;
        RECT 127.510 213.720 127.770 214.040 ;
        RECT 128.030 213.700 128.170 215.420 ;
        RECT 127.970 213.380 128.230 213.700 ;
        RECT 124.750 213.040 125.010 213.360 ;
        RECT 124.290 212.700 124.550 213.020 ;
        RECT 123.370 211.000 123.630 211.320 ;
        RECT 123.830 210.660 124.090 210.980 ;
        RECT 123.890 209.135 124.030 210.660 ;
        RECT 123.820 208.765 124.100 209.135 ;
        RECT 124.350 208.940 124.490 212.700 ;
        RECT 124.810 211.660 124.950 213.040 ;
        RECT 128.490 212.680 128.630 216.100 ;
        RECT 126.590 212.360 126.850 212.680 ;
        RECT 128.430 212.360 128.690 212.680 ;
        RECT 124.750 211.340 125.010 211.660 ;
        RECT 126.650 210.980 126.790 212.360 ;
        RECT 126.590 210.660 126.850 210.980 ;
        RECT 127.970 210.660 128.230 210.980 ;
        RECT 125.670 210.320 125.930 210.640 ;
        RECT 124.290 208.620 124.550 208.940 ;
        RECT 123.830 208.280 124.090 208.600 ;
        RECT 123.370 207.600 123.630 207.920 ;
        RECT 123.430 206.220 123.570 207.600 ;
        RECT 123.370 205.900 123.630 206.220 ;
        RECT 123.890 203.410 124.030 208.280 ;
        RECT 124.350 204.520 124.490 208.620 ;
        RECT 125.730 208.600 125.870 210.320 ;
        RECT 125.670 208.280 125.930 208.600 ;
        RECT 124.750 205.055 125.010 205.200 ;
        RECT 124.740 204.685 125.020 205.055 ;
        RECT 125.210 204.880 125.470 205.200 ;
        RECT 125.670 204.880 125.930 205.200 ;
        RECT 124.290 204.200 124.550 204.520 ;
        RECT 124.290 203.410 124.550 203.500 ;
        RECT 123.890 203.270 124.550 203.410 ;
        RECT 124.290 203.180 124.550 203.270 ;
        RECT 123.360 201.965 123.640 202.335 ;
        RECT 124.290 202.160 124.550 202.480 ;
        RECT 123.370 201.820 123.630 201.965 ;
        RECT 124.350 200.295 124.490 202.160 ;
        RECT 125.270 200.780 125.410 204.880 ;
        RECT 125.210 200.460 125.470 200.780 ;
        RECT 124.280 199.925 124.560 200.295 ;
        RECT 124.290 199.780 124.550 199.925 ;
        RECT 124.290 198.760 124.550 199.080 ;
        RECT 124.350 198.255 124.490 198.760 ;
        RECT 123.370 197.740 123.630 198.060 ;
        RECT 124.280 197.885 124.560 198.255 ;
        RECT 123.430 195.340 123.570 197.740 ;
        RECT 123.370 195.020 123.630 195.340 ;
        RECT 122.910 193.320 123.170 193.640 ;
        RECT 121.990 192.300 122.250 192.620 ;
        RECT 121.990 190.600 122.250 190.920 ;
        RECT 121.530 189.580 121.790 189.900 ;
        RECT 121.070 189.240 121.330 189.560 ;
        RECT 121.070 188.220 121.330 188.540 ;
        RECT 121.130 188.055 121.270 188.220 ;
        RECT 121.060 187.685 121.340 188.055 ;
        RECT 121.590 186.500 121.730 189.580 ;
        RECT 122.050 189.220 122.190 190.600 ;
        RECT 124.350 189.900 124.490 197.885 ;
        RECT 125.210 194.910 125.470 195.000 ;
        RECT 124.810 194.770 125.470 194.910 ;
        RECT 123.370 189.580 123.630 189.900 ;
        RECT 124.290 189.580 124.550 189.900 ;
        RECT 121.990 188.900 122.250 189.220 ;
        RECT 121.530 186.180 121.790 186.500 ;
        RECT 121.070 185.500 121.330 185.820 ;
        RECT 121.130 185.335 121.270 185.500 ;
        RECT 121.060 184.965 121.340 185.335 ;
        RECT 121.590 178.680 121.730 186.180 ;
        RECT 122.050 181.740 122.190 188.900 ;
        RECT 123.430 188.540 123.570 189.580 ;
        RECT 122.910 188.220 123.170 188.540 ;
        RECT 123.370 188.220 123.630 188.540 ;
        RECT 122.440 187.685 122.720 188.055 ;
        RECT 122.510 185.480 122.650 187.685 ;
        RECT 122.450 185.160 122.710 185.480 ;
        RECT 121.990 181.420 122.250 181.740 ;
        RECT 122.510 181.400 122.650 185.160 ;
        RECT 122.970 181.400 123.110 188.220 ;
        RECT 124.280 185.645 124.560 186.015 ;
        RECT 123.370 184.140 123.630 184.460 ;
        RECT 122.450 181.080 122.710 181.400 ;
        RECT 122.910 181.080 123.170 181.400 ;
        RECT 121.980 180.205 122.260 180.575 ;
        RECT 121.990 180.060 122.250 180.205 ;
        RECT 121.530 178.360 121.790 178.680 ;
        RECT 121.070 178.020 121.330 178.340 ;
        RECT 120.610 175.300 120.870 175.620 ;
        RECT 120.210 174.370 120.810 174.510 ;
        RECT 113.250 172.580 113.510 172.900 ;
        RECT 113.310 172.415 113.450 172.580 ;
        RECT 112.790 171.900 113.050 172.220 ;
        RECT 113.240 172.045 113.520 172.415 ;
        RECT 112.850 170.860 112.990 171.900 ;
        RECT 114.170 171.560 114.430 171.880 ;
        RECT 112.790 170.540 113.050 170.860 ;
        RECT 114.230 169.695 114.370 171.560 ;
        RECT 114.160 169.325 114.440 169.695 ;
        RECT 115.090 166.800 115.350 167.120 ;
        RECT 114.630 166.120 114.890 166.440 ;
        RECT 114.690 164.060 114.830 166.120 ;
        RECT 115.150 164.740 115.290 166.800 ;
        RECT 115.090 164.420 115.350 164.740 ;
        RECT 114.630 163.740 114.890 164.060 ;
        RECT 113.250 162.380 113.510 162.700 ;
        RECT 113.310 161.680 113.450 162.380 ;
        RECT 114.690 162.360 114.830 163.740 ;
        RECT 115.550 163.400 115.810 163.720 ;
        RECT 114.630 162.040 114.890 162.360 ;
        RECT 112.330 161.360 112.590 161.680 ;
        RECT 113.250 161.360 113.510 161.680 ;
        RECT 109.570 158.640 109.830 158.960 ;
        RECT 110.030 158.300 110.290 158.620 ;
        RECT 109.110 155.920 109.370 156.240 ;
        RECT 110.090 153.520 110.230 158.300 ;
        RECT 112.790 157.960 113.050 158.280 ;
        RECT 112.850 156.920 112.990 157.960 ;
        RECT 112.790 156.600 113.050 156.920 ;
        RECT 111.870 156.490 112.130 156.580 ;
        RECT 111.870 156.350 112.530 156.490 ;
        RECT 111.870 156.260 112.130 156.350 ;
        RECT 110.950 155.920 111.210 156.240 ;
        RECT 110.030 153.200 110.290 153.520 ;
        RECT 108.650 152.520 108.910 152.840 ;
        RECT 108.710 150.655 108.850 152.520 ;
        RECT 108.640 150.285 108.920 150.655 ;
        RECT 109.570 150.480 109.830 150.800 ;
        RECT 108.190 147.420 108.450 147.740 ;
        RECT 108.250 145.700 108.390 147.420 ;
        RECT 108.190 145.380 108.450 145.700 ;
        RECT 108.710 142.980 108.850 150.285 ;
        RECT 109.630 148.080 109.770 150.480 ;
        RECT 109.570 147.760 109.830 148.080 ;
        RECT 109.630 146.040 109.770 147.760 ;
        RECT 109.570 145.720 109.830 146.040 ;
        RECT 111.010 145.020 111.150 155.920 ;
        RECT 112.390 153.520 112.530 156.350 ;
        RECT 112.850 153.860 112.990 156.600 ;
        RECT 112.790 153.540 113.050 153.860 ;
        RECT 112.330 153.200 112.590 153.520 ;
        RECT 111.860 150.965 112.140 151.335 ;
        RECT 111.870 150.820 112.130 150.965 ;
        RECT 112.390 148.080 112.530 153.200 ;
        RECT 111.410 147.990 111.670 148.080 ;
        RECT 111.410 147.850 112.070 147.990 ;
        RECT 111.410 147.760 111.670 147.850 ;
        RECT 111.410 147.080 111.670 147.400 ;
        RECT 110.950 144.700 111.210 145.020 ;
        RECT 109.100 144.165 109.380 144.535 ;
        RECT 108.650 142.660 108.910 142.980 ;
        RECT 108.190 141.980 108.450 142.300 ;
        RECT 108.250 140.260 108.390 141.980 ;
        RECT 108.710 140.260 108.850 142.660 ;
        RECT 109.170 142.640 109.310 144.165 ;
        RECT 110.020 143.485 110.300 143.855 ;
        RECT 110.090 142.640 110.230 143.485 ;
        RECT 109.110 142.320 109.370 142.640 ;
        RECT 110.030 142.320 110.290 142.640 ;
        RECT 110.490 142.320 110.750 142.640 ;
        RECT 109.170 140.260 109.310 142.320 ;
        RECT 108.190 139.940 108.450 140.260 ;
        RECT 108.650 139.940 108.910 140.260 ;
        RECT 109.110 139.940 109.370 140.260 ;
        RECT 108.250 137.880 108.390 139.940 ;
        RECT 108.710 138.220 108.850 139.940 ;
        RECT 109.570 139.260 109.830 139.580 ;
        RECT 108.650 137.900 108.910 138.220 ;
        RECT 108.190 137.560 108.450 137.880 ;
        RECT 108.650 136.200 108.910 136.520 ;
        RECT 109.110 136.200 109.370 136.520 ;
        RECT 108.710 135.160 108.850 136.200 ;
        RECT 109.170 135.500 109.310 136.200 ;
        RECT 109.630 135.500 109.770 139.260 ;
        RECT 110.550 137.540 110.690 142.320 ;
        RECT 110.950 141.640 111.210 141.960 ;
        RECT 110.490 137.220 110.750 137.540 ;
        RECT 110.480 136.940 110.760 137.055 ;
        RECT 110.090 136.800 110.760 136.940 ;
        RECT 109.110 135.180 109.370 135.500 ;
        RECT 109.570 135.180 109.830 135.500 ;
        RECT 108.650 134.840 108.910 135.160 ;
        RECT 109.110 133.820 109.370 134.140 ;
        RECT 109.170 132.860 109.310 133.820 ;
        RECT 110.090 132.860 110.230 136.800 ;
        RECT 110.480 136.685 110.760 136.800 ;
        RECT 109.170 132.720 110.230 132.860 ;
        RECT 109.170 131.760 109.310 132.720 ;
        RECT 110.030 131.780 110.290 132.100 ;
        RECT 107.790 131.360 108.390 131.500 ;
        RECT 109.110 131.440 109.370 131.760 ;
        RECT 109.560 131.500 109.840 131.615 ;
        RECT 110.090 131.500 110.230 131.780 ;
        RECT 111.010 131.500 111.150 141.640 ;
        RECT 111.470 139.580 111.610 147.080 ;
        RECT 111.930 140.940 112.070 147.850 ;
        RECT 112.330 147.760 112.590 148.080 ;
        RECT 112.390 146.040 112.530 147.760 ;
        RECT 113.310 147.740 113.450 161.360 ;
        RECT 115.610 159.495 115.750 163.400 ;
        RECT 114.160 159.125 114.440 159.495 ;
        RECT 115.540 159.125 115.820 159.495 ;
        RECT 113.710 156.260 113.970 156.580 ;
        RECT 113.770 152.015 113.910 156.260 ;
        RECT 113.700 151.645 113.980 152.015 ;
        RECT 113.770 151.480 113.910 151.645 ;
        RECT 113.710 151.160 113.970 151.480 ;
        RECT 113.250 147.420 113.510 147.740 ;
        RECT 112.790 147.080 113.050 147.400 ;
        RECT 112.330 145.720 112.590 146.040 ;
        RECT 112.390 142.980 112.530 145.720 ;
        RECT 112.330 142.660 112.590 142.980 ;
        RECT 112.330 141.815 112.590 141.960 ;
        RECT 112.320 141.445 112.600 141.815 ;
        RECT 111.870 140.620 112.130 140.940 ;
        RECT 111.410 139.260 111.670 139.580 ;
        RECT 111.470 138.220 111.610 139.260 ;
        RECT 111.410 137.900 111.670 138.220 ;
        RECT 111.470 134.820 111.610 137.900 ;
        RECT 111.870 136.880 112.130 137.200 ;
        RECT 112.390 136.940 112.530 141.445 ;
        RECT 112.850 140.260 112.990 147.080 ;
        RECT 113.240 145.525 113.520 145.895 ;
        RECT 113.310 145.360 113.450 145.525 ;
        RECT 113.250 145.040 113.510 145.360 ;
        RECT 114.230 145.215 114.370 159.125 ;
        RECT 115.550 156.600 115.810 156.920 ;
        RECT 115.610 154.540 115.750 156.600 ;
        RECT 115.550 154.220 115.810 154.540 ;
        RECT 116.070 154.055 116.210 174.200 ;
        RECT 118.590 173.745 120.130 174.115 ;
        RECT 120.670 173.580 120.810 174.370 ;
        RECT 120.610 173.260 120.870 173.580 ;
        RECT 118.760 172.725 119.040 173.095 ;
        RECT 118.770 172.580 119.030 172.725 ;
        RECT 120.150 172.580 120.410 172.900 ;
        RECT 116.930 172.240 117.190 172.560 ;
        RECT 116.470 169.180 116.730 169.500 ;
        RECT 116.530 161.340 116.670 169.180 ;
        RECT 116.990 169.160 117.130 172.240 ;
        RECT 118.770 171.900 119.030 172.220 ;
        RECT 117.850 171.560 118.110 171.880 ;
        RECT 118.830 171.735 118.970 171.900 ;
        RECT 117.910 170.860 118.050 171.560 ;
        RECT 118.760 171.365 119.040 171.735 ;
        RECT 120.210 170.860 120.350 172.580 ;
        RECT 120.670 172.560 120.810 173.260 ;
        RECT 121.130 172.560 121.270 178.020 ;
        RECT 121.520 177.485 121.800 177.855 ;
        RECT 121.990 177.680 122.250 178.000 ;
        RECT 121.590 177.320 121.730 177.485 ;
        RECT 121.530 177.000 121.790 177.320 ;
        RECT 122.050 174.600 122.190 177.680 ;
        RECT 122.970 176.300 123.110 181.080 ;
        RECT 123.430 178.340 123.570 184.140 ;
        RECT 124.350 184.120 124.490 185.645 ;
        RECT 124.290 183.800 124.550 184.120 ;
        RECT 123.830 183.460 124.090 183.780 ;
        RECT 123.890 180.720 124.030 183.460 ;
        RECT 124.290 182.440 124.550 182.760 ;
        RECT 124.350 181.400 124.490 182.440 ;
        RECT 124.290 181.080 124.550 181.400 ;
        RECT 123.830 180.400 124.090 180.720 ;
        RECT 123.370 178.020 123.630 178.340 ;
        RECT 122.910 175.980 123.170 176.300 ;
        RECT 122.440 174.765 122.720 175.135 ;
        RECT 123.890 174.940 124.030 180.400 ;
        RECT 124.290 179.720 124.550 180.040 ;
        RECT 124.350 176.300 124.490 179.720 ;
        RECT 124.810 179.020 124.950 194.770 ;
        RECT 125.210 194.680 125.470 194.770 ;
        RECT 125.210 188.900 125.470 189.220 ;
        RECT 125.270 179.020 125.410 188.900 ;
        RECT 125.730 186.160 125.870 204.880 ;
        RECT 126.130 201.480 126.390 201.800 ;
        RECT 126.190 195.535 126.330 201.480 ;
        RECT 126.650 200.100 126.790 210.660 ;
        RECT 127.050 201.820 127.310 202.140 ;
        RECT 126.590 199.780 126.850 200.100 ;
        RECT 126.650 197.720 126.790 199.780 ;
        RECT 126.590 197.400 126.850 197.720 ;
        RECT 126.590 196.215 126.850 196.360 ;
        RECT 126.580 195.845 126.860 196.215 ;
        RECT 126.120 195.165 126.400 195.535 ;
        RECT 126.130 194.680 126.390 195.000 ;
        RECT 126.190 193.640 126.330 194.680 ;
        RECT 126.130 193.320 126.390 193.640 ;
        RECT 127.110 189.300 127.250 201.820 ;
        RECT 127.510 197.400 127.770 197.720 ;
        RECT 127.570 193.980 127.710 197.400 ;
        RECT 127.510 193.660 127.770 193.980 ;
        RECT 127.570 192.135 127.710 193.660 ;
        RECT 127.500 191.765 127.780 192.135 ;
        RECT 126.650 189.160 127.250 189.300 ;
        RECT 126.130 188.560 126.390 188.880 ;
        RECT 126.650 188.735 126.790 189.160 ;
        RECT 125.670 185.840 125.930 186.160 ;
        RECT 126.190 183.780 126.330 188.560 ;
        RECT 126.580 188.365 126.860 188.735 ;
        RECT 127.050 188.560 127.310 188.880 ;
        RECT 126.590 187.880 126.850 188.200 ;
        RECT 126.650 186.160 126.790 187.880 ;
        RECT 127.110 186.840 127.250 188.560 ;
        RECT 127.050 186.520 127.310 186.840 ;
        RECT 126.590 185.840 126.850 186.160 ;
        RECT 126.130 183.690 126.390 183.780 ;
        RECT 125.730 183.550 126.390 183.690 ;
        RECT 124.750 178.700 125.010 179.020 ;
        RECT 125.210 178.700 125.470 179.020 ;
        RECT 124.290 175.980 124.550 176.300 ;
        RECT 125.210 175.980 125.470 176.300 ;
        RECT 124.290 174.960 124.550 175.280 ;
        RECT 121.990 174.280 122.250 174.600 ;
        RECT 122.050 173.580 122.190 174.280 ;
        RECT 121.990 173.260 122.250 173.580 ;
        RECT 120.610 172.240 120.870 172.560 ;
        RECT 121.070 172.240 121.330 172.560 ;
        RECT 117.390 170.540 117.650 170.860 ;
        RECT 117.850 170.540 118.110 170.860 ;
        RECT 120.150 170.540 120.410 170.860 ;
        RECT 116.930 168.840 117.190 169.160 ;
        RECT 116.930 164.420 117.190 164.740 ;
        RECT 116.990 162.020 117.130 164.420 ;
        RECT 117.450 164.060 117.590 170.540 ;
        RECT 121.530 169.180 121.790 169.500 ;
        RECT 118.590 168.305 120.130 168.675 ;
        RECT 120.610 166.860 120.870 167.120 ;
        RECT 121.590 166.860 121.730 169.180 ;
        RECT 120.610 166.800 121.730 166.860 ;
        RECT 120.670 166.720 121.730 166.800 ;
        RECT 117.390 163.740 117.650 164.060 ;
        RECT 118.590 162.865 120.130 163.235 ;
        RECT 116.930 161.700 117.190 162.020 ;
        RECT 119.230 161.700 119.490 162.020 ;
        RECT 119.690 161.700 119.950 162.020 ;
        RECT 121.590 161.930 121.730 166.720 ;
        RECT 122.050 165.420 122.190 173.260 ;
        RECT 122.510 172.900 122.650 174.765 ;
        RECT 123.830 174.620 124.090 174.940 ;
        RECT 123.370 174.280 123.630 174.600 ;
        RECT 123.430 173.660 123.570 174.280 ;
        RECT 123.820 173.660 124.100 173.775 ;
        RECT 123.430 173.520 124.100 173.660 ;
        RECT 123.820 173.405 124.100 173.520 ;
        RECT 122.450 172.580 122.710 172.900 ;
        RECT 124.350 172.300 124.490 174.960 ;
        RECT 125.270 174.940 125.410 175.980 ;
        RECT 125.730 175.620 125.870 183.550 ;
        RECT 126.130 183.460 126.390 183.550 ;
        RECT 126.120 182.925 126.400 183.295 ;
        RECT 126.190 180.380 126.330 182.925 ;
        RECT 126.650 180.575 126.790 185.840 ;
        RECT 126.130 180.060 126.390 180.380 ;
        RECT 126.580 180.205 126.860 180.575 ;
        RECT 127.050 180.400 127.310 180.720 ;
        RECT 125.670 175.300 125.930 175.620 ;
        RECT 125.210 174.620 125.470 174.940 ;
        RECT 125.730 173.150 125.870 175.300 ;
        RECT 127.110 175.280 127.250 180.400 ;
        RECT 128.030 178.340 128.170 210.660 ;
        RECT 128.490 202.140 128.630 212.360 ;
        RECT 128.430 201.820 128.690 202.140 ;
        RECT 128.950 200.860 129.090 216.100 ;
        RECT 129.410 207.920 129.550 217.800 ;
        RECT 129.350 207.600 129.610 207.920 ;
        RECT 129.350 202.840 129.610 203.160 ;
        RECT 129.410 202.140 129.550 202.840 ;
        RECT 129.350 201.820 129.610 202.140 ;
        RECT 128.950 200.720 129.550 200.860 ;
        RECT 128.890 200.010 129.150 200.100 ;
        RECT 128.490 199.870 129.150 200.010 ;
        RECT 128.490 191.940 128.630 199.870 ;
        RECT 128.890 199.780 129.150 199.870 ;
        RECT 128.890 199.100 129.150 199.420 ;
        RECT 128.950 195.340 129.090 199.100 ;
        RECT 128.890 195.020 129.150 195.340 ;
        RECT 128.890 193.660 129.150 193.980 ;
        RECT 128.950 192.620 129.090 193.660 ;
        RECT 128.890 192.300 129.150 192.620 ;
        RECT 128.430 191.620 128.690 191.940 ;
        RECT 128.890 191.620 129.150 191.940 ;
        RECT 128.490 188.880 128.630 191.620 ;
        RECT 128.430 188.560 128.690 188.880 ;
        RECT 128.430 186.695 128.690 186.840 ;
        RECT 128.420 186.325 128.700 186.695 ;
        RECT 128.950 184.120 129.090 191.620 ;
        RECT 129.410 187.375 129.550 200.720 ;
        RECT 129.340 187.005 129.620 187.375 ;
        RECT 128.890 183.800 129.150 184.120 ;
        RECT 129.410 183.780 129.550 187.005 ;
        RECT 129.350 183.460 129.610 183.780 ;
        RECT 129.350 182.780 129.610 183.100 ;
        RECT 129.410 179.020 129.550 182.780 ;
        RECT 128.890 178.700 129.150 179.020 ;
        RECT 129.350 178.700 129.610 179.020 ;
        RECT 128.950 178.420 129.090 178.700 ;
        RECT 127.970 178.020 128.230 178.340 ;
        RECT 128.950 178.280 129.550 178.420 ;
        RECT 128.030 176.300 128.170 178.020 ;
        RECT 128.890 177.000 129.150 177.320 ;
        RECT 128.950 176.300 129.090 177.000 ;
        RECT 129.410 176.300 129.550 178.280 ;
        RECT 127.970 175.980 128.230 176.300 ;
        RECT 128.890 175.980 129.150 176.300 ;
        RECT 129.350 175.980 129.610 176.300 ;
        RECT 127.050 174.960 127.310 175.280 ;
        RECT 128.420 173.405 128.700 173.775 ;
        RECT 128.490 173.240 128.630 173.405 ;
        RECT 126.130 173.150 126.390 173.240 ;
        RECT 125.730 173.010 126.390 173.150 ;
        RECT 126.130 172.920 126.390 173.010 ;
        RECT 128.430 172.920 128.690 173.240 ;
        RECT 124.350 172.220 125.410 172.300 ;
        RECT 124.350 172.160 125.470 172.220 ;
        RECT 125.210 171.900 125.470 172.160 ;
        RECT 124.280 170.005 124.560 170.375 ;
        RECT 124.350 169.840 124.490 170.005 ;
        RECT 124.290 169.520 124.550 169.840 ;
        RECT 123.830 168.840 124.090 169.160 ;
        RECT 123.370 167.480 123.630 167.800 ;
        RECT 122.900 166.605 123.180 166.975 ;
        RECT 122.970 165.420 123.110 166.605 ;
        RECT 123.430 166.440 123.570 167.480 ;
        RECT 123.370 166.120 123.630 166.440 ;
        RECT 121.990 165.100 122.250 165.420 ;
        RECT 122.910 165.100 123.170 165.420 ;
        RECT 122.970 162.700 123.110 165.100 ;
        RECT 122.910 162.380 123.170 162.700 ;
        RECT 122.910 161.930 123.170 162.020 ;
        RECT 121.590 161.790 123.170 161.930 ;
        RECT 122.910 161.700 123.170 161.790 ;
        RECT 118.310 161.535 118.570 161.680 ;
        RECT 116.470 161.250 116.730 161.340 ;
        RECT 116.470 161.110 117.590 161.250 ;
        RECT 118.300 161.165 118.580 161.535 ;
        RECT 118.770 161.250 119.030 161.340 ;
        RECT 119.290 161.250 119.430 161.700 ;
        RECT 116.470 161.020 116.730 161.110 ;
        RECT 116.930 159.660 117.190 159.980 ;
        RECT 116.990 158.960 117.130 159.660 ;
        RECT 117.450 159.640 117.590 161.110 ;
        RECT 118.770 161.110 119.430 161.250 ;
        RECT 118.770 161.020 119.030 161.110 ;
        RECT 119.750 161.000 119.890 161.700 ;
        RECT 121.060 161.165 121.340 161.535 ;
        RECT 119.690 160.680 119.950 161.000 ;
        RECT 117.390 159.320 117.650 159.640 ;
        RECT 117.850 159.320 118.110 159.640 ;
        RECT 116.930 158.640 117.190 158.960 ;
        RECT 116.470 157.960 116.730 158.280 ;
        RECT 115.550 153.540 115.810 153.860 ;
        RECT 116.000 153.685 116.280 154.055 ;
        RECT 116.530 153.860 116.670 157.960 ;
        RECT 116.010 153.540 116.270 153.685 ;
        RECT 116.470 153.540 116.730 153.860 ;
        RECT 115.610 153.260 115.750 153.540 ;
        RECT 117.450 153.260 117.590 159.320 ;
        RECT 117.910 154.540 118.050 159.320 ;
        RECT 120.610 158.640 120.870 158.960 ;
        RECT 118.590 157.425 120.130 157.795 ;
        RECT 120.670 157.260 120.810 158.640 ;
        RECT 120.610 156.940 120.870 157.260 ;
        RECT 118.770 155.920 119.030 156.240 ;
        RECT 121.130 156.095 121.270 161.165 ;
        RECT 121.980 160.485 122.260 160.855 ;
        RECT 122.050 159.300 122.190 160.485 ;
        RECT 121.990 158.980 122.250 159.300 ;
        RECT 121.530 158.640 121.790 158.960 ;
        RECT 123.430 158.700 123.570 166.120 ;
        RECT 123.890 162.020 124.030 168.840 ;
        RECT 124.750 166.120 125.010 166.440 ;
        RECT 124.810 164.935 124.950 166.120 ;
        RECT 124.740 164.565 125.020 164.935 ;
        RECT 128.890 163.740 129.150 164.060 ;
        RECT 128.430 163.400 128.690 163.720 ;
        RECT 128.490 162.700 128.630 163.400 ;
        RECT 128.430 162.380 128.690 162.700 ;
        RECT 123.830 161.700 124.090 162.020 ;
        RECT 127.050 161.700 127.310 162.020 ;
        RECT 117.850 154.220 118.110 154.540 ;
        RECT 118.830 153.860 118.970 155.920 ;
        RECT 121.060 155.725 121.340 156.095 ;
        RECT 119.690 154.220 119.950 154.540 ;
        RECT 118.770 153.540 119.030 153.860 ;
        RECT 115.610 153.120 117.590 153.260 ;
        RECT 119.750 153.180 119.890 154.220 ;
        RECT 119.690 152.860 119.950 153.180 ;
        RECT 116.930 152.520 117.190 152.840 ;
        RECT 117.850 152.520 118.110 152.840 ;
        RECT 116.990 150.800 117.130 152.520 ;
        RECT 117.910 151.480 118.050 152.520 ;
        RECT 118.590 151.985 120.130 152.355 ;
        RECT 120.610 151.500 120.870 151.820 ;
        RECT 117.850 151.390 118.110 151.480 ;
        RECT 117.850 151.250 118.510 151.390 ;
        RECT 117.850 151.160 118.110 151.250 ;
        RECT 114.630 150.480 114.890 150.800 ;
        RECT 116.930 150.480 117.190 150.800 ;
        RECT 114.690 146.040 114.830 150.480 ;
        RECT 115.550 149.860 115.810 150.120 ;
        RECT 116.990 149.975 117.130 150.480 ;
        RECT 115.150 149.800 115.810 149.860 ;
        RECT 115.150 149.720 115.750 149.800 ;
        RECT 115.150 148.760 115.290 149.720 ;
        RECT 116.920 149.605 117.200 149.975 ;
        RECT 117.850 149.800 118.110 150.120 ;
        RECT 116.010 148.780 116.270 149.100 ;
        RECT 115.090 148.440 115.350 148.760 ;
        RECT 116.070 148.080 116.210 148.780 ;
        RECT 116.010 147.760 116.270 148.080 ;
        RECT 114.630 145.720 114.890 146.040 ;
        RECT 114.160 144.845 114.440 145.215 ;
        RECT 114.230 142.300 114.370 144.845 ;
        RECT 114.170 141.980 114.430 142.300 ;
        RECT 116.070 140.940 116.210 147.760 ;
        RECT 117.390 147.080 117.650 147.400 ;
        RECT 116.470 145.720 116.730 146.040 ;
        RECT 114.630 140.620 114.890 140.940 ;
        RECT 116.010 140.620 116.270 140.940 ;
        RECT 116.530 140.850 116.670 145.720 ;
        RECT 117.450 145.020 117.590 147.080 ;
        RECT 117.910 145.700 118.050 149.800 ;
        RECT 118.370 149.100 118.510 151.250 ;
        RECT 119.230 150.480 119.490 150.800 ;
        RECT 118.310 148.780 118.570 149.100 ;
        RECT 118.770 148.780 119.030 149.100 ;
        RECT 118.830 148.080 118.970 148.780 ;
        RECT 119.290 148.080 119.430 150.480 ;
        RECT 120.670 148.670 120.810 151.500 ;
        RECT 121.130 151.220 121.270 155.725 ;
        RECT 121.590 154.540 121.730 158.640 ;
        RECT 122.510 158.560 123.570 158.700 ;
        RECT 121.990 157.960 122.250 158.280 ;
        RECT 121.530 154.220 121.790 154.540 ;
        RECT 121.130 151.080 121.730 151.220 ;
        RECT 121.070 148.670 121.330 148.760 ;
        RECT 120.670 148.530 121.330 148.670 ;
        RECT 121.070 148.440 121.330 148.530 ;
        RECT 118.770 147.760 119.030 148.080 ;
        RECT 119.230 147.760 119.490 148.080 ;
        RECT 120.610 147.080 120.870 147.400 ;
        RECT 118.590 146.545 120.130 146.915 ;
        RECT 120.670 145.700 120.810 147.080 ;
        RECT 121.590 145.700 121.730 151.080 ;
        RECT 122.050 150.800 122.190 157.960 ;
        RECT 122.510 156.920 122.650 158.560 ;
        RECT 122.450 156.600 122.710 156.920 ;
        RECT 122.510 151.820 122.650 156.600 ;
        RECT 123.890 155.560 124.030 161.700 ;
        RECT 124.750 161.360 125.010 161.680 ;
        RECT 126.130 161.360 126.390 161.680 ;
        RECT 124.810 161.000 124.950 161.360 ;
        RECT 124.750 160.680 125.010 161.000 ;
        RECT 124.750 159.320 125.010 159.640 ;
        RECT 124.290 156.775 124.550 156.920 ;
        RECT 124.280 156.405 124.560 156.775 ;
        RECT 123.830 155.240 124.090 155.560 ;
        RECT 124.290 155.240 124.550 155.560 ;
        RECT 123.370 153.540 123.630 153.860 ;
        RECT 123.430 151.820 123.570 153.540 ;
        RECT 123.890 153.180 124.030 155.240 ;
        RECT 124.350 154.540 124.490 155.240 ;
        RECT 124.290 154.220 124.550 154.540 ;
        RECT 123.830 152.860 124.090 153.180 ;
        RECT 122.450 151.500 122.710 151.820 ;
        RECT 123.370 151.500 123.630 151.820 ;
        RECT 124.810 151.480 124.950 159.320 ;
        RECT 125.670 158.300 125.930 158.620 ;
        RECT 124.750 151.160 125.010 151.480 ;
        RECT 121.990 150.480 122.250 150.800 ;
        RECT 125.730 150.460 125.870 158.300 ;
        RECT 125.670 150.140 125.930 150.460 ;
        RECT 121.990 148.780 122.250 149.100 ;
        RECT 117.850 145.380 118.110 145.700 ;
        RECT 120.610 145.380 120.870 145.700 ;
        RECT 121.070 145.380 121.330 145.700 ;
        RECT 121.530 145.380 121.790 145.700 ;
        RECT 117.390 144.700 117.650 145.020 ;
        RECT 116.530 140.710 117.590 140.850 ;
        RECT 112.790 139.940 113.050 140.260 ;
        RECT 114.170 139.940 114.430 140.260 ;
        RECT 114.230 139.240 114.370 139.940 ;
        RECT 114.170 138.920 114.430 139.240 ;
        RECT 114.230 137.200 114.370 138.920 ;
        RECT 114.690 137.200 114.830 140.620 ;
        RECT 116.070 140.340 116.210 140.620 ;
        RECT 116.070 140.200 117.130 140.340 ;
        RECT 117.450 140.260 117.590 140.710 ;
        RECT 117.910 140.260 118.050 145.380 ;
        RECT 120.600 144.845 120.880 145.215 ;
        RECT 120.140 142.805 120.420 143.175 ;
        RECT 120.210 142.640 120.350 142.805 ;
        RECT 120.150 142.320 120.410 142.640 ;
        RECT 120.670 142.300 120.810 144.845 ;
        RECT 120.610 141.980 120.870 142.300 ;
        RECT 118.590 141.105 120.130 141.475 ;
        RECT 120.670 140.600 120.810 141.980 ;
        RECT 121.130 141.135 121.270 145.380 ;
        RECT 122.050 142.640 122.190 148.780 ;
        RECT 123.370 147.760 123.630 148.080 ;
        RECT 124.750 147.990 125.010 148.080 ;
        RECT 125.730 147.990 125.870 150.140 ;
        RECT 126.190 150.120 126.330 161.360 ;
        RECT 127.110 161.340 127.250 161.700 ;
        RECT 127.050 161.020 127.310 161.340 ;
        RECT 127.960 160.740 128.240 160.855 ;
        RECT 127.570 160.600 128.240 160.740 ;
        RECT 126.590 158.300 126.850 158.620 ;
        RECT 127.050 158.300 127.310 158.620 ;
        RECT 126.650 152.840 126.790 158.300 ;
        RECT 126.590 152.520 126.850 152.840 ;
        RECT 127.110 151.140 127.250 158.300 ;
        RECT 127.050 150.820 127.310 151.140 ;
        RECT 126.130 149.800 126.390 150.120 ;
        RECT 127.110 148.500 127.250 150.820 ;
        RECT 127.570 150.800 127.710 160.600 ;
        RECT 127.960 160.485 128.240 160.600 ;
        RECT 128.430 158.640 128.690 158.960 ;
        RECT 128.490 151.820 128.630 158.640 ;
        RECT 128.950 153.520 129.090 163.740 ;
        RECT 129.350 160.680 129.610 161.000 ;
        RECT 129.410 158.620 129.550 160.680 ;
        RECT 129.350 158.300 129.610 158.620 ;
        RECT 129.410 156.580 129.550 158.300 ;
        RECT 129.870 157.260 130.010 218.400 ;
        RECT 131.650 218.140 131.910 218.460 ;
        RECT 131.710 210.980 131.850 218.140 ;
        RECT 134.470 217.100 134.610 221.200 ;
        RECT 148.660 221.005 148.940 221.375 ;
        RECT 151.890 221.200 152.150 221.520 ;
        RECT 137.160 219.645 137.440 220.015 ;
        RECT 138.025 219.985 139.565 220.355 ;
        RECT 140.380 220.325 140.660 220.695 ;
        RECT 137.230 218.800 137.370 219.645 ;
        RECT 138.540 218.965 138.820 219.335 ;
        RECT 138.610 218.800 138.750 218.965 ;
        RECT 140.450 218.800 140.590 220.325 ;
        RECT 142.230 219.500 142.490 219.820 ;
        RECT 137.170 218.480 137.430 218.800 ;
        RECT 137.630 218.480 137.890 218.800 ;
        RECT 138.550 218.480 138.810 218.800 ;
        RECT 140.390 218.480 140.650 218.800 ;
        RECT 136.250 217.800 136.510 218.120 ;
        RECT 134.410 216.780 134.670 217.100 ;
        RECT 135.330 216.440 135.590 216.760 ;
        RECT 133.490 216.100 133.750 216.420 ;
        RECT 133.550 211.320 133.690 216.100 ;
        RECT 135.390 213.360 135.530 216.440 ;
        RECT 135.330 213.040 135.590 213.360 ;
        RECT 133.950 212.360 134.210 212.680 ;
        RECT 134.870 212.360 135.130 212.680 ;
        RECT 135.790 212.360 136.050 212.680 ;
        RECT 134.010 211.660 134.150 212.360 ;
        RECT 133.950 211.340 134.210 211.660 ;
        RECT 133.490 211.000 133.750 211.320 ;
        RECT 131.650 210.660 131.910 210.980 ;
        RECT 132.570 210.660 132.830 210.980 ;
        RECT 133.030 210.660 133.290 210.980 ;
        RECT 130.270 209.640 130.530 209.960 ;
        RECT 131.710 209.815 131.850 210.660 ;
        RECT 130.330 207.920 130.470 209.640 ;
        RECT 131.640 209.445 131.920 209.815 ;
        RECT 132.630 208.340 132.770 210.660 ;
        RECT 133.090 208.940 133.230 210.660 ;
        RECT 133.950 210.320 134.210 210.640 ;
        RECT 133.030 208.620 133.290 208.940 ;
        RECT 132.630 208.200 133.230 208.340 ;
        RECT 130.270 207.600 130.530 207.920 ;
        RECT 132.110 207.600 132.370 207.920 ;
        RECT 130.730 207.490 130.990 207.580 ;
        RECT 130.730 207.350 131.850 207.490 ;
        RECT 130.730 207.260 130.990 207.350 ;
        RECT 130.730 204.880 130.990 205.200 ;
        RECT 130.790 203.500 130.930 204.880 ;
        RECT 130.730 203.180 130.990 203.500 ;
        RECT 130.270 200.120 130.530 200.440 ;
        RECT 130.330 192.620 130.470 200.120 ;
        RECT 130.270 192.300 130.530 192.620 ;
        RECT 130.330 189.300 130.470 192.300 ;
        RECT 130.790 189.900 130.930 203.180 ;
        RECT 131.190 202.840 131.450 203.160 ;
        RECT 131.250 197.380 131.390 202.840 ;
        RECT 131.190 197.060 131.450 197.380 ;
        RECT 131.180 196.525 131.460 196.895 ;
        RECT 131.250 194.660 131.390 196.525 ;
        RECT 131.190 194.340 131.450 194.660 ;
        RECT 130.730 189.580 130.990 189.900 ;
        RECT 130.330 189.220 130.930 189.300 ;
        RECT 130.330 189.160 130.990 189.220 ;
        RECT 130.730 188.900 130.990 189.160 ;
        RECT 130.270 188.220 130.530 188.540 ;
        RECT 130.330 188.055 130.470 188.220 ;
        RECT 130.260 187.685 130.540 188.055 ;
        RECT 131.250 184.460 131.390 194.340 ;
        RECT 131.710 193.495 131.850 207.350 ;
        RECT 132.170 201.140 132.310 207.600 ;
        RECT 133.090 205.540 133.230 208.200 ;
        RECT 133.480 208.085 133.760 208.455 ;
        RECT 133.550 207.240 133.690 208.085 ;
        RECT 133.490 206.920 133.750 207.240 ;
        RECT 133.030 205.220 133.290 205.540 ;
        RECT 133.090 202.900 133.230 205.220 ;
        RECT 133.550 203.500 133.690 206.920 ;
        RECT 133.490 203.180 133.750 203.500 ;
        RECT 133.090 202.760 133.690 202.900 ;
        RECT 132.170 201.000 132.770 201.140 ;
        RECT 132.630 200.100 132.770 201.000 ;
        RECT 132.110 199.780 132.370 200.100 ;
        RECT 132.570 199.780 132.830 200.100 ;
        RECT 133.030 199.780 133.290 200.100 ;
        RECT 132.170 196.360 132.310 199.780 ;
        RECT 133.090 199.615 133.230 199.780 ;
        RECT 133.020 199.245 133.300 199.615 ;
        RECT 132.570 198.760 132.830 199.080 ;
        RECT 132.110 196.040 132.370 196.360 ;
        RECT 131.640 193.125 131.920 193.495 ;
        RECT 131.190 184.140 131.450 184.460 ;
        RECT 131.710 178.000 131.850 193.125 ;
        RECT 132.100 189.725 132.380 190.095 ;
        RECT 132.170 189.560 132.310 189.725 ;
        RECT 132.110 189.240 132.370 189.560 ;
        RECT 132.100 182.500 132.380 182.615 ;
        RECT 132.630 182.500 132.770 198.760 ;
        RECT 133.030 197.060 133.290 197.380 ;
        RECT 133.090 195.340 133.230 197.060 ;
        RECT 133.030 195.020 133.290 195.340 ;
        RECT 133.090 186.160 133.230 195.020 ;
        RECT 133.550 191.260 133.690 202.760 ;
        RECT 133.490 190.940 133.750 191.260 ;
        RECT 134.010 189.980 134.150 210.320 ;
        RECT 134.930 208.455 135.070 212.360 ;
        RECT 135.850 211.660 135.990 212.360 ;
        RECT 135.790 211.340 136.050 211.660 ;
        RECT 135.320 208.765 135.600 209.135 ;
        RECT 134.860 208.085 135.140 208.455 ;
        RECT 134.410 207.600 134.670 207.920 ;
        RECT 134.470 206.220 134.610 207.600 ;
        RECT 134.410 205.900 134.670 206.220 ;
        RECT 134.870 204.200 135.130 204.520 ;
        RECT 134.930 202.140 135.070 204.200 ;
        RECT 134.870 201.820 135.130 202.140 ;
        RECT 135.390 200.780 135.530 208.765 ;
        RECT 135.790 207.600 136.050 207.920 ;
        RECT 135.330 200.460 135.590 200.780 ;
        RECT 134.870 198.760 135.130 199.080 ;
        RECT 134.930 197.380 135.070 198.760 ;
        RECT 135.850 198.060 135.990 207.600 ;
        RECT 136.310 202.820 136.450 217.800 ;
        RECT 136.710 216.440 136.970 216.760 ;
        RECT 136.770 215.400 136.910 216.440 ;
        RECT 136.710 215.080 136.970 215.400 ;
        RECT 137.170 210.660 137.430 210.980 ;
        RECT 136.700 210.125 136.980 210.495 ;
        RECT 136.770 208.260 136.910 210.125 ;
        RECT 137.230 208.600 137.370 210.660 ;
        RECT 137.170 208.280 137.430 208.600 ;
        RECT 136.710 207.940 136.970 208.260 ;
        RECT 136.250 202.500 136.510 202.820 ;
        RECT 136.710 202.500 136.970 202.820 ;
        RECT 135.790 197.740 136.050 198.060 ;
        RECT 134.870 197.060 135.130 197.380 ;
        RECT 134.410 196.720 134.670 197.040 ;
        RECT 135.330 196.720 135.590 197.040 ;
        RECT 134.470 194.660 134.610 196.720 ;
        RECT 134.870 196.380 135.130 196.700 ;
        RECT 134.930 196.215 135.070 196.380 ;
        RECT 135.390 196.360 135.530 196.720 ;
        RECT 135.790 196.380 136.050 196.700 ;
        RECT 136.250 196.380 136.510 196.700 ;
        RECT 134.860 195.845 135.140 196.215 ;
        RECT 135.330 196.040 135.590 196.360 ;
        RECT 135.850 195.340 135.990 196.380 ;
        RECT 134.870 195.020 135.130 195.340 ;
        RECT 135.790 195.020 136.050 195.340 ;
        RECT 134.930 194.660 135.070 195.020 ;
        RECT 136.310 194.660 136.450 196.380 ;
        RECT 134.410 194.340 134.670 194.660 ;
        RECT 134.870 194.340 135.130 194.660 ;
        RECT 136.250 194.570 136.510 194.660 ;
        RECT 135.390 194.430 136.510 194.570 ;
        RECT 134.870 193.660 135.130 193.980 ;
        RECT 133.550 189.840 134.150 189.980 ;
        RECT 133.030 185.840 133.290 186.160 ;
        RECT 133.090 183.780 133.230 185.840 ;
        RECT 133.550 184.460 133.690 189.840 ;
        RECT 133.950 188.900 134.210 189.220 ;
        RECT 134.010 186.070 134.150 188.900 ;
        RECT 134.930 186.160 135.070 193.660 ;
        RECT 135.390 192.815 135.530 194.430 ;
        RECT 136.250 194.340 136.510 194.430 ;
        RECT 135.790 193.660 136.050 193.980 ;
        RECT 135.320 192.445 135.600 192.815 ;
        RECT 135.330 191.960 135.590 192.280 ;
        RECT 134.410 186.070 134.670 186.160 ;
        RECT 134.010 185.930 134.670 186.070 ;
        RECT 134.410 185.840 134.670 185.930 ;
        RECT 134.870 185.840 135.130 186.160 ;
        RECT 133.950 185.160 134.210 185.480 ;
        RECT 134.410 185.160 134.670 185.480 ;
        RECT 133.490 184.140 133.750 184.460 ;
        RECT 134.010 183.780 134.150 185.160 ;
        RECT 133.030 183.460 133.290 183.780 ;
        RECT 133.950 183.460 134.210 183.780 ;
        RECT 134.470 182.760 134.610 185.160 ;
        RECT 132.100 182.360 132.770 182.500 ;
        RECT 134.410 182.440 134.670 182.760 ;
        RECT 134.930 182.670 135.070 185.840 ;
        RECT 135.390 183.180 135.530 191.960 ;
        RECT 135.850 186.500 135.990 193.660 ;
        RECT 135.790 186.180 136.050 186.500 ;
        RECT 135.780 184.965 136.060 185.335 ;
        RECT 135.850 184.460 135.990 184.965 ;
        RECT 135.790 184.140 136.050 184.460 ;
        RECT 135.390 183.040 135.990 183.180 ;
        RECT 134.930 182.530 135.530 182.670 ;
        RECT 132.100 182.245 132.380 182.360 ;
        RECT 134.860 181.565 135.140 181.935 ;
        RECT 132.560 180.885 132.840 181.255 ;
        RECT 132.630 180.380 132.770 180.885 ;
        RECT 132.570 180.060 132.830 180.380 ;
        RECT 133.490 180.060 133.750 180.380 ;
        RECT 133.550 178.340 133.690 180.060 ;
        RECT 132.110 178.020 132.370 178.340 ;
        RECT 133.490 178.020 133.750 178.340 ;
        RECT 131.650 177.680 131.910 178.000 ;
        RECT 131.650 174.620 131.910 174.940 ;
        RECT 131.710 173.095 131.850 174.620 ;
        RECT 131.640 172.725 131.920 173.095 ;
        RECT 132.170 172.560 132.310 178.020 ;
        RECT 134.930 178.000 135.070 181.565 ;
        RECT 135.390 180.040 135.530 182.530 ;
        RECT 135.330 179.720 135.590 180.040 ;
        RECT 134.870 177.680 135.130 178.000 ;
        RECT 135.330 177.855 135.590 178.000 ;
        RECT 134.410 174.620 134.670 174.940 ;
        RECT 134.470 172.560 134.610 174.620 ;
        RECT 134.930 174.600 135.070 177.680 ;
        RECT 135.320 177.485 135.600 177.855 ;
        RECT 135.330 174.960 135.590 175.280 ;
        RECT 134.870 174.280 135.130 174.600 ;
        RECT 132.110 172.240 132.370 172.560 ;
        RECT 134.410 172.240 134.670 172.560 ;
        RECT 133.020 170.685 133.300 171.055 ;
        RECT 134.470 170.860 134.610 172.240 ;
        RECT 134.870 171.560 135.130 171.880 ;
        RECT 134.930 170.860 135.070 171.560 ;
        RECT 131.650 169.180 131.910 169.500 ;
        RECT 131.710 167.800 131.850 169.180 ;
        RECT 133.090 167.800 133.230 170.685 ;
        RECT 134.410 170.540 134.670 170.860 ;
        RECT 134.870 170.540 135.130 170.860 ;
        RECT 133.950 169.520 134.210 169.840 ;
        RECT 131.650 167.480 131.910 167.800 ;
        RECT 133.030 167.480 133.290 167.800 ;
        RECT 133.030 166.800 133.290 167.120 ;
        RECT 132.570 164.760 132.830 165.080 ;
        RECT 132.630 164.255 132.770 164.760 ;
        RECT 130.270 163.740 130.530 164.060 ;
        RECT 132.560 163.885 132.840 164.255 ;
        RECT 130.330 162.700 130.470 163.740 ;
        RECT 132.630 162.700 132.770 163.885 ;
        RECT 130.270 162.380 130.530 162.700 ;
        RECT 132.570 162.380 132.830 162.700 ;
        RECT 133.090 161.680 133.230 166.800 ;
        RECT 134.010 166.780 134.150 169.520 ;
        RECT 134.470 167.460 134.610 170.540 ;
        RECT 135.390 167.460 135.530 174.960 ;
        RECT 134.410 167.140 134.670 167.460 ;
        RECT 135.330 167.140 135.590 167.460 ;
        RECT 133.950 166.460 134.210 166.780 ;
        RECT 134.010 164.740 134.150 166.460 ;
        RECT 133.950 164.420 134.210 164.740 ;
        RECT 130.270 161.360 130.530 161.680 ;
        RECT 133.030 161.360 133.290 161.680 ;
        RECT 133.490 161.360 133.750 161.680 ;
        RECT 130.330 160.855 130.470 161.360 ;
        RECT 130.260 160.485 130.540 160.855 ;
        RECT 133.550 158.960 133.690 161.360 ;
        RECT 131.180 158.445 131.460 158.815 ;
        RECT 133.490 158.640 133.750 158.960 ;
        RECT 130.270 157.960 130.530 158.280 ;
        RECT 129.810 156.940 130.070 157.260 ;
        RECT 129.350 156.260 129.610 156.580 ;
        RECT 128.890 153.200 129.150 153.520 ;
        RECT 128.950 151.820 129.090 153.200 ;
        RECT 128.430 151.500 128.690 151.820 ;
        RECT 128.890 151.500 129.150 151.820 ;
        RECT 129.870 151.335 130.010 156.940 ;
        RECT 129.350 150.820 129.610 151.140 ;
        RECT 129.800 150.965 130.080 151.335 ;
        RECT 127.510 150.480 127.770 150.800 ;
        RECT 129.410 150.655 129.550 150.820 ;
        RECT 124.750 147.850 125.870 147.990 ;
        RECT 126.190 148.360 127.250 148.500 ;
        RECT 127.570 148.420 127.710 150.480 ;
        RECT 129.340 150.285 129.620 150.655 ;
        RECT 128.890 148.440 129.150 148.760 ;
        RECT 126.190 147.935 126.330 148.360 ;
        RECT 127.510 148.100 127.770 148.420 ;
        RECT 124.750 147.760 125.010 147.850 ;
        RECT 122.450 145.380 122.710 145.700 ;
        RECT 121.990 142.320 122.250 142.640 ;
        RECT 122.050 141.815 122.190 142.320 ;
        RECT 121.980 141.445 122.260 141.815 ;
        RECT 121.060 140.765 121.340 141.135 ;
        RECT 122.510 140.940 122.650 145.380 ;
        RECT 123.430 144.680 123.570 147.760 ;
        RECT 124.810 146.040 124.950 147.760 ;
        RECT 126.120 147.565 126.400 147.935 ;
        RECT 126.590 147.420 126.850 147.740 ;
        RECT 126.130 147.080 126.390 147.400 ;
        RECT 124.750 145.720 125.010 146.040 ;
        RECT 125.670 145.040 125.930 145.360 ;
        RECT 123.830 144.700 124.090 145.020 ;
        RECT 123.370 144.360 123.630 144.680 ;
        RECT 123.890 142.980 124.030 144.700 ;
        RECT 125.730 143.320 125.870 145.040 ;
        RECT 125.670 143.000 125.930 143.320 ;
        RECT 123.830 142.660 124.090 142.980 ;
        RECT 125.730 142.640 125.870 143.000 ;
        RECT 123.370 142.320 123.630 142.640 ;
        RECT 124.750 142.495 125.010 142.640 ;
        RECT 120.610 140.280 120.870 140.600 ;
        RECT 116.010 139.600 116.270 139.920 ;
        RECT 116.470 139.600 116.730 139.920 ;
        RECT 115.550 138.920 115.810 139.240 ;
        RECT 115.090 137.560 115.350 137.880 ;
        RECT 111.930 135.695 112.070 136.880 ;
        RECT 112.390 136.800 112.990 136.940 ;
        RECT 114.170 136.880 114.430 137.200 ;
        RECT 114.630 136.880 114.890 137.200 ;
        RECT 112.330 136.200 112.590 136.520 ;
        RECT 111.860 135.325 112.140 135.695 ;
        RECT 111.410 134.500 111.670 134.820 ;
        RECT 112.390 132.440 112.530 136.200 ;
        RECT 112.850 135.160 112.990 136.800 ;
        RECT 112.790 134.840 113.050 135.160 ;
        RECT 114.230 134.820 114.370 136.880 ;
        RECT 115.150 135.500 115.290 137.560 ;
        RECT 115.610 135.500 115.750 138.920 ;
        RECT 116.070 136.860 116.210 139.600 ;
        RECT 116.530 137.540 116.670 139.600 ;
        RECT 116.470 137.220 116.730 137.540 ;
        RECT 116.990 136.860 117.130 140.200 ;
        RECT 117.390 139.940 117.650 140.260 ;
        RECT 117.850 139.940 118.110 140.260 ;
        RECT 117.850 138.920 118.110 139.240 ;
        RECT 116.010 136.540 116.270 136.860 ;
        RECT 116.930 136.540 117.190 136.860 ;
        RECT 117.910 135.500 118.050 138.920 ;
        RECT 121.130 138.220 121.270 140.765 ;
        RECT 122.450 140.620 122.710 140.940 ;
        RECT 121.530 139.775 121.790 139.920 ;
        RECT 121.520 139.405 121.800 139.775 ;
        RECT 122.910 139.600 123.170 139.920 ;
        RECT 122.450 138.920 122.710 139.240 ;
        RECT 121.070 137.900 121.330 138.220 ;
        RECT 121.990 137.560 122.250 137.880 ;
        RECT 119.680 136.940 119.960 137.055 ;
        RECT 119.290 136.860 119.960 136.940 ;
        RECT 122.050 136.860 122.190 137.560 ;
        RECT 119.230 136.800 119.960 136.860 ;
        RECT 119.230 136.540 119.490 136.800 ;
        RECT 119.680 136.685 119.960 136.800 ;
        RECT 121.990 136.540 122.250 136.860 ;
        RECT 119.690 136.430 119.950 136.520 ;
        RECT 119.690 136.290 121.270 136.430 ;
        RECT 119.690 136.200 119.950 136.290 ;
        RECT 118.590 135.665 120.130 136.035 ;
        RECT 121.130 135.500 121.270 136.290 ;
        RECT 115.090 135.180 115.350 135.500 ;
        RECT 115.550 135.180 115.810 135.500 ;
        RECT 117.850 135.180 118.110 135.500 ;
        RECT 121.070 135.180 121.330 135.500 ;
        RECT 121.990 135.180 122.250 135.500 ;
        RECT 114.170 134.500 114.430 134.820 ;
        RECT 114.630 134.500 114.890 134.820 ;
        RECT 117.380 134.645 117.660 135.015 ;
        RECT 114.690 132.780 114.830 134.500 ;
        RECT 116.010 133.820 116.270 134.140 ;
        RECT 114.630 132.460 114.890 132.780 ;
        RECT 112.330 132.120 112.590 132.440 ;
        RECT 107.270 130.760 107.530 131.080 ;
        RECT 107.730 130.760 107.990 131.080 ;
        RECT 107.330 130.060 107.470 130.760 ;
        RECT 107.270 129.740 107.530 130.060 ;
        RECT 107.270 129.290 107.530 129.380 ;
        RECT 104.970 129.060 105.230 129.205 ;
        RECT 106.870 129.150 107.530 129.290 ;
        RECT 107.270 129.060 107.530 129.150 ;
        RECT 104.510 128.720 104.770 129.040 ;
        RECT 104.050 128.040 104.310 128.360 ;
        RECT 98.070 126.340 98.330 126.660 ;
        RECT 98.530 126.340 98.790 126.660 ;
        RECT 99.050 126.600 101.490 126.740 ;
        RECT 103.590 126.680 103.850 127.000 ;
        RECT 98.130 123.940 98.270 126.340 ;
        RECT 99.050 126.320 99.190 126.600 ;
        RECT 101.350 126.320 101.490 126.600 ;
        RECT 98.990 126.000 99.250 126.320 ;
        RECT 99.910 126.000 100.170 126.320 ;
        RECT 99.970 125.640 100.110 126.000 ;
        RECT 100.360 125.805 100.640 126.175 ;
        RECT 101.290 126.000 101.550 126.320 ;
        RECT 100.430 125.640 100.570 125.805 ;
        RECT 99.910 125.320 100.170 125.640 ;
        RECT 100.370 125.320 100.630 125.640 ;
        RECT 99.970 123.940 100.110 125.320 ;
        RECT 104.110 123.940 104.250 128.040 ;
        RECT 104.570 125.240 104.710 128.720 ;
        RECT 107.330 128.215 107.470 129.060 ;
        RECT 107.260 127.845 107.540 128.215 ;
        RECT 107.330 126.060 107.470 127.845 ;
        RECT 107.790 126.320 107.930 130.760 ;
        RECT 106.410 125.980 107.470 126.060 ;
        RECT 107.730 126.000 107.990 126.320 ;
        RECT 108.250 126.060 108.390 131.360 ;
        RECT 109.560 131.360 110.230 131.500 ;
        RECT 109.560 131.245 109.840 131.360 ;
        RECT 109.110 130.760 109.370 131.080 ;
        RECT 109.170 130.060 109.310 130.760 ;
        RECT 110.090 130.060 110.230 131.360 ;
        RECT 110.550 131.360 111.150 131.500 ;
        RECT 108.650 129.740 108.910 130.060 ;
        RECT 109.110 129.740 109.370 130.060 ;
        RECT 110.030 129.740 110.290 130.060 ;
        RECT 108.710 126.855 108.850 129.740 ;
        RECT 109.570 129.060 109.830 129.380 ;
        RECT 109.110 128.720 109.370 129.040 ;
        RECT 109.630 128.780 109.770 129.060 ;
        RECT 109.170 127.000 109.310 128.720 ;
        RECT 109.630 128.700 110.230 128.780 ;
        RECT 109.630 128.640 110.290 128.700 ;
        RECT 110.030 128.380 110.290 128.640 ;
        RECT 110.550 127.340 110.690 131.360 ;
        RECT 111.410 130.760 111.670 131.080 ;
        RECT 110.490 127.020 110.750 127.340 ;
        RECT 108.640 126.485 108.920 126.855 ;
        RECT 109.110 126.680 109.370 127.000 ;
        RECT 108.650 126.340 108.910 126.485 ;
        RECT 106.350 125.920 107.470 125.980 ;
        RECT 108.250 125.920 108.850 126.060 ;
        RECT 106.350 125.660 106.610 125.920 ;
        RECT 107.270 125.380 107.530 125.640 ;
        RECT 107.270 125.320 108.390 125.380 ;
        RECT 107.330 125.240 108.390 125.320 ;
        RECT 104.570 125.100 105.170 125.240 ;
        RECT 104.510 123.960 104.770 124.280 ;
        RECT 95.310 123.620 95.570 123.940 ;
        RECT 96.230 123.620 96.490 123.940 ;
        RECT 96.690 123.620 96.950 123.940 ;
        RECT 97.150 123.620 97.410 123.940 ;
        RECT 98.070 123.620 98.330 123.940 ;
        RECT 99.910 123.620 100.170 123.940 ;
        RECT 104.050 123.620 104.310 123.940 ;
        RECT 94.850 123.280 95.110 123.600 ;
        RECT 94.850 122.600 95.110 122.920 ;
        RECT 90.710 121.580 90.970 121.900 ;
        RECT 94.390 121.580 94.650 121.900 ;
        RECT 87.490 121.240 87.750 121.560 ;
        RECT 82.890 120.560 83.150 120.880 ;
        RECT 94.910 120.200 95.050 122.600 ;
        RECT 95.310 120.900 95.570 121.220 ;
        RECT 78.750 119.880 79.010 120.200 ;
        RECT 94.850 119.880 95.110 120.200 ;
        RECT 79.720 119.345 81.260 119.715 ;
        RECT 70.930 118.520 71.190 118.840 ;
        RECT 95.370 118.160 95.510 120.900 ;
        RECT 95.770 119.880 96.030 120.200 ;
        RECT 95.830 118.500 95.970 119.880 ;
        RECT 96.290 119.180 96.430 123.620 ;
        RECT 98.130 123.260 99.190 123.340 ;
        RECT 101.750 123.280 102.010 123.600 ;
        RECT 98.130 123.200 99.250 123.260 ;
        RECT 96.690 121.580 96.950 121.900 ;
        RECT 96.750 119.180 96.890 121.580 ;
        RECT 98.130 121.560 98.270 123.200 ;
        RECT 98.990 122.940 99.250 123.200 ;
        RECT 99.155 122.065 100.695 122.435 ;
        RECT 98.070 121.240 98.330 121.560 ;
        RECT 101.810 120.880 101.950 123.280 ;
        RECT 104.570 121.900 104.710 123.960 ;
        RECT 105.030 123.940 105.170 125.100 ;
        RECT 106.810 124.300 107.070 124.620 ;
        RECT 104.970 123.620 105.230 123.940 ;
        RECT 106.350 123.620 106.610 123.940 ;
        RECT 106.410 121.900 106.550 123.620 ;
        RECT 104.510 121.580 104.770 121.900 ;
        RECT 106.350 121.580 106.610 121.900 ;
        RECT 98.530 120.560 98.790 120.880 ;
        RECT 101.750 120.560 102.010 120.880 ;
        RECT 104.050 120.560 104.310 120.880 ;
        RECT 96.230 118.860 96.490 119.180 ;
        RECT 96.690 118.860 96.950 119.180 ;
        RECT 98.590 118.500 98.730 120.560 ;
        RECT 102.210 120.220 102.470 120.540 ;
        RECT 102.270 119.180 102.410 120.220 ;
        RECT 104.110 120.200 104.250 120.560 ;
        RECT 104.050 119.880 104.310 120.200 ;
        RECT 106.870 119.180 107.010 124.300 ;
        RECT 107.730 124.190 107.990 124.280 ;
        RECT 108.250 124.190 108.390 125.240 ;
        RECT 107.730 124.050 108.390 124.190 ;
        RECT 107.730 123.960 107.990 124.050 ;
        RECT 107.270 123.280 107.530 123.600 ;
        RECT 107.330 121.300 107.470 123.280 ;
        RECT 107.330 121.160 107.930 121.300 ;
        RECT 107.790 120.880 107.930 121.160 ;
        RECT 107.730 120.560 107.990 120.880 ;
        RECT 108.710 120.540 108.850 125.920 ;
        RECT 110.490 125.660 110.750 125.980 ;
        RECT 110.030 125.320 110.290 125.640 ;
        RECT 109.570 124.300 109.830 124.620 ;
        RECT 109.110 122.600 109.370 122.920 ;
        RECT 108.650 120.220 108.910 120.540 ;
        RECT 102.210 118.860 102.470 119.180 ;
        RECT 106.810 118.860 107.070 119.180 ;
        RECT 109.170 118.840 109.310 122.600 ;
        RECT 109.630 121.220 109.770 124.300 ;
        RECT 110.090 123.940 110.230 125.320 ;
        RECT 110.030 123.620 110.290 123.940 ;
        RECT 110.550 123.260 110.690 125.660 ;
        RECT 111.470 125.240 111.610 130.760 ;
        RECT 114.690 129.380 114.830 132.460 ;
        RECT 116.070 132.440 116.210 133.820 ;
        RECT 116.930 133.480 117.190 133.800 ;
        RECT 116.010 132.120 116.270 132.440 ;
        RECT 115.080 131.245 115.360 131.615 ;
        RECT 115.150 131.080 115.290 131.245 ;
        RECT 115.090 130.760 115.350 131.080 ;
        RECT 116.070 130.060 116.210 132.120 ;
        RECT 116.470 131.615 116.730 131.760 ;
        RECT 116.460 131.245 116.740 131.615 ;
        RECT 116.010 129.740 116.270 130.060 ;
        RECT 114.630 129.060 114.890 129.380 ;
        RECT 111.870 125.660 112.130 125.980 ;
        RECT 111.010 125.100 111.610 125.240 ;
        RECT 111.010 123.940 111.150 125.100 ;
        RECT 111.930 124.620 112.070 125.660 ;
        RECT 114.690 125.240 114.830 129.060 ;
        RECT 116.470 128.720 116.730 129.040 ;
        RECT 115.550 128.040 115.810 128.360 ;
        RECT 115.610 127.340 115.750 128.040 ;
        RECT 116.530 127.340 116.670 128.720 ;
        RECT 115.090 127.020 115.350 127.340 ;
        RECT 115.550 127.020 115.810 127.340 ;
        RECT 116.470 127.020 116.730 127.340 ;
        RECT 115.150 126.060 115.290 127.020 ;
        RECT 116.990 126.320 117.130 133.480 ;
        RECT 117.450 132.440 117.590 134.645 ;
        RECT 119.230 133.480 119.490 133.800 ;
        RECT 117.390 132.120 117.650 132.440 ;
        RECT 119.290 132.010 119.430 133.480 ;
        RECT 120.610 132.460 120.870 132.780 ;
        RECT 118.830 131.870 119.430 132.010 ;
        RECT 118.830 131.080 118.970 131.870 ;
        RECT 117.850 130.760 118.110 131.080 ;
        RECT 118.770 130.760 119.030 131.080 ;
        RECT 117.910 129.460 118.050 130.760 ;
        RECT 118.590 130.225 120.130 130.595 ;
        RECT 119.230 129.740 119.490 130.060 ;
        RECT 117.910 129.320 118.970 129.460 ;
        RECT 118.310 128.950 118.570 129.040 ;
        RECT 117.450 128.810 118.570 128.950 ;
        RECT 116.010 126.060 116.270 126.320 ;
        RECT 115.150 126.000 116.270 126.060 ;
        RECT 116.930 126.000 117.190 126.320 ;
        RECT 115.150 125.920 116.210 126.000 ;
        RECT 114.690 125.100 117.130 125.240 ;
        RECT 116.990 124.620 117.130 125.100 ;
        RECT 111.870 124.300 112.130 124.620 ;
        RECT 116.930 124.300 117.190 124.620 ;
        RECT 110.950 123.620 111.210 123.940 ;
        RECT 117.450 123.260 117.590 128.810 ;
        RECT 118.310 128.720 118.570 128.810 ;
        RECT 117.850 128.040 118.110 128.360 ;
        RECT 117.910 123.940 118.050 128.040 ;
        RECT 118.830 127.000 118.970 129.320 ;
        RECT 118.770 126.680 119.030 127.000 ;
        RECT 119.290 126.320 119.430 129.740 ;
        RECT 120.150 129.060 120.410 129.380 ;
        RECT 120.210 128.895 120.350 129.060 ;
        RECT 120.140 128.525 120.420 128.895 ;
        RECT 120.670 127.340 120.810 132.460 ;
        RECT 122.050 132.295 122.190 135.180 ;
        RECT 122.510 134.820 122.650 138.920 ;
        RECT 122.450 134.500 122.710 134.820 ;
        RECT 121.980 131.925 122.260 132.295 ;
        RECT 122.050 129.720 122.190 131.925 ;
        RECT 121.990 129.400 122.250 129.720 ;
        RECT 122.970 129.630 123.110 139.600 ;
        RECT 123.430 132.440 123.570 142.320 ;
        RECT 124.740 142.125 125.020 142.495 ;
        RECT 125.670 142.320 125.930 142.640 ;
        RECT 125.670 141.640 125.930 141.960 ;
        RECT 125.730 140.940 125.870 141.640 ;
        RECT 126.190 140.940 126.330 147.080 ;
        RECT 126.650 142.640 126.790 147.420 ;
        RECT 127.050 145.720 127.310 146.040 ;
        RECT 127.110 144.535 127.250 145.720 ;
        RECT 127.570 145.360 127.710 148.100 ;
        RECT 127.970 147.080 128.230 147.400 ;
        RECT 128.430 147.080 128.690 147.400 ;
        RECT 128.030 146.380 128.170 147.080 ;
        RECT 127.970 146.060 128.230 146.380 ;
        RECT 127.510 145.040 127.770 145.360 ;
        RECT 127.960 144.845 128.240 145.215 ;
        RECT 127.040 144.165 127.320 144.535 ;
        RECT 127.500 142.805 127.780 143.175 ;
        RECT 126.590 142.550 126.850 142.640 ;
        RECT 126.590 142.410 127.250 142.550 ;
        RECT 126.590 142.320 126.850 142.410 ;
        RECT 126.590 141.640 126.850 141.960 ;
        RECT 125.670 140.620 125.930 140.940 ;
        RECT 126.130 140.620 126.390 140.940 ;
        RECT 124.280 140.085 124.560 140.455 ;
        RECT 124.290 139.940 124.550 140.085 ;
        RECT 124.750 139.600 125.010 139.920 ;
        RECT 124.810 138.220 124.950 139.600 ;
        RECT 125.210 138.920 125.470 139.240 ;
        RECT 124.750 137.900 125.010 138.220 ;
        RECT 123.830 137.560 124.090 137.880 ;
        RECT 123.890 134.335 124.030 137.560 ;
        RECT 123.820 134.220 124.100 134.335 ;
        RECT 123.820 134.080 124.950 134.220 ;
        RECT 123.820 133.965 124.100 134.080 ;
        RECT 123.370 132.120 123.630 132.440 ;
        RECT 124.290 131.440 124.550 131.760 ;
        RECT 123.830 130.760 124.090 131.080 ;
        RECT 122.510 129.490 123.110 129.630 ;
        RECT 122.510 128.360 122.650 129.490 ;
        RECT 123.370 129.290 123.630 129.380 ;
        RECT 122.970 129.150 123.630 129.290 ;
        RECT 122.450 128.040 122.710 128.360 ;
        RECT 120.610 127.020 120.870 127.340 ;
        RECT 121.070 126.570 121.330 126.660 ;
        RECT 119.750 126.430 122.190 126.570 ;
        RECT 119.230 126.000 119.490 126.320 ;
        RECT 119.750 125.980 119.890 126.430 ;
        RECT 121.070 126.340 121.330 126.430 ;
        RECT 119.690 125.660 119.950 125.980 ;
        RECT 121.070 125.660 121.330 125.980 ;
        RECT 120.610 125.320 120.870 125.640 ;
        RECT 118.590 124.785 120.130 125.155 ;
        RECT 120.670 124.530 120.810 125.320 ;
        RECT 120.210 124.390 120.810 124.530 ;
        RECT 117.850 123.620 118.110 123.940 ;
        RECT 120.210 123.600 120.350 124.390 ;
        RECT 120.150 123.280 120.410 123.600 ;
        RECT 121.130 123.260 121.270 125.660 ;
        RECT 121.530 123.620 121.790 123.940 ;
        RECT 110.490 122.940 110.750 123.260 ;
        RECT 117.390 122.940 117.650 123.260 ;
        RECT 121.070 122.940 121.330 123.260 ;
        RECT 111.410 122.600 111.670 122.920 ;
        RECT 111.470 121.900 111.610 122.600 ;
        RECT 111.410 121.580 111.670 121.900 ;
        RECT 117.450 121.560 117.590 122.940 ;
        RECT 121.590 122.920 121.730 123.620 ;
        RECT 118.770 122.600 119.030 122.920 ;
        RECT 121.530 122.600 121.790 122.920 ;
        RECT 118.830 121.900 118.970 122.600 ;
        RECT 122.050 121.900 122.190 126.430 ;
        RECT 122.970 123.940 123.110 129.150 ;
        RECT 123.370 129.060 123.630 129.150 ;
        RECT 123.360 126.485 123.640 126.855 ;
        RECT 123.370 126.340 123.630 126.485 ;
        RECT 123.370 125.660 123.630 125.980 ;
        RECT 122.910 123.620 123.170 123.940 ;
        RECT 122.970 121.900 123.110 123.620 ;
        RECT 123.430 123.510 123.570 125.660 ;
        RECT 123.890 124.280 124.030 130.760 ;
        RECT 124.350 129.720 124.490 131.440 ;
        RECT 124.290 129.400 124.550 129.720 ;
        RECT 124.810 128.780 124.950 134.080 ;
        RECT 125.270 131.615 125.410 138.920 ;
        RECT 125.730 137.620 125.870 140.620 ;
        RECT 126.190 140.260 126.330 140.620 ;
        RECT 126.130 139.940 126.390 140.260 ;
        RECT 126.120 137.620 126.400 137.735 ;
        RECT 125.730 137.480 126.400 137.620 ;
        RECT 125.730 135.500 125.870 137.480 ;
        RECT 126.120 137.365 126.400 137.480 ;
        RECT 125.670 135.180 125.930 135.500 ;
        RECT 126.130 134.840 126.390 135.160 ;
        RECT 125.670 134.500 125.930 134.820 ;
        RECT 125.730 131.760 125.870 134.500 ;
        RECT 125.200 131.245 125.480 131.615 ;
        RECT 125.670 131.440 125.930 131.760 ;
        RECT 124.350 128.640 124.950 128.780 ;
        RECT 124.350 128.215 124.490 128.640 ;
        RECT 124.280 127.845 124.560 128.215 ;
        RECT 124.750 128.040 125.010 128.360 ;
        RECT 124.350 127.340 124.490 127.845 ;
        RECT 124.810 127.340 124.950 128.040 ;
        RECT 124.290 127.020 124.550 127.340 ;
        RECT 124.750 127.020 125.010 127.340 ;
        RECT 124.750 126.000 125.010 126.320 ;
        RECT 124.810 124.280 124.950 126.000 ;
        RECT 125.270 125.980 125.410 131.245 ;
        RECT 125.660 129.885 125.940 130.255 ;
        RECT 125.730 129.380 125.870 129.885 ;
        RECT 125.670 129.060 125.930 129.380 ;
        RECT 126.190 128.895 126.330 134.840 ;
        RECT 126.650 134.480 126.790 141.640 ;
        RECT 127.110 137.200 127.250 142.410 ;
        RECT 127.570 140.170 127.710 142.805 ;
        RECT 128.030 142.640 128.170 144.845 ;
        RECT 128.490 143.855 128.630 147.080 ;
        RECT 128.420 143.485 128.700 143.855 ;
        RECT 128.950 142.640 129.090 148.440 ;
        RECT 129.350 145.100 129.610 145.360 ;
        RECT 129.870 145.100 130.010 150.965 ;
        RECT 129.350 145.040 130.010 145.100 ;
        RECT 129.410 144.960 130.010 145.040 ;
        RECT 130.330 144.590 130.470 157.960 ;
        RECT 130.730 155.920 130.990 156.240 ;
        RECT 130.790 154.540 130.930 155.920 ;
        RECT 131.250 154.540 131.390 158.445 ;
        RECT 131.650 157.960 131.910 158.280 ;
        RECT 132.110 157.960 132.370 158.280 ;
        RECT 130.730 154.220 130.990 154.540 ;
        RECT 131.190 154.220 131.450 154.540 ;
        RECT 131.710 148.760 131.850 157.960 ;
        RECT 132.170 157.260 132.310 157.960 ;
        RECT 132.110 156.940 132.370 157.260 ;
        RECT 133.030 155.580 133.290 155.900 ;
        RECT 132.570 151.050 132.830 151.140 ;
        RECT 133.090 151.050 133.230 155.580 ;
        RECT 133.550 153.180 133.690 158.640 ;
        RECT 135.850 158.620 135.990 183.040 ;
        RECT 136.310 177.660 136.450 194.340 ;
        RECT 136.250 177.340 136.510 177.660 ;
        RECT 136.310 173.580 136.450 177.340 ;
        RECT 136.770 176.300 136.910 202.500 ;
        RECT 137.230 197.040 137.370 208.280 ;
        RECT 137.170 196.720 137.430 197.040 ;
        RECT 137.230 195.340 137.370 196.720 ;
        RECT 137.170 195.020 137.430 195.340 ;
        RECT 137.690 191.940 137.830 218.480 ;
        RECT 139.010 216.100 139.270 216.420 ;
        RECT 139.470 216.330 139.730 216.420 ;
        RECT 139.470 216.190 140.130 216.330 ;
        RECT 139.470 216.100 139.730 216.190 ;
        RECT 139.070 215.400 139.210 216.100 ;
        RECT 139.010 215.080 139.270 215.400 ;
        RECT 138.025 214.545 139.565 214.915 ;
        RECT 138.025 209.105 139.565 209.475 ;
        RECT 138.025 203.665 139.565 204.035 ;
        RECT 139.000 202.645 139.280 203.015 ;
        RECT 139.070 202.140 139.210 202.645 ;
        RECT 139.010 201.820 139.270 202.140 ;
        RECT 138.025 198.225 139.565 198.595 ;
        RECT 139.990 198.060 140.130 216.190 ;
        RECT 141.770 215.760 142.030 216.080 ;
        RECT 140.390 215.080 140.650 215.400 ;
        RECT 140.450 210.980 140.590 215.080 ;
        RECT 141.830 212.680 141.970 215.760 ;
        RECT 142.290 213.700 142.430 219.500 ;
        RECT 144.070 218.820 144.330 219.140 ;
        RECT 142.690 216.100 142.950 216.420 ;
        RECT 142.230 213.380 142.490 213.700 ;
        RECT 141.770 212.360 142.030 212.680 ;
        RECT 140.390 210.660 140.650 210.980 ;
        RECT 142.750 210.300 142.890 216.100 ;
        RECT 143.150 213.040 143.410 213.360 ;
        RECT 144.130 213.100 144.270 218.820 ;
        RECT 148.730 218.800 148.870 221.005 ;
        RECT 150.040 220.325 150.320 220.695 ;
        RECT 151.420 220.325 151.700 220.695 ;
        RECT 150.110 218.800 150.250 220.325 ;
        RECT 151.490 218.800 151.630 220.325 ;
        RECT 144.990 218.540 145.250 218.800 ;
        RECT 144.990 218.480 145.650 218.540 ;
        RECT 145.910 218.480 146.170 218.800 ;
        RECT 148.670 218.480 148.930 218.800 ;
        RECT 150.050 218.480 150.310 218.800 ;
        RECT 151.430 218.480 151.690 218.800 ;
        RECT 145.050 218.400 145.650 218.480 ;
        RECT 144.990 217.800 145.250 218.120 ;
        RECT 140.390 209.980 140.650 210.300 ;
        RECT 142.690 209.980 142.950 210.300 ;
        RECT 140.450 203.160 140.590 209.980 ;
        RECT 143.210 207.150 143.350 213.040 ;
        RECT 143.670 212.960 144.270 213.100 ;
        RECT 143.670 212.420 143.810 212.960 ;
        RECT 143.670 212.280 144.270 212.420 ;
        RECT 142.750 207.010 143.350 207.150 ;
        RECT 140.850 204.200 141.110 204.520 ;
        RECT 140.390 202.840 140.650 203.160 ;
        RECT 140.390 200.460 140.650 200.780 ;
        RECT 139.930 197.740 140.190 198.060 ;
        RECT 138.090 196.720 138.350 197.040 ;
        RECT 138.150 193.980 138.290 196.720 ;
        RECT 138.090 193.660 138.350 193.980 ;
        RECT 138.025 192.785 139.565 193.155 ;
        RECT 137.630 191.620 137.890 191.940 ;
        RECT 137.170 190.940 137.430 191.260 ;
        RECT 137.230 189.220 137.370 190.940 ;
        RECT 137.630 190.600 137.890 190.920 ;
        RECT 137.690 189.900 137.830 190.600 ;
        RECT 137.630 189.580 137.890 189.900 ;
        RECT 138.540 189.725 138.820 190.095 ;
        RECT 138.610 189.560 138.750 189.725 ;
        RECT 138.550 189.240 138.810 189.560 ;
        RECT 137.170 188.900 137.430 189.220 ;
        RECT 137.630 188.900 137.890 189.220 ;
        RECT 139.930 189.130 140.190 189.220 ;
        RECT 140.450 189.130 140.590 200.460 ;
        RECT 140.910 191.940 141.050 204.200 ;
        RECT 141.760 201.965 142.040 202.335 ;
        RECT 141.830 200.100 141.970 201.965 ;
        RECT 142.230 200.120 142.490 200.440 ;
        RECT 141.770 199.780 142.030 200.100 ;
        RECT 141.310 197.400 141.570 197.720 ;
        RECT 141.370 194.660 141.510 197.400 ;
        RECT 141.830 196.700 141.970 199.780 ;
        RECT 141.770 196.380 142.030 196.700 ;
        RECT 141.310 194.340 141.570 194.660 ;
        RECT 141.770 193.320 142.030 193.640 ;
        RECT 140.850 191.620 141.110 191.940 ;
        RECT 139.930 188.990 140.590 189.130 ;
        RECT 139.930 188.900 140.190 188.990 ;
        RECT 141.310 188.900 141.570 189.220 ;
        RECT 137.690 187.180 137.830 188.900 ;
        RECT 138.025 187.345 139.565 187.715 ;
        RECT 137.630 186.860 137.890 187.180 ;
        RECT 139.990 186.500 140.130 188.900 ;
        RECT 140.850 186.860 141.110 187.180 ;
        RECT 139.930 186.180 140.190 186.500 ;
        RECT 140.390 185.500 140.650 185.820 ;
        RECT 137.170 183.800 137.430 184.120 ;
        RECT 137.230 181.740 137.370 183.800 ;
        RECT 139.930 182.440 140.190 182.760 ;
        RECT 138.025 181.905 139.565 182.275 ;
        RECT 137.170 181.420 137.430 181.740 ;
        RECT 137.160 178.165 137.440 178.535 ;
        RECT 138.550 178.360 138.810 178.680 ;
        RECT 137.170 178.020 137.430 178.165 ;
        RECT 136.710 175.980 136.970 176.300 ;
        RECT 137.230 175.280 137.370 178.020 ;
        RECT 138.610 178.000 138.750 178.360 ;
        RECT 138.550 177.680 138.810 178.000 ;
        RECT 138.025 176.465 139.565 176.835 ;
        RECT 139.990 176.300 140.130 182.440 ;
        RECT 140.450 178.680 140.590 185.500 ;
        RECT 140.390 178.360 140.650 178.680 ;
        RECT 139.930 175.980 140.190 176.300 ;
        RECT 140.910 175.960 141.050 186.860 ;
        RECT 141.370 184.460 141.510 188.900 ;
        RECT 141.310 184.140 141.570 184.460 ;
        RECT 141.310 180.740 141.570 181.060 ;
        RECT 137.620 175.445 137.900 175.815 ;
        RECT 140.850 175.640 141.110 175.960 ;
        RECT 137.630 175.300 137.890 175.445 ;
        RECT 141.370 175.280 141.510 180.740 ;
        RECT 141.830 180.380 141.970 193.320 ;
        RECT 142.290 185.900 142.430 200.120 ;
        RECT 142.750 199.760 142.890 207.010 ;
        RECT 143.150 202.160 143.410 202.480 ;
        RECT 142.690 199.440 142.950 199.760 ;
        RECT 142.750 195.250 142.890 199.440 ;
        RECT 143.210 199.420 143.350 202.160 ;
        RECT 143.610 199.780 143.870 200.100 ;
        RECT 143.150 199.100 143.410 199.420 ;
        RECT 143.210 197.380 143.350 199.100 ;
        RECT 143.150 197.060 143.410 197.380 ;
        RECT 142.750 195.110 143.350 195.250 ;
        RECT 142.690 194.340 142.950 194.660 ;
        RECT 142.750 188.200 142.890 194.340 ;
        RECT 143.210 192.280 143.350 195.110 ;
        RECT 143.670 194.855 143.810 199.780 ;
        RECT 143.600 194.485 143.880 194.855 ;
        RECT 144.130 193.980 144.270 212.280 ;
        RECT 145.050 207.920 145.190 217.800 ;
        RECT 145.510 216.760 145.650 218.400 ;
        RECT 145.970 217.100 146.110 218.480 ;
        RECT 148.210 218.140 148.470 218.460 ;
        RECT 146.830 217.800 147.090 218.120 ;
        RECT 145.910 216.780 146.170 217.100 ;
        RECT 145.450 216.440 145.710 216.760 ;
        RECT 145.510 214.380 145.650 216.440 ;
        RECT 145.450 214.060 145.710 214.380 ;
        RECT 145.910 212.700 146.170 213.020 ;
        RECT 145.970 211.660 146.110 212.700 ;
        RECT 145.910 211.340 146.170 211.660 ;
        RECT 145.450 208.280 145.710 208.600 ;
        RECT 144.520 207.405 144.800 207.775 ;
        RECT 144.990 207.600 145.250 207.920 ;
        RECT 144.590 205.540 144.730 207.405 ;
        RECT 145.510 206.300 145.650 208.280 ;
        RECT 146.890 207.920 147.030 217.800 ;
        RECT 147.290 214.060 147.550 214.380 ;
        RECT 147.350 211.660 147.490 214.060 ;
        RECT 147.750 212.700 148.010 213.020 ;
        RECT 147.290 211.340 147.550 211.660 ;
        RECT 147.290 208.620 147.550 208.940 ;
        RECT 145.910 207.600 146.170 207.920 ;
        RECT 146.370 207.600 146.630 207.920 ;
        RECT 146.830 207.600 147.090 207.920 ;
        RECT 145.050 206.160 145.650 206.300 ;
        RECT 144.530 205.220 144.790 205.540 ;
        RECT 144.530 204.200 144.790 204.520 ;
        RECT 144.590 200.780 144.730 204.200 ;
        RECT 144.530 200.460 144.790 200.780 ;
        RECT 144.530 197.060 144.790 197.380 ;
        RECT 144.590 193.980 144.730 197.060 ;
        RECT 144.070 193.660 144.330 193.980 ;
        RECT 144.530 193.660 144.790 193.980 ;
        RECT 143.150 191.960 143.410 192.280 ;
        RECT 143.610 191.280 143.870 191.600 ;
        RECT 143.150 188.900 143.410 189.220 ;
        RECT 142.690 187.880 142.950 188.200 ;
        RECT 142.290 185.760 142.890 185.900 ;
        RECT 142.230 185.160 142.490 185.480 ;
        RECT 142.290 183.295 142.430 185.160 ;
        RECT 142.750 183.780 142.890 185.760 ;
        RECT 142.690 183.460 142.950 183.780 ;
        RECT 142.220 182.925 142.500 183.295 ;
        RECT 143.210 181.060 143.350 188.900 ;
        RECT 143.670 183.780 143.810 191.280 ;
        RECT 143.610 183.460 143.870 183.780 ;
        RECT 143.150 180.740 143.410 181.060 ;
        RECT 141.770 180.060 142.030 180.380 ;
        RECT 143.140 180.205 143.420 180.575 ;
        RECT 141.830 178.680 141.970 180.060 ;
        RECT 141.770 178.360 142.030 178.680 ;
        RECT 143.210 177.660 143.350 180.205 ;
        RECT 143.150 177.340 143.410 177.660 ;
        RECT 137.170 174.960 137.430 175.280 ;
        RECT 141.310 174.960 141.570 175.280 ;
        RECT 136.250 173.260 136.510 173.580 ;
        RECT 145.050 173.540 145.190 206.160 ;
        RECT 145.970 205.735 146.110 207.600 ;
        RECT 146.430 206.220 146.570 207.600 ;
        RECT 146.370 205.900 146.630 206.220 ;
        RECT 145.450 205.220 145.710 205.540 ;
        RECT 145.900 205.365 146.180 205.735 ;
        RECT 145.510 197.380 145.650 205.220 ;
        RECT 146.370 203.180 146.630 203.500 ;
        RECT 145.910 200.120 146.170 200.440 ;
        RECT 145.970 197.720 146.110 200.120 ;
        RECT 145.910 197.400 146.170 197.720 ;
        RECT 145.450 197.060 145.710 197.380 ;
        RECT 145.970 194.660 146.110 197.400 ;
        RECT 145.910 194.340 146.170 194.660 ;
        RECT 146.430 193.640 146.570 203.180 ;
        RECT 147.350 199.080 147.490 208.620 ;
        RECT 147.810 203.500 147.950 212.700 ;
        RECT 148.270 207.920 148.410 218.140 ;
        RECT 151.430 217.800 151.690 218.120 ;
        RECT 151.490 215.255 151.630 217.800 ;
        RECT 151.420 214.885 151.700 215.255 ;
        RECT 148.660 213.525 148.940 213.895 ;
        RECT 148.730 211.320 148.870 213.525 ;
        RECT 150.970 213.380 151.230 213.700 ;
        RECT 149.590 213.040 149.850 213.360 ;
        RECT 148.670 211.000 148.930 211.320 ;
        RECT 149.650 208.940 149.790 213.040 ;
        RECT 150.510 212.360 150.770 212.680 ;
        RECT 149.590 208.620 149.850 208.940 ;
        RECT 148.210 207.600 148.470 207.920 ;
        RECT 149.130 207.600 149.390 207.920 ;
        RECT 147.750 203.180 148.010 203.500 ;
        RECT 147.290 198.760 147.550 199.080 ;
        RECT 146.830 196.720 147.090 197.040 ;
        RECT 146.890 194.660 147.030 196.720 ;
        RECT 146.830 194.340 147.090 194.660 ;
        RECT 146.370 193.320 146.630 193.640 ;
        RECT 146.890 192.620 147.030 194.340 ;
        RECT 146.830 192.300 147.090 192.620 ;
        RECT 146.830 188.900 147.090 189.220 ;
        RECT 146.890 187.180 147.030 188.900 ;
        RECT 146.830 186.860 147.090 187.180 ;
        RECT 145.450 183.460 145.710 183.780 ;
        RECT 145.510 178.340 145.650 183.460 ;
        RECT 145.450 178.020 145.710 178.340 ;
        RECT 147.350 177.320 147.490 198.760 ;
        RECT 147.750 194.340 148.010 194.660 ;
        RECT 147.810 189.900 147.950 194.340 ;
        RECT 148.210 192.300 148.470 192.620 ;
        RECT 147.750 189.580 148.010 189.900 ;
        RECT 148.270 189.220 148.410 192.300 ;
        RECT 148.670 190.940 148.930 191.260 ;
        RECT 148.730 189.415 148.870 190.940 ;
        RECT 148.210 188.900 148.470 189.220 ;
        RECT 148.660 189.045 148.940 189.415 ;
        RECT 148.670 188.900 148.930 189.045 ;
        RECT 148.270 183.780 148.410 188.900 ;
        RECT 149.190 188.880 149.330 207.600 ;
        RECT 149.590 204.880 149.850 205.200 ;
        RECT 149.650 200.780 149.790 204.880 ;
        RECT 150.570 202.480 150.710 212.360 ;
        RECT 151.030 207.920 151.170 213.380 ;
        RECT 151.950 213.100 152.090 221.200 ;
        RECT 154.190 220.520 154.450 220.840 ;
        RECT 154.250 217.100 154.390 220.520 ;
        RECT 157.460 217.265 159.000 217.635 ;
        RECT 154.190 216.780 154.450 217.100 ;
        RECT 152.810 215.760 153.070 216.080 ;
        RECT 152.350 215.080 152.610 215.400 ;
        RECT 152.410 214.380 152.550 215.080 ;
        RECT 152.350 214.060 152.610 214.380 ;
        RECT 152.870 214.040 153.010 215.760 ;
        RECT 152.810 213.720 153.070 214.040 ;
        RECT 154.250 213.700 154.390 216.780 ;
        RECT 154.650 216.100 154.910 216.420 ;
        RECT 154.190 213.380 154.450 213.700 ;
        RECT 151.430 212.700 151.690 213.020 ;
        RECT 151.950 212.960 152.550 213.100 ;
        RECT 153.730 213.040 153.990 213.360 ;
        RECT 151.490 208.600 151.630 212.700 ;
        RECT 152.410 210.980 152.550 212.960 ;
        RECT 153.790 211.740 153.930 213.040 ;
        RECT 153.790 211.660 154.390 211.740 ;
        RECT 153.730 211.600 154.390 211.660 ;
        RECT 153.730 211.340 153.990 211.600 ;
        RECT 152.350 210.660 152.610 210.980 ;
        RECT 153.730 210.660 153.990 210.980 ;
        RECT 151.430 208.280 151.690 208.600 ;
        RECT 150.970 207.600 151.230 207.920 ;
        RECT 151.030 203.500 151.170 207.600 ;
        RECT 152.410 203.500 152.550 210.660 ;
        RECT 153.270 207.830 153.530 207.920 ;
        RECT 152.870 207.690 153.530 207.830 ;
        RECT 150.970 203.180 151.230 203.500 ;
        RECT 152.350 203.180 152.610 203.500 ;
        RECT 150.510 202.160 150.770 202.480 ;
        RECT 150.050 201.820 150.310 202.140 ;
        RECT 149.590 200.460 149.850 200.780 ;
        RECT 149.130 188.560 149.390 188.880 ;
        RECT 149.190 184.460 149.330 188.560 ;
        RECT 149.130 184.140 149.390 184.460 ;
        RECT 150.110 183.780 150.250 201.820 ;
        RECT 152.350 201.480 152.610 201.800 ;
        RECT 150.960 200.605 151.240 200.975 ;
        RECT 151.030 200.100 151.170 200.605 ;
        RECT 152.410 200.100 152.550 201.480 ;
        RECT 150.970 199.780 151.230 200.100 ;
        RECT 152.350 199.780 152.610 200.100 ;
        RECT 151.430 199.100 151.690 199.420 ;
        RECT 150.970 196.040 151.230 196.360 ;
        RECT 151.030 192.620 151.170 196.040 ;
        RECT 150.970 192.300 151.230 192.620 ;
        RECT 150.970 191.620 151.230 191.940 ;
        RECT 151.030 189.220 151.170 191.620 ;
        RECT 150.970 188.900 151.230 189.220 ;
        RECT 151.030 187.180 151.170 188.900 ;
        RECT 150.970 186.860 151.230 187.180 ;
        RECT 150.510 184.140 150.770 184.460 ;
        RECT 150.570 183.975 150.710 184.140 ;
        RECT 148.210 183.460 148.470 183.780 ;
        RECT 150.050 183.460 150.310 183.780 ;
        RECT 150.500 183.605 150.780 183.975 ;
        RECT 150.570 183.440 150.710 183.605 ;
        RECT 150.510 183.120 150.770 183.440 ;
        RECT 149.130 182.440 149.390 182.760 ;
        RECT 149.190 178.340 149.330 182.440 ;
        RECT 151.030 180.720 151.170 186.860 ;
        RECT 150.970 180.400 151.230 180.720 ;
        RECT 149.130 178.020 149.390 178.340 ;
        RECT 147.290 177.000 147.550 177.320 ;
        RECT 149.190 176.300 149.330 178.020 ;
        RECT 151.490 176.300 151.630 199.100 ;
        RECT 152.350 197.060 152.610 197.380 ;
        RECT 151.890 196.380 152.150 196.700 ;
        RECT 151.950 194.660 152.090 196.380 ;
        RECT 151.890 194.340 152.150 194.660 ;
        RECT 151.890 191.280 152.150 191.600 ;
        RECT 151.950 189.560 152.090 191.280 ;
        RECT 152.410 190.920 152.550 197.060 ;
        RECT 152.870 196.360 153.010 207.690 ;
        RECT 153.270 207.600 153.530 207.690 ;
        RECT 153.270 206.920 153.530 207.240 ;
        RECT 153.330 206.220 153.470 206.920 ;
        RECT 153.270 205.900 153.530 206.220 ;
        RECT 153.270 202.160 153.530 202.480 ;
        RECT 153.330 198.060 153.470 202.160 ;
        RECT 153.270 197.740 153.530 198.060 ;
        RECT 152.810 196.040 153.070 196.360 ;
        RECT 152.870 195.340 153.010 196.040 ;
        RECT 152.810 195.020 153.070 195.340 ;
        RECT 153.270 194.340 153.530 194.660 ;
        RECT 152.350 190.600 152.610 190.920 ;
        RECT 151.890 189.240 152.150 189.560 ;
        RECT 151.890 188.560 152.150 188.880 ;
        RECT 151.950 184.120 152.090 188.560 ;
        RECT 152.410 185.820 152.550 190.600 ;
        RECT 152.810 188.900 153.070 189.220 ;
        RECT 152.870 186.160 153.010 188.900 ;
        RECT 152.810 185.840 153.070 186.160 ;
        RECT 152.350 185.500 152.610 185.820 ;
        RECT 152.350 184.140 152.610 184.460 ;
        RECT 151.890 183.800 152.150 184.120 ;
        RECT 151.890 182.440 152.150 182.760 ;
        RECT 151.950 180.720 152.090 182.440 ;
        RECT 151.890 180.400 152.150 180.720 ;
        RECT 149.130 175.980 149.390 176.300 ;
        RECT 151.430 175.980 151.690 176.300 ;
        RECT 151.950 175.280 152.090 180.400 ;
        RECT 152.410 179.020 152.550 184.140 ;
        RECT 152.870 181.740 153.010 185.840 ;
        RECT 152.810 181.420 153.070 181.740 ;
        RECT 152.350 178.700 152.610 179.020 ;
        RECT 153.330 176.300 153.470 194.340 ;
        RECT 153.790 191.600 153.930 210.660 ;
        RECT 154.250 208.260 154.390 211.600 ;
        RECT 154.190 207.940 154.450 208.260 ;
        RECT 154.190 197.400 154.450 197.720 ;
        RECT 153.730 191.280 153.990 191.600 ;
        RECT 154.250 187.180 154.390 197.400 ;
        RECT 154.190 186.860 154.450 187.180 ;
        RECT 154.250 183.780 154.390 186.860 ;
        RECT 154.710 184.460 154.850 216.100 ;
        RECT 155.110 213.040 155.370 213.360 ;
        RECT 155.170 211.320 155.310 213.040 ;
        RECT 157.460 211.825 159.000 212.195 ;
        RECT 155.110 211.000 155.370 211.320 ;
        RECT 155.110 207.940 155.370 208.260 ;
        RECT 154.650 184.140 154.910 184.460 ;
        RECT 155.170 183.780 155.310 207.940 ;
        RECT 157.460 206.385 159.000 206.755 ;
        RECT 157.460 200.945 159.000 201.315 ;
        RECT 157.460 195.505 159.000 195.875 ;
        RECT 157.460 190.065 159.000 190.435 ;
        RECT 155.570 186.180 155.830 186.500 ;
        RECT 155.630 184.460 155.770 186.180 ;
        RECT 157.460 184.625 159.000 184.995 ;
        RECT 155.570 184.140 155.830 184.460 ;
        RECT 154.190 183.460 154.450 183.780 ;
        RECT 155.110 183.460 155.370 183.780 ;
        RECT 154.250 179.020 154.390 183.460 ;
        RECT 155.170 179.020 155.310 183.460 ;
        RECT 157.460 179.185 159.000 179.555 ;
        RECT 154.190 178.700 154.450 179.020 ;
        RECT 155.110 178.700 155.370 179.020 ;
        RECT 153.270 175.980 153.530 176.300 ;
        RECT 151.890 174.960 152.150 175.280 ;
        RECT 157.460 173.745 159.000 174.115 ;
        RECT 144.590 173.400 145.190 173.540 ;
        RECT 138.025 171.025 139.565 171.395 ;
        RECT 137.630 168.840 137.890 169.160 ;
        RECT 143.150 168.840 143.410 169.160 ;
        RECT 137.690 164.060 137.830 168.840 ;
        RECT 143.210 167.460 143.350 168.840 ;
        RECT 143.150 167.140 143.410 167.460 ;
        RECT 140.850 166.800 141.110 167.120 ;
        RECT 138.025 165.585 139.565 165.955 ;
        RECT 137.630 163.740 137.890 164.060 ;
        RECT 138.550 163.740 138.810 164.060 ;
        RECT 137.690 162.100 137.830 163.740 ;
        RECT 138.610 162.700 138.750 163.740 ;
        RECT 138.550 162.380 138.810 162.700 ;
        RECT 137.230 161.960 137.830 162.100 ;
        RECT 135.790 158.300 136.050 158.620 ;
        RECT 133.950 157.960 134.210 158.280 ;
        RECT 134.010 155.560 134.150 157.960 ;
        RECT 137.230 156.920 137.370 161.960 ;
        RECT 138.080 161.845 138.360 162.215 ;
        RECT 138.150 161.680 138.290 161.845 ;
        RECT 138.090 161.360 138.350 161.680 ;
        RECT 138.025 160.145 139.565 160.515 ;
        RECT 139.000 159.125 139.280 159.495 ;
        RECT 140.910 159.300 141.050 166.800 ;
        RECT 144.070 164.080 144.330 164.400 ;
        RECT 144.130 162.360 144.270 164.080 ;
        RECT 144.070 162.040 144.330 162.360 ;
        RECT 144.590 159.300 144.730 173.400 ;
        RECT 148.660 172.045 148.940 172.415 ;
        RECT 148.730 168.140 148.870 172.045 ;
        RECT 149.580 170.005 149.860 170.375 ;
        RECT 148.670 167.820 148.930 168.140 ;
        RECT 149.650 167.460 149.790 170.005 ;
        RECT 157.460 168.305 159.000 168.675 ;
        RECT 149.590 167.140 149.850 167.460 ;
        RECT 147.750 166.120 148.010 166.440 ;
        RECT 150.970 166.120 151.230 166.440 ;
        RECT 145.450 164.080 145.710 164.400 ;
        RECT 144.990 163.740 145.250 164.060 ;
        RECT 145.050 162.700 145.190 163.740 ;
        RECT 144.990 162.380 145.250 162.700 ;
        RECT 139.070 158.280 139.210 159.125 ;
        RECT 140.850 158.980 141.110 159.300 ;
        RECT 144.530 158.980 144.790 159.300 ;
        RECT 137.630 157.960 137.890 158.280 ;
        RECT 139.010 157.960 139.270 158.280 ;
        RECT 141.770 157.960 142.030 158.280 ;
        RECT 137.170 156.600 137.430 156.920 ;
        RECT 133.950 155.240 134.210 155.560 ;
        RECT 137.690 154.540 137.830 157.960 ;
        RECT 141.830 157.260 141.970 157.960 ;
        RECT 141.770 156.940 142.030 157.260 ;
        RECT 145.510 156.920 145.650 164.080 ;
        RECT 147.810 162.360 147.950 166.120 ;
        RECT 151.030 164.400 151.170 166.120 ;
        RECT 150.970 164.080 151.230 164.400 ;
        RECT 147.750 162.040 148.010 162.360 ;
        RECT 151.030 159.980 151.170 164.080 ;
        RECT 157.460 162.865 159.000 163.235 ;
        RECT 150.970 159.660 151.230 159.980 ;
        RECT 157.460 157.425 159.000 157.795 ;
        RECT 145.450 156.600 145.710 156.920 ;
        RECT 143.150 155.920 143.410 156.240 ;
        RECT 138.025 154.705 139.565 155.075 ;
        RECT 143.210 154.540 143.350 155.920 ;
        RECT 137.630 154.220 137.890 154.540 ;
        RECT 143.150 154.220 143.410 154.540 ;
        RECT 137.170 153.880 137.430 154.200 ;
        RECT 133.490 152.860 133.750 153.180 ;
        RECT 132.570 150.910 133.230 151.050 ;
        RECT 132.570 150.820 132.830 150.910 ;
        RECT 131.650 148.670 131.910 148.760 ;
        RECT 131.650 148.530 132.310 148.670 ;
        RECT 131.650 148.440 131.910 148.530 ;
        RECT 131.190 147.760 131.450 148.080 ;
        RECT 130.730 147.080 130.990 147.400 ;
        RECT 130.790 145.700 130.930 147.080 ;
        RECT 131.250 145.700 131.390 147.760 ;
        RECT 131.650 146.060 131.910 146.380 ;
        RECT 130.730 145.380 130.990 145.700 ;
        RECT 131.190 145.380 131.450 145.700 ;
        RECT 131.710 145.360 131.850 146.060 ;
        RECT 131.650 145.040 131.910 145.360 ;
        RECT 130.730 144.590 130.990 144.680 ;
        RECT 130.330 144.450 130.990 144.590 ;
        RECT 130.730 144.360 130.990 144.450 ;
        RECT 131.190 144.360 131.450 144.680 ;
        RECT 131.650 144.360 131.910 144.680 ;
        RECT 129.350 143.340 129.610 143.660 ;
        RECT 127.970 142.320 128.230 142.640 ;
        RECT 128.430 142.320 128.690 142.640 ;
        RECT 128.890 142.320 129.150 142.640 ;
        RECT 128.030 141.960 128.170 142.320 ;
        RECT 127.970 141.640 128.230 141.960 ;
        RECT 128.490 141.815 128.630 142.320 ;
        RECT 128.420 141.445 128.700 141.815 ;
        RECT 127.970 140.170 128.230 140.260 ;
        RECT 127.570 140.030 128.230 140.170 ;
        RECT 127.970 139.940 128.230 140.030 ;
        RECT 127.510 139.095 127.770 139.240 ;
        RECT 127.500 138.725 127.780 139.095 ;
        RECT 127.050 136.880 127.310 137.200 ;
        RECT 126.590 134.160 126.850 134.480 ;
        RECT 126.650 132.100 126.790 134.160 ;
        RECT 128.030 134.140 128.170 139.940 ;
        RECT 128.950 138.220 129.090 142.320 ;
        RECT 128.890 137.900 129.150 138.220 ;
        RECT 128.890 135.180 129.150 135.500 ;
        RECT 128.950 135.015 129.090 135.180 ;
        RECT 128.430 134.500 128.690 134.820 ;
        RECT 128.880 134.645 129.160 135.015 ;
        RECT 127.970 133.820 128.230 134.140 ;
        RECT 127.050 133.480 127.310 133.800 ;
        RECT 127.510 133.480 127.770 133.800 ;
        RECT 126.590 131.780 126.850 132.100 ;
        RECT 126.120 128.525 126.400 128.895 ;
        RECT 125.210 125.660 125.470 125.980 ;
        RECT 126.590 125.660 126.850 125.980 ;
        RECT 123.830 124.190 124.090 124.280 ;
        RECT 123.830 124.050 124.490 124.190 ;
        RECT 123.830 123.960 124.090 124.050 ;
        RECT 123.830 123.510 124.090 123.600 ;
        RECT 123.430 123.370 124.090 123.510 ;
        RECT 123.830 123.280 124.090 123.370 ;
        RECT 123.370 122.600 123.630 122.920 ;
        RECT 118.770 121.580 119.030 121.900 ;
        RECT 121.990 121.580 122.250 121.900 ;
        RECT 122.910 121.580 123.170 121.900 ;
        RECT 117.390 121.240 117.650 121.560 ;
        RECT 109.570 120.900 109.830 121.220 ;
        RECT 123.430 119.940 123.570 122.600 ;
        RECT 123.890 120.830 124.030 123.280 ;
        RECT 124.350 121.220 124.490 124.050 ;
        RECT 124.750 123.960 125.010 124.280 ;
        RECT 126.130 123.850 126.390 123.940 ;
        RECT 126.650 123.850 126.790 125.660 ;
        RECT 127.110 124.620 127.250 133.480 ;
        RECT 127.570 131.760 127.710 133.480 ;
        RECT 127.510 131.440 127.770 131.760 ;
        RECT 127.960 131.245 128.240 131.615 ;
        RECT 127.970 131.100 128.230 131.245 ;
        RECT 128.490 129.380 128.630 134.500 ;
        RECT 129.410 132.780 129.550 143.340 ;
        RECT 129.810 143.000 130.070 143.320 ;
        RECT 129.870 140.260 130.010 143.000 ;
        RECT 130.790 140.260 130.930 144.360 ;
        RECT 131.250 143.660 131.390 144.360 ;
        RECT 131.190 143.340 131.450 143.660 ;
        RECT 131.190 141.640 131.450 141.960 ;
        RECT 131.250 141.135 131.390 141.640 ;
        RECT 131.180 140.765 131.460 141.135 ;
        RECT 131.190 140.620 131.450 140.765 ;
        RECT 129.810 139.940 130.070 140.260 ;
        RECT 130.730 139.940 130.990 140.260 ;
        RECT 129.810 138.920 130.070 139.240 ;
        RECT 130.270 138.920 130.530 139.240 ;
        RECT 129.870 138.220 130.010 138.920 ;
        RECT 129.810 137.900 130.070 138.220 ;
        RECT 129.800 136.685 130.080 137.055 ;
        RECT 129.810 136.540 130.070 136.685 ;
        RECT 130.330 133.710 130.470 138.920 ;
        RECT 131.710 135.500 131.850 144.360 ;
        RECT 132.170 140.940 132.310 148.530 ;
        RECT 132.630 148.420 132.770 150.820 ;
        RECT 132.570 148.100 132.830 148.420 ;
        RECT 133.950 148.100 134.210 148.420 ;
        RECT 133.490 147.650 133.750 147.740 ;
        RECT 133.090 147.510 133.750 147.650 ;
        RECT 133.090 146.380 133.230 147.510 ;
        RECT 133.490 147.420 133.750 147.510 ;
        RECT 133.090 146.060 133.450 146.380 ;
        RECT 133.090 141.960 133.230 146.060 ;
        RECT 134.010 145.700 134.150 148.100 ;
        RECT 134.410 147.080 134.670 147.400 ;
        RECT 133.950 145.380 134.210 145.700 ;
        RECT 133.480 143.485 133.760 143.855 ;
        RECT 133.550 142.640 133.690 143.485 ;
        RECT 133.490 142.320 133.750 142.640 ;
        RECT 133.030 141.640 133.290 141.960 ;
        RECT 132.110 140.620 132.370 140.940 ;
        RECT 132.100 140.085 132.380 140.455 ;
        RECT 131.650 135.180 131.910 135.500 ;
        RECT 131.710 134.820 131.850 135.180 ;
        RECT 131.650 134.500 131.910 134.820 ;
        RECT 131.650 133.820 131.910 134.140 ;
        RECT 132.170 134.050 132.310 140.085 ;
        RECT 132.570 139.775 132.830 139.920 ;
        RECT 132.560 139.405 132.840 139.775 ;
        RECT 133.550 139.580 133.690 142.320 ;
        RECT 133.030 139.260 133.290 139.580 ;
        RECT 133.490 139.260 133.750 139.580 ;
        RECT 132.570 138.920 132.830 139.240 ;
        RECT 132.630 138.220 132.770 138.920 ;
        RECT 132.570 137.900 132.830 138.220 ;
        RECT 132.630 135.160 132.770 137.900 ;
        RECT 133.090 137.200 133.230 139.260 ;
        RECT 133.550 138.220 133.690 139.260 ;
        RECT 133.490 137.900 133.750 138.220 ;
        RECT 133.030 136.880 133.290 137.200 ;
        RECT 133.490 136.540 133.750 136.860 ;
        RECT 132.570 134.840 132.830 135.160 ;
        RECT 132.570 134.050 132.830 134.140 ;
        RECT 132.170 133.910 132.830 134.050 ;
        RECT 132.570 133.820 132.830 133.910 ;
        RECT 131.190 133.710 131.450 133.800 ;
        RECT 130.330 133.570 131.450 133.710 ;
        RECT 129.350 132.460 129.610 132.780 ;
        RECT 129.410 129.380 129.550 132.460 ;
        RECT 130.330 130.060 130.470 133.570 ;
        RECT 131.190 133.480 131.450 133.570 ;
        RECT 131.710 132.010 131.850 133.820 ;
        RECT 133.550 133.800 133.690 136.540 ;
        RECT 134.470 135.160 134.610 147.080 ;
        RECT 135.790 144.360 136.050 144.680 ;
        RECT 135.850 142.640 135.990 144.360 ;
        RECT 135.790 142.320 136.050 142.640 ;
        RECT 136.710 142.320 136.970 142.640 ;
        RECT 134.870 141.640 135.130 141.960 ;
        RECT 134.930 140.260 135.070 141.640 ;
        RECT 134.870 139.940 135.130 140.260 ;
        RECT 134.930 136.520 135.070 139.940 ;
        RECT 135.330 139.600 135.590 139.920 ;
        RECT 135.390 139.095 135.530 139.600 ;
        RECT 135.320 138.725 135.600 139.095 ;
        RECT 134.870 136.200 135.130 136.520 ;
        RECT 134.410 135.015 134.670 135.160 ;
        RECT 133.950 134.500 134.210 134.820 ;
        RECT 134.400 134.645 134.680 135.015 ;
        RECT 133.490 133.480 133.750 133.800 ;
        RECT 132.110 132.010 132.370 132.100 ;
        RECT 131.710 131.870 132.370 132.010 ;
        RECT 132.110 131.780 132.370 131.870 ;
        RECT 132.570 131.440 132.830 131.760 ;
        RECT 130.270 129.740 130.530 130.060 ;
        RECT 132.630 129.380 132.770 131.440 ;
        RECT 133.490 131.100 133.750 131.420 ;
        RECT 133.550 130.060 133.690 131.100 ;
        RECT 133.490 129.740 133.750 130.060 ;
        RECT 128.430 129.060 128.690 129.380 ;
        RECT 129.350 129.060 129.610 129.380 ;
        RECT 132.570 129.060 132.830 129.380 ;
        RECT 134.010 129.040 134.150 134.500 ;
        RECT 134.400 133.965 134.680 134.335 ;
        RECT 134.470 131.760 134.610 133.965 ;
        RECT 134.870 133.480 135.130 133.800 ;
        RECT 134.930 131.760 135.070 133.480 ;
        RECT 135.390 131.760 135.530 138.725 ;
        RECT 135.780 137.365 136.060 137.735 ;
        RECT 135.850 136.520 135.990 137.365 ;
        RECT 136.770 136.860 136.910 142.320 ;
        RECT 136.710 136.540 136.970 136.860 ;
        RECT 135.790 136.430 136.050 136.520 ;
        RECT 135.790 136.290 136.450 136.430 ;
        RECT 135.790 136.200 136.050 136.290 ;
        RECT 136.310 131.760 136.450 136.290 ;
        RECT 134.410 131.440 134.670 131.760 ;
        RECT 134.870 131.440 135.130 131.760 ;
        RECT 135.330 131.440 135.590 131.760 ;
        RECT 135.790 131.615 136.050 131.760 ;
        RECT 134.410 130.760 134.670 131.080 ;
        RECT 133.950 128.720 134.210 129.040 ;
        RECT 134.470 128.700 134.610 130.760 ;
        RECT 128.430 128.380 128.690 128.700 ;
        RECT 134.410 128.380 134.670 128.700 ;
        RECT 128.490 127.340 128.630 128.380 ;
        RECT 128.430 127.020 128.690 127.340 ;
        RECT 134.930 127.000 135.070 131.440 ;
        RECT 135.780 131.245 136.060 131.615 ;
        RECT 136.250 131.440 136.510 131.760 ;
        RECT 137.230 129.380 137.370 153.880 ;
        RECT 140.850 153.200 141.110 153.520 ;
        RECT 139.930 152.520 140.190 152.840 ;
        RECT 138.025 149.265 139.565 149.635 ;
        RECT 139.990 147.400 140.130 152.520 ;
        RECT 140.390 150.480 140.650 150.800 ;
        RECT 139.930 147.080 140.190 147.400 ;
        RECT 140.450 146.380 140.590 150.480 ;
        RECT 140.390 146.060 140.650 146.380 ;
        RECT 138.025 143.825 139.565 144.195 ;
        RECT 140.910 143.660 141.050 153.200 ;
        RECT 145.510 151.820 145.650 156.600 ;
        RECT 157.460 151.985 159.000 152.355 ;
        RECT 141.310 151.500 141.570 151.820 ;
        RECT 145.450 151.500 145.710 151.820 ;
        RECT 141.370 148.760 141.510 151.500 ;
        RECT 143.610 150.820 143.870 151.140 ;
        RECT 141.760 150.285 142.040 150.655 ;
        RECT 141.770 150.140 142.030 150.285 ;
        RECT 141.310 148.440 141.570 148.760 ;
        RECT 141.370 145.700 141.510 148.440 ;
        RECT 141.310 145.380 141.570 145.700 ;
        RECT 141.830 143.740 141.970 150.140 ;
        RECT 142.690 149.800 142.950 150.120 ;
        RECT 142.750 146.040 142.890 149.800 ;
        RECT 142.690 145.720 142.950 146.040 ;
        RECT 143.150 144.360 143.410 144.680 ;
        RECT 141.830 143.660 142.430 143.740 ;
        RECT 143.210 143.660 143.350 144.360 ;
        RECT 140.850 143.340 141.110 143.660 ;
        RECT 141.770 143.600 142.430 143.660 ;
        RECT 141.770 143.340 142.030 143.600 ;
        RECT 138.080 142.125 138.360 142.495 ;
        RECT 140.390 142.320 140.650 142.640 ;
        RECT 138.090 141.980 138.350 142.125 ;
        RECT 139.930 141.980 140.190 142.300 ;
        RECT 138.025 138.385 139.565 138.755 ;
        RECT 138.090 136.200 138.350 136.520 ;
        RECT 138.150 134.335 138.290 136.200 ;
        RECT 137.630 133.820 137.890 134.140 ;
        RECT 138.080 133.965 138.360 134.335 ;
        RECT 137.690 131.420 137.830 133.820 ;
        RECT 138.025 132.945 139.565 133.315 ;
        RECT 139.990 131.760 140.130 141.980 ;
        RECT 140.450 140.600 140.590 142.320 ;
        RECT 141.770 141.980 142.030 142.300 ;
        RECT 140.390 140.280 140.650 140.600 ;
        RECT 140.450 137.540 140.590 140.280 ;
        RECT 140.390 137.220 140.650 137.540 ;
        RECT 141.830 137.200 141.970 141.980 ;
        RECT 142.290 140.260 142.430 143.600 ;
        RECT 143.150 143.340 143.410 143.660 ;
        RECT 143.670 142.640 143.810 150.820 ;
        RECT 144.990 148.780 145.250 149.100 ;
        RECT 144.070 147.420 144.330 147.740 ;
        RECT 143.610 142.320 143.870 142.640 ;
        RECT 144.130 140.940 144.270 147.420 ;
        RECT 145.050 146.380 145.190 148.780 ;
        RECT 157.460 146.545 159.000 146.915 ;
        RECT 144.990 146.060 145.250 146.380 ;
        RECT 146.830 142.320 147.090 142.640 ;
        RECT 144.990 141.640 145.250 141.960 ;
        RECT 144.070 140.620 144.330 140.940 ;
        RECT 142.230 139.940 142.490 140.260 ;
        RECT 142.290 139.240 142.430 139.940 ;
        RECT 145.050 139.920 145.190 141.640 ;
        RECT 146.890 140.940 147.030 142.320 ;
        RECT 148.210 141.640 148.470 141.960 ;
        RECT 146.830 140.620 147.090 140.940 ;
        RECT 148.270 140.260 148.410 141.640 ;
        RECT 157.460 141.105 159.000 141.475 ;
        RECT 148.210 139.940 148.470 140.260 ;
        RECT 144.990 139.600 145.250 139.920 ;
        RECT 145.450 139.260 145.710 139.580 ;
        RECT 142.230 138.920 142.490 139.240 ;
        RECT 143.150 138.920 143.410 139.240 ;
        RECT 143.210 138.220 143.350 138.920 ;
        RECT 143.150 137.900 143.410 138.220 ;
        RECT 141.770 136.880 142.030 137.200 ;
        RECT 140.390 136.540 140.650 136.860 ;
        RECT 139.930 131.440 140.190 131.760 ;
        RECT 137.630 131.100 137.890 131.420 ;
        RECT 137.170 129.060 137.430 129.380 ;
        RECT 135.790 128.720 136.050 129.040 ;
        RECT 135.850 127.340 135.990 128.720 ;
        RECT 135.790 127.020 136.050 127.340 ;
        RECT 134.870 126.680 135.130 127.000 ;
        RECT 137.230 126.660 137.370 129.060 ;
        RECT 138.025 127.505 139.565 127.875 ;
        RECT 137.170 126.340 137.430 126.660 ;
        RECT 127.970 126.000 128.230 126.320 ;
        RECT 127.050 124.300 127.310 124.620 ;
        RECT 126.130 123.710 126.790 123.850 ;
        RECT 126.130 123.620 126.390 123.710 ;
        RECT 126.650 121.900 126.790 123.710 ;
        RECT 127.510 123.620 127.770 123.940 ;
        RECT 127.570 121.900 127.710 123.620 ;
        RECT 128.030 123.600 128.170 126.000 ;
        RECT 132.110 125.320 132.370 125.640 ;
        RECT 136.710 125.320 136.970 125.640 ;
        RECT 132.170 123.940 132.310 125.320 ;
        RECT 133.030 124.300 133.290 124.620 ;
        RECT 128.430 123.620 128.690 123.940 ;
        RECT 129.810 123.620 130.070 123.940 ;
        RECT 132.110 123.620 132.370 123.940 ;
        RECT 127.970 123.280 128.230 123.600 ;
        RECT 126.590 121.580 126.850 121.900 ;
        RECT 127.510 121.580 127.770 121.900 ;
        RECT 128.490 121.560 128.630 123.620 ;
        RECT 129.870 121.900 130.010 123.620 ;
        RECT 130.730 123.280 130.990 123.600 ;
        RECT 129.810 121.580 130.070 121.900 ;
        RECT 130.790 121.560 130.930 123.280 ;
        RECT 132.570 122.940 132.830 123.260 ;
        RECT 128.430 121.240 128.690 121.560 ;
        RECT 130.730 121.240 130.990 121.560 ;
        RECT 124.290 120.900 124.550 121.220 ;
        RECT 131.190 120.900 131.450 121.220 ;
        RECT 123.830 120.510 124.090 120.830 ;
        RECT 124.290 120.220 124.550 120.540 ;
        RECT 124.350 119.940 124.490 120.220 ;
        RECT 123.430 119.800 124.490 119.940 ;
        RECT 118.590 119.345 120.130 119.715 ;
        RECT 131.250 119.180 131.390 120.900 ;
        RECT 132.630 120.540 132.770 122.940 ;
        RECT 133.090 121.900 133.230 124.300 ;
        RECT 136.770 123.260 136.910 125.320 ;
        RECT 136.710 122.940 136.970 123.260 ;
        RECT 138.025 122.065 139.565 122.435 ;
        RECT 133.030 121.580 133.290 121.900 ;
        RECT 139.990 121.220 140.130 131.440 ;
        RECT 140.450 131.420 140.590 136.540 ;
        RECT 141.310 136.200 141.570 136.520 ;
        RECT 140.390 131.100 140.650 131.420 ;
        RECT 140.850 131.100 141.110 131.420 ;
        RECT 140.910 130.060 141.050 131.100 ;
        RECT 141.370 130.255 141.510 136.200 ;
        RECT 140.850 129.740 141.110 130.060 ;
        RECT 141.300 129.885 141.580 130.255 ;
        RECT 143.210 126.855 143.350 137.900 ;
        RECT 145.510 137.200 145.650 139.260 ;
        RECT 147.750 138.920 148.010 139.240 ;
        RECT 147.810 137.200 147.950 138.920 ;
        RECT 145.450 136.880 145.710 137.200 ;
        RECT 147.750 136.880 148.010 137.200 ;
        RECT 148.210 136.200 148.470 136.520 ;
        RECT 148.270 133.800 148.410 136.200 ;
        RECT 157.460 135.665 159.000 136.035 ;
        RECT 148.210 133.480 148.470 133.800 ;
        RECT 157.460 130.225 159.000 130.595 ;
        RECT 143.140 126.485 143.420 126.855 ;
        RECT 157.460 124.785 159.000 125.155 ;
        RECT 139.930 120.900 140.190 121.220 ;
        RECT 132.570 120.220 132.830 120.540 ;
        RECT 157.460 119.345 159.000 119.715 ;
        RECT 131.190 118.860 131.450 119.180 ;
        RECT 109.110 118.520 109.370 118.840 ;
        RECT 95.770 118.180 96.030 118.500 ;
        RECT 98.530 118.180 98.790 118.500 ;
        RECT 95.310 117.840 95.570 118.160 ;
        RECT 21.415 116.625 22.955 116.995 ;
        RECT 60.285 116.625 61.825 116.995 ;
        RECT 99.155 116.625 100.695 116.995 ;
        RECT 138.025 116.625 139.565 116.995 ;
        RECT 40.850 113.905 42.390 114.275 ;
        RECT 79.720 113.905 81.260 114.275 ;
        RECT 118.590 113.905 120.130 114.275 ;
        RECT 157.460 113.905 159.000 114.275 ;
        RECT 11.340 111.590 11.640 111.600 ;
        RECT 11.305 111.310 11.675 111.590 ;
        RECT 11.340 110.700 11.640 111.310 ;
        RECT 16.130 111.270 16.430 111.280 ;
        RECT 16.095 110.990 16.465 111.270 ;
        RECT 29.740 111.000 30.040 111.010 ;
        RECT 16.130 110.490 16.430 110.990 ;
        RECT 18.700 110.980 19.000 110.990 ;
        RECT 26.060 110.980 26.360 110.990 ;
        RECT 18.665 110.700 19.035 110.980 ;
        RECT 23.740 110.950 24.040 110.960 ;
        RECT 18.700 110.320 19.000 110.700 ;
        RECT 23.705 110.670 24.075 110.950 ;
        RECT 26.025 110.700 26.395 110.980 ;
        RECT 29.705 110.720 30.075 111.000 ;
        RECT 23.740 110.390 24.040 110.670 ;
        RECT 26.060 110.450 26.360 110.700 ;
        RECT 29.740 110.390 30.040 110.720 ;
        RECT 3.980 109.100 4.280 109.110 ;
        RECT 3.945 108.820 4.315 109.100 ;
        RECT 3.980 108.170 4.280 108.820 ;
        RECT 6.680 108.490 6.980 108.500 ;
        RECT 6.645 108.210 7.015 108.490 ;
        RECT 6.680 107.560 6.980 108.210 ;
        RECT 31.450 99.510 32.450 99.540 ;
        RECT 3.490 98.510 32.450 99.510 ;
        RECT 31.450 98.480 32.450 98.510 ;
        RECT 6.320 97.510 7.320 97.540 ;
        RECT 31.350 97.510 32.350 97.540 ;
        RECT 6.320 96.510 32.350 97.510 ;
        RECT 6.320 96.480 7.320 96.510 ;
        RECT 31.350 96.480 32.350 96.510 ;
        RECT 31.450 95.700 32.450 95.730 ;
        RECT 11.000 94.700 32.450 95.700 ;
        RECT 31.450 94.670 32.450 94.700 ;
        RECT 15.790 92.590 32.480 93.590 ;
        RECT 21.100 90.390 32.380 91.390 ;
        RECT 31.450 89.490 32.450 89.520 ;
        RECT 23.300 88.490 32.450 89.490 ;
        RECT 31.450 88.460 32.450 88.490 ;
        RECT 31.750 87.580 32.750 87.610 ;
        RECT 26.810 86.580 32.750 87.580 ;
        RECT 31.750 86.550 32.750 86.580 ;
        RECT 103.000 81.975 104.000 82.000 ;
        RECT 102.980 81.025 104.020 81.975 ;
        RECT 103.000 77.670 104.000 81.025 ;
        RECT 137.870 35.700 138.530 36.300 ;
        RECT 137.900 26.400 138.500 35.700 ;
        RECT 147.325 26.400 147.875 26.420 ;
        RECT 137.900 25.800 147.900 26.400 ;
        RECT 147.325 25.780 147.875 25.800 ;
      LAYER met3 ;
        RECT 68.595 222.020 68.925 222.035 ;
        RECT 73.860 222.020 74.240 222.030 ;
        RECT 68.595 221.720 74.240 222.020 ;
        RECT 68.595 221.705 68.925 221.720 ;
        RECT 73.860 221.710 74.240 221.720 ;
        RECT 22.595 221.350 22.925 221.355 ;
        RECT 22.340 221.340 22.925 221.350 ;
        RECT 48.100 221.340 48.480 221.350 ;
        RECT 62.615 221.340 62.945 221.355 ;
        RECT 22.340 221.040 23.150 221.340 ;
        RECT 48.100 221.040 62.945 221.340 ;
        RECT 22.340 221.030 22.925 221.040 ;
        RECT 48.100 221.030 48.480 221.040 ;
        RECT 22.595 221.025 22.925 221.030 ;
        RECT 62.615 221.025 62.945 221.040 ;
        RECT 68.595 221.340 68.925 221.355 ;
        RECT 81.220 221.340 81.600 221.350 ;
        RECT 68.595 221.040 81.600 221.340 ;
        RECT 68.595 221.025 68.925 221.040 ;
        RECT 81.220 221.030 81.600 221.040 ;
        RECT 125.380 221.340 125.760 221.350 ;
        RECT 130.235 221.340 130.565 221.355 ;
        RECT 125.380 221.040 130.565 221.340 ;
        RECT 125.380 221.030 125.760 221.040 ;
        RECT 130.235 221.025 130.565 221.040 ;
        RECT 143.780 221.340 144.160 221.350 ;
        RECT 148.635 221.340 148.965 221.355 ;
        RECT 143.780 221.040 148.965 221.340 ;
        RECT 143.780 221.030 144.160 221.040 ;
        RECT 148.635 221.025 148.965 221.040 ;
        RECT 33.380 220.660 33.760 220.670 ;
        RECT 35.015 220.660 35.345 220.675 ;
        RECT 33.380 220.360 35.345 220.660 ;
        RECT 33.380 220.350 33.760 220.360 ;
        RECT 35.015 220.345 35.345 220.360 ;
        RECT 37.060 220.660 37.440 220.670 ;
        RECT 44.215 220.660 44.545 220.675 ;
        RECT 37.060 220.360 44.545 220.660 ;
        RECT 37.060 220.350 37.440 220.360 ;
        RECT 44.215 220.345 44.545 220.360 ;
        RECT 62.820 220.660 63.200 220.670 ;
        RECT 69.055 220.660 69.385 220.675 ;
        RECT 62.820 220.360 69.385 220.660 ;
        RECT 62.820 220.350 63.200 220.360 ;
        RECT 69.055 220.345 69.385 220.360 ;
        RECT 121.700 220.660 122.080 220.670 ;
        RECT 123.335 220.660 123.665 220.675 ;
        RECT 121.700 220.360 123.665 220.660 ;
        RECT 121.700 220.350 122.080 220.360 ;
        RECT 123.335 220.345 123.665 220.360 ;
        RECT 129.060 220.660 129.440 220.670 ;
        RECT 132.995 220.660 133.325 220.675 ;
        RECT 140.355 220.670 140.685 220.675 ;
        RECT 129.060 220.360 133.325 220.660 ;
        RECT 129.060 220.350 129.440 220.360 ;
        RECT 132.995 220.345 133.325 220.360 ;
        RECT 140.100 220.660 140.685 220.670 ;
        RECT 147.460 220.660 147.840 220.670 ;
        RECT 150.015 220.660 150.345 220.675 ;
        RECT 151.395 220.670 151.725 220.675 ;
        RECT 151.140 220.660 151.725 220.670 ;
        RECT 140.100 220.360 140.910 220.660 ;
        RECT 147.460 220.360 150.345 220.660 ;
        RECT 150.940 220.360 151.725 220.660 ;
        RECT 140.100 220.350 140.685 220.360 ;
        RECT 147.460 220.350 147.840 220.360 ;
        RECT 140.355 220.345 140.685 220.350 ;
        RECT 150.015 220.345 150.345 220.360 ;
        RECT 151.140 220.350 151.725 220.360 ;
        RECT 151.395 220.345 151.725 220.350 ;
        RECT 21.395 220.005 22.975 220.335 ;
        RECT 60.265 220.005 61.845 220.335 ;
        RECT 99.135 220.005 100.715 220.335 ;
        RECT 138.005 220.005 139.585 220.335 ;
        RECT 66.755 219.990 67.085 219.995 ;
        RECT 66.500 219.980 67.085 219.990 ;
        RECT 66.300 219.680 67.085 219.980 ;
        RECT 66.500 219.670 67.085 219.680 ;
        RECT 132.740 219.980 133.120 219.990 ;
        RECT 137.135 219.980 137.465 219.995 ;
        RECT 132.740 219.680 137.465 219.980 ;
        RECT 132.740 219.670 133.120 219.680 ;
        RECT 66.755 219.665 67.085 219.670 ;
        RECT 137.135 219.665 137.465 219.680 ;
        RECT 18.660 219.300 19.040 219.310 ;
        RECT 24.895 219.300 25.225 219.315 ;
        RECT 18.660 219.000 25.225 219.300 ;
        RECT 18.660 218.990 19.040 219.000 ;
        RECT 24.895 218.985 25.225 219.000 ;
        RECT 67.675 219.300 68.005 219.315 ;
        RECT 70.180 219.300 70.560 219.310 ;
        RECT 67.675 219.000 70.560 219.300 ;
        RECT 67.675 218.985 68.005 219.000 ;
        RECT 70.180 218.990 70.560 219.000 ;
        RECT 73.655 219.300 73.985 219.315 ;
        RECT 88.580 219.300 88.960 219.310 ;
        RECT 73.655 219.000 88.960 219.300 ;
        RECT 73.655 218.985 73.985 219.000 ;
        RECT 88.580 218.990 88.960 219.000 ;
        RECT 136.420 219.300 136.800 219.310 ;
        RECT 138.515 219.300 138.845 219.315 ;
        RECT 136.420 219.000 138.845 219.300 ;
        RECT 136.420 218.990 136.800 219.000 ;
        RECT 138.515 218.985 138.845 219.000 ;
        RECT 75.495 218.620 75.825 218.635 ;
        RECT 77.540 218.620 77.920 218.630 ;
        RECT 75.495 218.320 77.920 218.620 ;
        RECT 75.495 218.305 75.825 218.320 ;
        RECT 77.540 218.310 77.920 218.320 ;
        RECT 78.715 218.620 79.045 218.635 ;
        RECT 95.735 218.620 96.065 218.635 ;
        RECT 78.715 218.320 96.065 218.620 ;
        RECT 78.715 218.305 79.045 218.320 ;
        RECT 95.735 218.305 96.065 218.320 ;
        RECT 3.940 217.940 4.320 217.950 ;
        RECT 6.495 217.940 6.825 217.955 ;
        RECT 30.875 217.940 31.205 217.955 ;
        RECT 3.940 217.640 31.205 217.940 ;
        RECT 3.940 217.630 4.320 217.640 ;
        RECT 6.495 217.625 6.825 217.640 ;
        RECT 30.875 217.625 31.205 217.640 ;
        RECT 66.295 217.940 66.625 217.955 ;
        RECT 70.895 217.940 71.225 217.955 ;
        RECT 66.295 217.640 71.225 217.940 ;
        RECT 66.295 217.625 66.625 217.640 ;
        RECT 70.895 217.625 71.225 217.640 ;
        RECT 92.515 217.940 92.845 217.955 ;
        RECT 116.895 217.940 117.225 217.955 ;
        RECT 92.515 217.640 117.225 217.940 ;
        RECT 92.515 217.625 92.845 217.640 ;
        RECT 116.895 217.625 117.225 217.640 ;
        RECT 40.830 217.285 42.410 217.615 ;
        RECT 79.700 217.285 81.280 217.615 ;
        RECT 118.570 217.285 120.150 217.615 ;
        RECT 157.440 217.285 159.020 217.615 ;
        RECT 7.620 217.260 8.000 217.270 ;
        RECT 10.635 217.260 10.965 217.275 ;
        RECT 7.620 216.960 10.965 217.260 ;
        RECT 7.620 216.950 8.000 216.960 ;
        RECT 10.635 216.945 10.965 216.960 ;
        RECT 14.980 217.260 15.360 217.270 ;
        RECT 19.835 217.260 20.165 217.275 ;
        RECT 14.980 216.960 20.165 217.260 ;
        RECT 14.980 216.950 15.360 216.960 ;
        RECT 19.835 216.945 20.165 216.960 ;
        RECT 29.700 217.260 30.080 217.270 ;
        RECT 32.255 217.260 32.585 217.275 ;
        RECT 29.700 216.960 32.585 217.260 ;
        RECT 29.700 216.950 30.080 216.960 ;
        RECT 32.255 216.945 32.585 216.960 ;
        RECT 52.035 216.590 52.365 216.595 ;
        RECT 51.780 216.580 52.365 216.590 ;
        RECT 51.580 216.280 52.365 216.580 ;
        RECT 51.780 216.270 52.365 216.280 ;
        RECT 52.035 216.265 52.365 216.270 ;
        RECT 61.695 216.580 62.025 216.595 ;
        RECT 63.740 216.580 64.120 216.590 ;
        RECT 61.695 216.280 64.120 216.580 ;
        RECT 61.695 216.265 62.025 216.280 ;
        RECT 63.740 216.270 64.120 216.280 ;
        RECT 96.195 216.580 96.525 216.595 ;
        RECT 96.860 216.580 97.240 216.590 ;
        RECT 96.195 216.280 97.240 216.580 ;
        RECT 96.195 216.265 96.525 216.280 ;
        RECT 96.860 216.270 97.240 216.280 ;
        RECT 114.135 216.580 114.465 216.595 ;
        RECT 127.015 216.580 127.345 216.595 ;
        RECT 114.135 216.280 127.345 216.580 ;
        RECT 114.135 216.265 114.465 216.280 ;
        RECT 127.015 216.265 127.345 216.280 ;
        RECT 57.095 215.900 57.425 215.915 ;
        RECT 75.495 215.900 75.825 215.915 ;
        RECT 57.095 215.600 75.825 215.900 ;
        RECT 57.095 215.585 57.425 215.600 ;
        RECT 75.495 215.585 75.825 215.600 ;
        RECT 82.395 215.900 82.725 215.915 ;
        RECT 103.555 215.900 103.885 215.915 ;
        RECT 82.395 215.600 103.885 215.900 ;
        RECT 82.395 215.585 82.725 215.600 ;
        RECT 103.555 215.585 103.885 215.600 ;
        RECT 7.875 215.220 8.205 215.235 ;
        RECT 11.300 215.220 11.680 215.230 ;
        RECT 16.615 215.220 16.945 215.235 ;
        RECT 31.795 215.230 32.125 215.235 ;
        RECT 7.875 214.920 16.945 215.220 ;
        RECT 7.875 214.905 8.205 214.920 ;
        RECT 11.300 214.910 11.680 214.920 ;
        RECT 16.615 214.905 16.945 214.920 ;
        RECT 31.540 215.220 32.125 215.230 ;
        RECT 51.575 215.220 51.905 215.235 ;
        RECT 54.540 215.220 54.920 215.230 ;
        RECT 31.540 214.920 32.350 215.220 ;
        RECT 51.575 214.920 54.920 215.220 ;
        RECT 31.540 214.910 32.125 214.920 ;
        RECT 31.795 214.905 32.125 214.910 ;
        RECT 51.575 214.905 51.905 214.920 ;
        RECT 54.540 214.910 54.920 214.920 ;
        RECT 92.055 215.220 92.385 215.235 ;
        RECT 97.575 215.220 97.905 215.235 ;
        RECT 92.055 214.920 97.905 215.220 ;
        RECT 92.055 214.905 92.385 214.920 ;
        RECT 97.575 214.905 97.905 214.920 ;
        RECT 107.695 215.220 108.025 215.235 ;
        RECT 123.335 215.220 123.665 215.235 ;
        RECT 107.695 214.920 123.665 215.220 ;
        RECT 107.695 214.905 108.025 214.920 ;
        RECT 123.335 214.905 123.665 214.920 ;
        RECT 150.220 215.220 150.600 215.230 ;
        RECT 151.395 215.220 151.725 215.235 ;
        RECT 150.220 214.920 151.725 215.220 ;
        RECT 150.220 214.910 150.600 214.920 ;
        RECT 151.395 214.905 151.725 214.920 ;
        RECT 21.395 214.565 22.975 214.895 ;
        RECT 60.265 214.565 61.845 214.895 ;
        RECT 99.135 214.565 100.715 214.895 ;
        RECT 138.005 214.565 139.585 214.895 ;
        RECT 39.615 214.550 39.945 214.555 ;
        RECT 39.615 214.540 40.200 214.550 ;
        RECT 43.295 214.540 43.625 214.555 ;
        RECT 58.935 214.550 59.265 214.555 ;
        RECT 48.100 214.540 48.480 214.550 ;
        RECT 39.615 214.240 40.400 214.540 ;
        RECT 43.295 214.240 48.480 214.540 ;
        RECT 39.615 214.230 40.200 214.240 ;
        RECT 39.615 214.225 39.945 214.230 ;
        RECT 43.295 214.225 43.625 214.240 ;
        RECT 48.100 214.230 48.480 214.240 ;
        RECT 58.935 214.540 59.520 214.550 ;
        RECT 68.595 214.540 68.925 214.555 ;
        RECT 84.900 214.540 85.280 214.550 ;
        RECT 58.935 214.240 59.720 214.540 ;
        RECT 68.380 214.240 85.280 214.540 ;
        RECT 58.935 214.230 59.520 214.240 ;
        RECT 58.935 214.225 59.265 214.230 ;
        RECT 68.380 214.225 68.925 214.240 ;
        RECT 84.900 214.230 85.280 214.240 ;
        RECT 39.155 213.860 39.485 213.875 ;
        RECT 68.380 213.860 68.680 214.225 ;
        RECT 39.155 213.560 68.680 213.860 ;
        RECT 79.635 213.860 79.965 213.875 ;
        RECT 116.435 213.860 116.765 213.875 ;
        RECT 79.635 213.560 116.765 213.860 ;
        RECT 39.155 213.545 39.485 213.560 ;
        RECT 79.635 213.545 79.965 213.560 ;
        RECT 116.435 213.545 116.765 213.560 ;
        RECT 118.735 213.860 119.065 213.875 ;
        RECT 148.635 213.860 148.965 213.875 ;
        RECT 118.735 213.560 148.965 213.860 ;
        RECT 118.735 213.545 119.065 213.560 ;
        RECT 148.635 213.545 148.965 213.560 ;
        RECT 84.695 213.180 85.025 213.195 ;
        RECT 88.580 213.180 88.960 213.190 ;
        RECT 115.515 213.180 115.845 213.195 ;
        RECT 84.695 212.880 115.845 213.180 ;
        RECT 84.695 212.865 85.025 212.880 ;
        RECT 88.580 212.870 88.960 212.880 ;
        RECT 115.515 212.865 115.845 212.880 ;
        RECT 89.295 212.500 89.625 212.515 ;
        RECT 106.775 212.500 107.105 212.515 ;
        RECT 89.295 212.200 107.105 212.500 ;
        RECT 89.295 212.185 89.625 212.200 ;
        RECT 106.775 212.185 107.105 212.200 ;
        RECT 107.695 212.500 108.025 212.515 ;
        RECT 111.375 212.500 111.705 212.515 ;
        RECT 107.695 212.200 111.705 212.500 ;
        RECT 107.695 212.185 108.025 212.200 ;
        RECT 111.375 212.185 111.705 212.200 ;
        RECT 40.830 211.845 42.410 212.175 ;
        RECT 79.700 211.845 81.280 212.175 ;
        RECT 118.570 211.845 120.150 212.175 ;
        RECT 157.440 211.845 159.020 212.175 ;
        RECT 96.195 211.820 96.525 211.835 ;
        RECT 105.395 211.820 105.725 211.835 ;
        RECT 96.195 211.520 105.725 211.820 ;
        RECT 96.195 211.505 96.525 211.520 ;
        RECT 105.395 211.505 105.725 211.520 ;
        RECT 53.875 211.140 54.205 211.155 ;
        RECT 93.435 211.140 93.765 211.155 ;
        RECT 53.875 210.840 93.765 211.140 ;
        RECT 53.875 210.825 54.205 210.840 ;
        RECT 93.435 210.825 93.765 210.840 ;
        RECT 98.495 211.140 98.825 211.155 ;
        RECT 106.775 211.140 107.105 211.155 ;
        RECT 98.495 210.840 107.105 211.140 ;
        RECT 98.495 210.825 98.825 210.840 ;
        RECT 106.775 210.825 107.105 210.840 ;
        RECT 75.495 210.460 75.825 210.475 ;
        RECT 113.675 210.460 114.005 210.475 ;
        RECT 75.495 210.160 114.005 210.460 ;
        RECT 75.495 210.145 75.825 210.160 ;
        RECT 113.675 210.145 114.005 210.160 ;
        RECT 115.055 210.460 115.385 210.475 ;
        RECT 136.675 210.460 137.005 210.475 ;
        RECT 115.055 210.160 137.005 210.460 ;
        RECT 115.055 210.145 115.385 210.160 ;
        RECT 136.675 210.145 137.005 210.160 ;
        RECT 50.655 209.790 50.985 209.795 ;
        RECT 50.655 209.780 51.240 209.790 ;
        RECT 88.835 209.780 89.165 209.795 ;
        RECT 50.430 209.480 51.240 209.780 ;
        RECT 50.655 209.470 51.240 209.480 ;
        RECT 75.740 209.480 89.165 209.780 ;
        RECT 50.655 209.465 50.985 209.470 ;
        RECT 21.395 209.125 22.975 209.455 ;
        RECT 60.265 209.125 61.845 209.455 ;
        RECT 32.715 209.100 33.045 209.115 ;
        RECT 55.715 209.100 56.045 209.115 ;
        RECT 32.715 208.800 56.045 209.100 ;
        RECT 32.715 208.785 33.045 208.800 ;
        RECT 55.715 208.785 56.045 208.800 ;
        RECT 21.215 208.420 21.545 208.435 ;
        RECT 26.940 208.420 27.320 208.430 ;
        RECT 21.215 208.120 27.320 208.420 ;
        RECT 21.215 208.105 21.545 208.120 ;
        RECT 26.940 208.110 27.320 208.120 ;
        RECT 47.435 208.420 47.765 208.435 ;
        RECT 50.195 208.420 50.525 208.435 ;
        RECT 66.295 208.420 66.625 208.435 ;
        RECT 67.420 208.420 67.800 208.430 ;
        RECT 75.740 208.420 76.040 209.480 ;
        RECT 88.835 209.465 89.165 209.480 ;
        RECT 92.975 209.780 93.305 209.795 ;
        RECT 94.355 209.780 94.685 209.795 ;
        RECT 92.975 209.480 94.685 209.780 ;
        RECT 92.975 209.465 93.305 209.480 ;
        RECT 94.355 209.465 94.685 209.480 ;
        RECT 106.775 209.780 107.105 209.795 ;
        RECT 131.615 209.780 131.945 209.795 ;
        RECT 106.775 209.480 131.945 209.780 ;
        RECT 106.775 209.465 107.105 209.480 ;
        RECT 131.615 209.465 131.945 209.480 ;
        RECT 99.135 209.125 100.715 209.455 ;
        RECT 138.005 209.125 139.585 209.455 ;
        RECT 86.075 209.100 86.405 209.115 ;
        RECT 107.235 209.110 107.565 209.115 ;
        RECT 106.980 209.100 107.565 209.110 ;
        RECT 109.535 209.110 109.865 209.115 ;
        RECT 117.355 209.110 117.685 209.115 ;
        RECT 109.535 209.100 110.120 209.110 ;
        RECT 117.100 209.100 117.685 209.110 ;
        RECT 86.075 208.800 90.760 209.100 ;
        RECT 86.075 208.785 86.405 208.800 ;
        RECT 47.435 208.120 67.800 208.420 ;
        RECT 47.435 208.105 47.765 208.120 ;
        RECT 50.195 208.105 50.525 208.120 ;
        RECT 66.295 208.105 66.625 208.120 ;
        RECT 67.420 208.110 67.800 208.120 ;
        RECT 68.380 208.120 76.040 208.420 ;
        RECT 82.855 208.420 83.185 208.435 ;
        RECT 90.460 208.420 90.760 208.800 ;
        RECT 106.980 208.800 107.790 209.100 ;
        RECT 109.535 208.800 110.320 209.100 ;
        RECT 116.900 208.800 117.685 209.100 ;
        RECT 106.980 208.790 107.565 208.800 ;
        RECT 107.235 208.785 107.565 208.790 ;
        RECT 109.535 208.790 110.120 208.800 ;
        RECT 117.100 208.790 117.685 208.800 ;
        RECT 109.535 208.785 109.865 208.790 ;
        RECT 117.355 208.785 117.685 208.790 ;
        RECT 123.795 209.100 124.125 209.115 ;
        RECT 135.295 209.100 135.625 209.115 ;
        RECT 123.795 208.800 135.625 209.100 ;
        RECT 123.795 208.785 124.125 208.800 ;
        RECT 135.295 208.785 135.625 208.800 ;
        RECT 133.455 208.420 133.785 208.435 ;
        RECT 82.855 208.120 89.840 208.420 ;
        RECT 90.460 208.120 133.785 208.420 ;
        RECT 26.020 207.740 26.400 207.750 ;
        RECT 33.175 207.740 33.505 207.755 ;
        RECT 26.020 207.440 33.505 207.740 ;
        RECT 26.020 207.430 26.400 207.440 ;
        RECT 33.175 207.425 33.505 207.440 ;
        RECT 53.415 207.740 53.745 207.755 ;
        RECT 55.460 207.740 55.840 207.750 ;
        RECT 53.415 207.440 55.840 207.740 ;
        RECT 53.415 207.425 53.745 207.440 ;
        RECT 55.460 207.430 55.840 207.440 ;
        RECT 57.095 207.740 57.425 207.755 ;
        RECT 68.380 207.740 68.680 208.120 ;
        RECT 82.855 208.105 83.185 208.120 ;
        RECT 57.095 207.440 68.680 207.740 ;
        RECT 69.515 207.740 69.845 207.755 ;
        RECT 86.075 207.740 86.405 207.755 ;
        RECT 69.515 207.440 86.405 207.740 ;
        RECT 89.540 207.740 89.840 208.120 ;
        RECT 133.455 208.105 133.785 208.120 ;
        RECT 134.835 208.420 135.165 208.435 ;
        RECT 135.500 208.420 135.880 208.430 ;
        RECT 134.835 208.120 135.880 208.420 ;
        RECT 134.835 208.105 135.165 208.120 ;
        RECT 135.500 208.110 135.880 208.120 ;
        RECT 144.495 207.740 144.825 207.755 ;
        RECT 89.540 207.440 144.825 207.740 ;
        RECT 57.095 207.425 57.425 207.440 ;
        RECT 69.515 207.425 69.845 207.440 ;
        RECT 86.075 207.425 86.405 207.440 ;
        RECT 144.495 207.425 144.825 207.440 ;
        RECT 58.015 207.060 58.345 207.075 ;
        RECT 76.415 207.060 76.745 207.075 ;
        RECT 58.015 206.760 76.745 207.060 ;
        RECT 58.015 206.745 58.345 206.760 ;
        RECT 76.415 206.745 76.745 206.760 ;
        RECT 83.775 207.060 84.105 207.075 ;
        RECT 104.015 207.060 104.345 207.075 ;
        RECT 115.975 207.060 116.305 207.075 ;
        RECT 83.775 206.760 116.305 207.060 ;
        RECT 83.775 206.745 84.105 206.760 ;
        RECT 104.015 206.745 104.345 206.760 ;
        RECT 115.975 206.745 116.305 206.760 ;
        RECT 40.830 206.405 42.410 206.735 ;
        RECT 79.700 206.405 81.280 206.735 ;
        RECT 118.570 206.405 120.150 206.735 ;
        RECT 157.440 206.405 159.020 206.735 ;
        RECT 55.715 206.380 56.045 206.395 ;
        RECT 68.595 206.380 68.925 206.395 ;
        RECT 75.955 206.380 76.285 206.395 ;
        RECT 55.715 206.080 59.480 206.380 ;
        RECT 55.715 206.065 56.045 206.080 ;
        RECT 12.475 205.700 12.805 205.715 ;
        RECT 21.675 205.700 22.005 205.715 ;
        RECT 57.555 205.700 57.885 205.715 ;
        RECT 59.180 205.710 59.480 206.080 ;
        RECT 68.595 206.080 76.285 206.380 ;
        RECT 68.595 206.065 68.925 206.080 ;
        RECT 75.955 206.065 76.285 206.080 ;
        RECT 83.315 206.380 83.645 206.395 ;
        RECT 83.980 206.380 84.360 206.390 ;
        RECT 83.315 206.080 84.360 206.380 ;
        RECT 83.315 206.065 83.645 206.080 ;
        RECT 83.980 206.070 84.360 206.080 ;
        RECT 86.075 206.380 86.405 206.395 ;
        RECT 101.255 206.380 101.585 206.395 ;
        RECT 102.380 206.380 102.760 206.390 ;
        RECT 86.075 206.080 99.040 206.380 ;
        RECT 86.075 206.065 86.405 206.080 ;
        RECT 12.475 205.400 57.885 205.700 ;
        RECT 12.475 205.385 12.805 205.400 ;
        RECT 21.675 205.385 22.005 205.400 ;
        RECT 57.555 205.385 57.885 205.400 ;
        RECT 59.140 205.390 59.520 205.710 ;
        RECT 92.515 205.700 92.845 205.715 ;
        RECT 97.115 205.700 97.445 205.715 ;
        RECT 92.515 205.400 97.445 205.700 ;
        RECT 98.740 205.700 99.040 206.080 ;
        RECT 101.255 206.080 102.760 206.380 ;
        RECT 101.255 206.065 101.585 206.080 ;
        RECT 102.380 206.070 102.760 206.080 ;
        RECT 103.095 206.380 103.425 206.395 ;
        RECT 107.235 206.380 107.565 206.395 ;
        RECT 103.095 206.080 107.565 206.380 ;
        RECT 103.095 206.065 103.425 206.080 ;
        RECT 107.235 206.065 107.565 206.080 ;
        RECT 145.875 205.700 146.205 205.715 ;
        RECT 98.740 205.400 146.205 205.700 ;
        RECT 92.515 205.385 92.845 205.400 ;
        RECT 97.115 205.385 97.445 205.400 ;
        RECT 145.875 205.385 146.205 205.400 ;
        RECT 21.215 205.020 21.545 205.035 ;
        RECT 29.495 205.020 29.825 205.035 ;
        RECT 45.595 205.020 45.925 205.035 ;
        RECT 21.215 204.720 45.925 205.020 ;
        RECT 21.215 204.705 21.545 204.720 ;
        RECT 29.495 204.705 29.825 204.720 ;
        RECT 45.595 204.705 45.925 204.720 ;
        RECT 55.255 205.020 55.585 205.035 ;
        RECT 124.715 205.020 125.045 205.035 ;
        RECT 55.255 204.720 125.045 205.020 ;
        RECT 55.255 204.705 55.585 204.720 ;
        RECT 124.715 204.705 125.045 204.720 ;
        RECT 71.355 204.340 71.685 204.355 ;
        RECT 84.235 204.340 84.565 204.355 ;
        RECT 71.355 204.040 84.565 204.340 ;
        RECT 71.355 204.025 71.685 204.040 ;
        RECT 84.235 204.025 84.565 204.040 ;
        RECT 21.395 203.685 22.975 204.015 ;
        RECT 60.265 203.685 61.845 204.015 ;
        RECT 99.135 203.685 100.715 204.015 ;
        RECT 138.005 203.685 139.585 204.015 ;
        RECT 64.915 203.660 65.245 203.675 ;
        RECT 73.195 203.660 73.525 203.675 ;
        RECT 64.915 203.360 73.525 203.660 ;
        RECT 64.915 203.345 65.245 203.360 ;
        RECT 73.195 203.345 73.525 203.360 ;
        RECT 83.315 203.660 83.645 203.675 ;
        RECT 96.655 203.660 96.985 203.675 ;
        RECT 83.315 203.360 96.985 203.660 ;
        RECT 83.315 203.345 83.645 203.360 ;
        RECT 96.655 203.345 96.985 203.360 ;
        RECT 101.255 203.660 101.585 203.675 ;
        RECT 106.315 203.660 106.645 203.675 ;
        RECT 101.255 203.360 106.645 203.660 ;
        RECT 101.255 203.345 101.585 203.360 ;
        RECT 106.315 203.345 106.645 203.360 ;
        RECT 27.195 202.980 27.525 202.995 ;
        RECT 38.235 202.980 38.565 202.995 ;
        RECT 45.135 202.980 45.465 202.995 ;
        RECT 27.195 202.680 45.465 202.980 ;
        RECT 27.195 202.665 27.525 202.680 ;
        RECT 38.235 202.665 38.565 202.680 ;
        RECT 45.135 202.665 45.465 202.680 ;
        RECT 49.020 202.980 49.400 202.990 ;
        RECT 49.735 202.980 50.065 202.995 ;
        RECT 49.020 202.680 50.065 202.980 ;
        RECT 49.020 202.670 49.400 202.680 ;
        RECT 49.735 202.665 50.065 202.680 ;
        RECT 66.755 202.980 67.085 202.995 ;
        RECT 81.935 202.980 82.265 202.995 ;
        RECT 66.755 202.680 82.265 202.980 ;
        RECT 66.755 202.665 67.085 202.680 ;
        RECT 81.935 202.665 82.265 202.680 ;
        RECT 95.735 202.980 96.065 202.995 ;
        RECT 100.795 202.980 101.125 202.995 ;
        RECT 95.735 202.680 101.125 202.980 ;
        RECT 95.735 202.665 96.065 202.680 ;
        RECT 100.795 202.665 101.125 202.680 ;
        RECT 114.595 202.980 114.925 202.995 ;
        RECT 138.975 202.980 139.305 202.995 ;
        RECT 114.595 202.680 139.305 202.980 ;
        RECT 114.595 202.665 114.925 202.680 ;
        RECT 138.975 202.665 139.305 202.680 ;
        RECT 18.915 202.300 19.245 202.315 ;
        RECT 22.135 202.300 22.465 202.315 ;
        RECT 18.915 202.000 22.465 202.300 ;
        RECT 18.915 201.985 19.245 202.000 ;
        RECT 22.135 201.985 22.465 202.000 ;
        RECT 32.255 202.300 32.585 202.315 ;
        RECT 66.755 202.300 67.085 202.315 ;
        RECT 32.255 202.000 67.085 202.300 ;
        RECT 32.255 201.985 32.585 202.000 ;
        RECT 66.755 201.985 67.085 202.000 ;
        RECT 89.295 202.300 89.625 202.315 ;
        RECT 91.340 202.300 91.720 202.310 ;
        RECT 123.335 202.300 123.665 202.315 ;
        RECT 141.735 202.300 142.065 202.315 ;
        RECT 89.295 202.000 142.065 202.300 ;
        RECT 89.295 201.985 89.625 202.000 ;
        RECT 91.340 201.990 91.720 202.000 ;
        RECT 123.335 201.985 123.665 202.000 ;
        RECT 141.735 201.985 142.065 202.000 ;
        RECT 13.395 201.620 13.725 201.635 ;
        RECT 19.835 201.620 20.165 201.635 ;
        RECT 13.395 201.320 20.165 201.620 ;
        RECT 13.395 201.305 13.725 201.320 ;
        RECT 19.835 201.305 20.165 201.320 ;
        RECT 42.835 201.620 43.165 201.635 ;
        RECT 54.335 201.620 54.665 201.635 ;
        RECT 42.835 201.320 54.665 201.620 ;
        RECT 42.835 201.305 43.165 201.320 ;
        RECT 54.335 201.305 54.665 201.320 ;
        RECT 58.935 201.620 59.265 201.635 ;
        RECT 73.195 201.620 73.525 201.635 ;
        RECT 58.935 201.320 73.525 201.620 ;
        RECT 58.935 201.305 59.265 201.320 ;
        RECT 73.195 201.305 73.525 201.320 ;
        RECT 82.855 201.620 83.185 201.635 ;
        RECT 93.180 201.620 93.560 201.630 ;
        RECT 94.815 201.620 95.145 201.635 ;
        RECT 82.855 201.320 95.145 201.620 ;
        RECT 82.855 201.305 83.185 201.320 ;
        RECT 93.180 201.310 93.560 201.320 ;
        RECT 94.815 201.305 95.145 201.320 ;
        RECT 97.115 201.620 97.445 201.635 ;
        RECT 113.215 201.620 113.545 201.635 ;
        RECT 97.115 201.320 113.545 201.620 ;
        RECT 97.115 201.305 97.445 201.320 ;
        RECT 113.215 201.305 113.545 201.320 ;
        RECT 40.830 200.965 42.410 201.295 ;
        RECT 79.700 200.965 81.280 201.295 ;
        RECT 118.570 200.965 120.150 201.295 ;
        RECT 157.440 200.965 159.020 201.295 ;
        RECT 50.655 200.940 50.985 200.955 ;
        RECT 43.540 200.640 50.985 200.940 ;
        RECT 40.535 200.260 40.865 200.275 ;
        RECT 43.540 200.260 43.840 200.640 ;
        RECT 50.655 200.625 50.985 200.640 ;
        RECT 55.715 200.940 56.045 200.955 ;
        RECT 59.855 200.940 60.185 200.955 ;
        RECT 55.715 200.640 60.185 200.940 ;
        RECT 55.715 200.625 56.045 200.640 ;
        RECT 59.855 200.625 60.185 200.640 ;
        RECT 82.855 200.940 83.185 200.955 ;
        RECT 94.815 200.940 95.145 200.955 ;
        RECT 82.855 200.640 95.145 200.940 ;
        RECT 82.855 200.625 83.185 200.640 ;
        RECT 94.815 200.625 95.145 200.640 ;
        RECT 97.115 200.940 97.445 200.955 ;
        RECT 117.815 200.940 118.145 200.955 ;
        RECT 97.115 200.640 118.145 200.940 ;
        RECT 97.115 200.625 97.445 200.640 ;
        RECT 117.815 200.625 118.145 200.640 ;
        RECT 121.495 200.940 121.825 200.955 ;
        RECT 150.935 200.940 151.265 200.955 ;
        RECT 121.495 200.640 151.265 200.940 ;
        RECT 121.495 200.625 121.825 200.640 ;
        RECT 150.935 200.625 151.265 200.640 ;
        RECT 40.535 199.960 43.840 200.260 ;
        RECT 50.655 200.260 50.985 200.275 ;
        RECT 56.175 200.260 56.505 200.275 ;
        RECT 50.655 199.960 56.505 200.260 ;
        RECT 40.535 199.945 40.865 199.960 ;
        RECT 50.655 199.945 50.985 199.960 ;
        RECT 56.175 199.945 56.505 199.960 ;
        RECT 67.675 200.260 68.005 200.275 ;
        RECT 78.255 200.260 78.585 200.275 ;
        RECT 67.675 199.960 78.585 200.260 ;
        RECT 67.675 199.945 68.005 199.960 ;
        RECT 78.255 199.945 78.585 199.960 ;
        RECT 83.775 200.260 84.105 200.275 ;
        RECT 88.835 200.260 89.165 200.275 ;
        RECT 124.255 200.260 124.585 200.275 ;
        RECT 83.775 199.960 124.585 200.260 ;
        RECT 83.775 199.945 84.105 199.960 ;
        RECT 88.835 199.945 89.165 199.960 ;
        RECT 124.255 199.945 124.585 199.960 ;
        RECT 27.195 199.580 27.525 199.595 ;
        RECT 70.435 199.580 70.765 199.595 ;
        RECT 92.515 199.580 92.845 199.595 ;
        RECT 96.655 199.580 96.985 199.595 ;
        RECT 106.775 199.580 107.105 199.595 ;
        RECT 108.155 199.580 108.485 199.595 ;
        RECT 27.195 199.280 88.920 199.580 ;
        RECT 27.195 199.265 27.525 199.280 ;
        RECT 70.435 199.265 70.765 199.280 ;
        RECT 39.155 198.900 39.485 198.915 ;
        RECT 54.795 198.900 55.125 198.915 ;
        RECT 39.155 198.600 55.125 198.900 ;
        RECT 88.620 198.900 88.920 199.280 ;
        RECT 92.515 199.280 96.985 199.580 ;
        RECT 92.515 199.265 92.845 199.280 ;
        RECT 96.655 199.265 96.985 199.280 ;
        RECT 97.820 199.280 108.485 199.580 ;
        RECT 97.820 198.900 98.120 199.280 ;
        RECT 106.775 199.265 107.105 199.280 ;
        RECT 108.155 199.265 108.485 199.280 ;
        RECT 116.435 199.580 116.765 199.595 ;
        RECT 132.995 199.580 133.325 199.595 ;
        RECT 116.435 199.280 133.325 199.580 ;
        RECT 116.435 199.265 116.765 199.280 ;
        RECT 132.995 199.265 133.325 199.280 ;
        RECT 88.620 198.600 98.120 198.900 ;
        RECT 102.635 198.900 102.965 198.915 ;
        RECT 121.035 198.900 121.365 198.915 ;
        RECT 102.635 198.600 121.365 198.900 ;
        RECT 39.155 198.585 39.485 198.600 ;
        RECT 54.795 198.585 55.125 198.600 ;
        RECT 102.635 198.585 102.965 198.600 ;
        RECT 121.035 198.585 121.365 198.600 ;
        RECT 21.395 198.245 22.975 198.575 ;
        RECT 60.265 198.245 61.845 198.575 ;
        RECT 99.135 198.245 100.715 198.575 ;
        RECT 138.005 198.245 139.585 198.575 ;
        RECT 46.055 198.220 46.385 198.235 ;
        RECT 52.495 198.220 52.825 198.235 ;
        RECT 46.055 197.920 52.825 198.220 ;
        RECT 46.055 197.905 46.385 197.920 ;
        RECT 52.495 197.905 52.825 197.920 ;
        RECT 73.195 198.220 73.525 198.235 ;
        RECT 76.415 198.220 76.745 198.235 ;
        RECT 85.615 198.230 85.945 198.235 ;
        RECT 85.615 198.220 86.200 198.230 ;
        RECT 73.195 197.920 86.200 198.220 ;
        RECT 73.195 197.905 73.525 197.920 ;
        RECT 76.415 197.905 76.745 197.920 ;
        RECT 85.615 197.910 86.200 197.920 ;
        RECT 85.615 197.905 85.945 197.910 ;
        RECT 90.675 197.905 91.005 198.235 ;
        RECT 101.255 198.220 101.585 198.235 ;
        RECT 124.255 198.220 124.585 198.235 ;
        RECT 101.255 197.920 124.585 198.220 ;
        RECT 101.255 197.905 101.585 197.920 ;
        RECT 124.255 197.905 124.585 197.920 ;
        RECT 25.355 197.540 25.685 197.555 ;
        RECT 53.620 197.540 54.000 197.550 ;
        RECT 54.335 197.540 54.665 197.555 ;
        RECT 25.355 197.240 54.665 197.540 ;
        RECT 25.355 197.225 25.685 197.240 ;
        RECT 53.620 197.230 54.000 197.240 ;
        RECT 54.335 197.225 54.665 197.240 ;
        RECT 86.075 197.540 86.405 197.555 ;
        RECT 90.690 197.540 90.990 197.905 ;
        RECT 98.035 197.550 98.365 197.555 ;
        RECT 97.780 197.540 98.365 197.550 ;
        RECT 86.075 197.240 90.990 197.540 ;
        RECT 97.580 197.240 98.365 197.540 ;
        RECT 86.075 197.225 86.405 197.240 ;
        RECT 97.780 197.230 98.365 197.240 ;
        RECT 98.035 197.225 98.365 197.230 ;
        RECT 99.415 197.540 99.745 197.555 ;
        RECT 120.115 197.540 120.445 197.555 ;
        RECT 99.415 197.240 120.445 197.540 ;
        RECT 99.415 197.225 99.745 197.240 ;
        RECT 120.115 197.225 120.445 197.240 ;
        RECT 42.375 196.860 42.705 196.875 ;
        RECT 59.855 196.860 60.185 196.875 ;
        RECT 103.095 196.860 103.425 196.875 ;
        RECT 111.375 196.860 111.705 196.875 ;
        RECT 112.755 196.860 113.085 196.875 ;
        RECT 131.155 196.860 131.485 196.875 ;
        RECT 42.375 196.560 59.480 196.860 ;
        RECT 42.375 196.545 42.705 196.560 ;
        RECT 46.515 196.180 46.845 196.195 ;
        RECT 54.795 196.180 55.125 196.195 ;
        RECT 46.515 195.880 55.125 196.180 ;
        RECT 59.180 196.180 59.480 196.560 ;
        RECT 59.855 196.560 103.425 196.860 ;
        RECT 59.855 196.545 60.185 196.560 ;
        RECT 103.095 196.545 103.425 196.560 ;
        RECT 104.030 196.560 111.705 196.860 ;
        RECT 59.855 196.180 60.185 196.195 ;
        RECT 59.180 195.880 60.185 196.180 ;
        RECT 46.515 195.865 46.845 195.880 ;
        RECT 54.795 195.865 55.125 195.880 ;
        RECT 59.855 195.865 60.185 195.880 ;
        RECT 92.055 196.180 92.385 196.195 ;
        RECT 94.355 196.180 94.685 196.195 ;
        RECT 104.030 196.180 104.330 196.560 ;
        RECT 111.375 196.545 111.705 196.560 ;
        RECT 112.540 196.560 131.485 196.860 ;
        RECT 112.540 196.545 113.085 196.560 ;
        RECT 131.155 196.545 131.485 196.560 ;
        RECT 92.055 195.880 104.330 196.180 ;
        RECT 104.935 196.180 105.265 196.195 ;
        RECT 112.540 196.180 112.840 196.545 ;
        RECT 104.935 195.880 112.840 196.180 ;
        RECT 126.555 196.180 126.885 196.195 ;
        RECT 134.835 196.180 135.165 196.195 ;
        RECT 126.555 195.880 135.165 196.180 ;
        RECT 92.055 195.865 92.385 195.880 ;
        RECT 94.355 195.865 94.685 195.880 ;
        RECT 104.935 195.865 105.265 195.880 ;
        RECT 126.555 195.865 126.885 195.880 ;
        RECT 134.835 195.865 135.165 195.880 ;
        RECT 40.830 195.525 42.410 195.855 ;
        RECT 79.700 195.525 81.280 195.855 ;
        RECT 118.570 195.525 120.150 195.855 ;
        RECT 157.440 195.525 159.020 195.855 ;
        RECT 46.975 195.500 47.305 195.515 ;
        RECT 48.100 195.500 48.480 195.510 ;
        RECT 46.975 195.200 48.480 195.500 ;
        RECT 46.975 195.185 47.305 195.200 ;
        RECT 48.100 195.190 48.480 195.200 ;
        RECT 82.395 195.500 82.725 195.515 ;
        RECT 87.455 195.500 87.785 195.515 ;
        RECT 111.375 195.500 111.705 195.515 ;
        RECT 82.395 195.200 111.705 195.500 ;
        RECT 82.395 195.185 82.725 195.200 ;
        RECT 87.455 195.185 87.785 195.200 ;
        RECT 111.375 195.185 111.705 195.200 ;
        RECT 120.575 195.500 120.905 195.515 ;
        RECT 126.095 195.500 126.425 195.515 ;
        RECT 120.575 195.200 126.425 195.500 ;
        RECT 120.575 195.185 120.905 195.200 ;
        RECT 126.095 195.185 126.425 195.200 ;
        RECT 33.175 194.820 33.505 194.835 ;
        RECT 52.955 194.820 53.285 194.835 ;
        RECT 33.175 194.520 53.285 194.820 ;
        RECT 33.175 194.505 33.505 194.520 ;
        RECT 52.955 194.505 53.285 194.520 ;
        RECT 58.935 194.820 59.265 194.835 ;
        RECT 67.675 194.820 68.005 194.835 ;
        RECT 58.935 194.520 68.005 194.820 ;
        RECT 58.935 194.505 59.265 194.520 ;
        RECT 67.675 194.505 68.005 194.520 ;
        RECT 82.855 194.820 83.185 194.835 ;
        RECT 143.575 194.820 143.905 194.835 ;
        RECT 82.855 194.520 143.905 194.820 ;
        RECT 82.855 194.505 83.185 194.520 ;
        RECT 143.575 194.505 143.905 194.520 ;
        RECT 60.315 194.140 60.645 194.155 ;
        RECT 84.695 194.140 85.025 194.155 ;
        RECT 60.315 193.840 85.025 194.140 ;
        RECT 60.315 193.825 60.645 193.840 ;
        RECT 84.695 193.825 85.025 193.840 ;
        RECT 106.315 194.140 106.645 194.155 ;
        RECT 106.980 194.140 107.360 194.150 ;
        RECT 106.315 193.840 107.360 194.140 ;
        RECT 106.315 193.825 106.645 193.840 ;
        RECT 106.980 193.830 107.360 193.840 ;
        RECT 109.535 194.140 109.865 194.155 ;
        RECT 119.655 194.140 119.985 194.155 ;
        RECT 109.535 193.840 119.985 194.140 ;
        RECT 109.535 193.825 109.865 193.840 ;
        RECT 119.655 193.825 119.985 193.840 ;
        RECT 42.375 193.460 42.705 193.475 ;
        RECT 53.415 193.460 53.745 193.475 ;
        RECT 42.375 193.160 53.745 193.460 ;
        RECT 42.375 193.145 42.705 193.160 ;
        RECT 53.415 193.145 53.745 193.160 ;
        RECT 67.420 193.460 67.800 193.470 ;
        RECT 72.275 193.460 72.605 193.475 ;
        RECT 67.420 193.160 72.605 193.460 ;
        RECT 67.420 193.150 67.800 193.160 ;
        RECT 72.275 193.145 72.605 193.160 ;
        RECT 83.315 193.460 83.645 193.475 ;
        RECT 89.295 193.460 89.625 193.475 ;
        RECT 83.315 193.160 89.625 193.460 ;
        RECT 83.315 193.145 83.645 193.160 ;
        RECT 89.295 193.145 89.625 193.160 ;
        RECT 107.695 193.460 108.025 193.475 ;
        RECT 131.615 193.460 131.945 193.475 ;
        RECT 107.695 193.160 131.945 193.460 ;
        RECT 107.695 193.145 108.025 193.160 ;
        RECT 131.615 193.145 131.945 193.160 ;
        RECT 21.395 192.805 22.975 193.135 ;
        RECT 60.265 192.805 61.845 193.135 ;
        RECT 99.135 192.805 100.715 193.135 ;
        RECT 138.005 192.805 139.585 193.135 ;
        RECT 94.100 192.780 94.480 192.790 ;
        RECT 98.035 192.780 98.365 192.795 ;
        RECT 72.980 192.480 98.365 192.780 ;
        RECT 26.735 192.100 27.065 192.115 ;
        RECT 52.035 192.100 52.365 192.115 ;
        RECT 26.735 191.800 52.365 192.100 ;
        RECT 26.735 191.785 27.065 191.800 ;
        RECT 52.035 191.785 52.365 191.800 ;
        RECT 58.015 192.100 58.345 192.115 ;
        RECT 72.980 192.100 73.280 192.480 ;
        RECT 94.100 192.470 94.480 192.480 ;
        RECT 98.035 192.465 98.365 192.480 ;
        RECT 102.175 192.780 102.505 192.795 ;
        RECT 135.295 192.780 135.625 192.795 ;
        RECT 102.175 192.480 135.625 192.780 ;
        RECT 102.175 192.465 102.505 192.480 ;
        RECT 135.295 192.465 135.625 192.480 ;
        RECT 58.015 191.800 73.280 192.100 ;
        RECT 73.655 192.100 73.985 192.115 ;
        RECT 127.475 192.100 127.805 192.115 ;
        RECT 73.655 191.800 127.805 192.100 ;
        RECT 58.015 191.785 58.345 191.800 ;
        RECT 73.655 191.785 73.985 191.800 ;
        RECT 127.475 191.785 127.805 191.800 ;
        RECT 74.575 191.420 74.905 191.435 ;
        RECT 103.555 191.420 103.885 191.435 ;
        RECT 154.820 191.420 155.200 191.430 ;
        RECT 74.575 191.120 87.310 191.420 ;
        RECT 74.575 191.105 74.905 191.120 ;
        RECT 87.010 190.755 87.310 191.120 ;
        RECT 103.555 191.120 155.200 191.420 ;
        RECT 103.555 191.105 103.885 191.120 ;
        RECT 154.820 191.110 155.200 191.120 ;
        RECT 86.995 190.740 87.325 190.755 ;
        RECT 105.855 190.740 106.185 190.755 ;
        RECT 86.995 190.440 106.185 190.740 ;
        RECT 86.995 190.425 87.325 190.440 ;
        RECT 105.855 190.425 106.185 190.440 ;
        RECT 107.695 190.740 108.025 190.755 ;
        RECT 117.815 190.740 118.145 190.755 ;
        RECT 107.695 190.440 118.145 190.740 ;
        RECT 107.695 190.425 108.025 190.440 ;
        RECT 117.815 190.425 118.145 190.440 ;
        RECT 40.830 190.085 42.410 190.415 ;
        RECT 79.700 190.085 81.280 190.415 ;
        RECT 118.570 190.085 120.150 190.415 ;
        RECT 157.440 190.085 159.020 190.415 ;
        RECT 85.615 190.060 85.945 190.075 ;
        RECT 86.995 190.060 87.325 190.075 ;
        RECT 85.615 189.760 87.325 190.060 ;
        RECT 85.615 189.745 85.945 189.760 ;
        RECT 86.995 189.745 87.325 189.760 ;
        RECT 88.835 190.060 89.165 190.075 ;
        RECT 100.335 190.060 100.665 190.075 ;
        RECT 88.835 189.760 100.665 190.060 ;
        RECT 88.835 189.745 89.165 189.760 ;
        RECT 100.335 189.745 100.665 189.760 ;
        RECT 101.715 190.060 102.045 190.075 ;
        RECT 116.895 190.060 117.225 190.075 ;
        RECT 101.715 189.760 117.225 190.060 ;
        RECT 101.715 189.745 102.045 189.760 ;
        RECT 116.895 189.745 117.225 189.760 ;
        RECT 132.075 190.060 132.405 190.075 ;
        RECT 138.515 190.060 138.845 190.075 ;
        RECT 132.075 189.760 138.845 190.060 ;
        RECT 132.075 189.745 132.405 189.760 ;
        RECT 138.515 189.745 138.845 189.760 ;
        RECT 48.355 189.380 48.685 189.395 ;
        RECT 78.715 189.380 79.045 189.395 ;
        RECT 97.575 189.380 97.905 189.395 ;
        RECT 116.895 189.390 117.225 189.395 ;
        RECT 116.895 189.380 117.480 189.390 ;
        RECT 148.635 189.380 148.965 189.395 ;
        RECT 48.355 189.080 50.050 189.380 ;
        RECT 48.355 189.065 48.685 189.080 ;
        RECT 49.750 188.715 50.050 189.080 ;
        RECT 78.715 189.080 115.370 189.380 ;
        RECT 116.690 189.080 148.965 189.380 ;
        RECT 78.715 189.065 79.045 189.080 ;
        RECT 97.575 189.065 97.905 189.080 ;
        RECT 49.735 188.385 50.065 188.715 ;
        RECT 73.655 188.700 73.985 188.715 ;
        RECT 114.135 188.700 114.465 188.715 ;
        RECT 73.655 188.400 114.465 188.700 ;
        RECT 115.070 188.700 115.370 189.080 ;
        RECT 116.895 189.070 117.480 189.080 ;
        RECT 116.895 189.065 117.225 189.070 ;
        RECT 148.635 189.065 148.965 189.080 ;
        RECT 126.555 188.700 126.885 188.715 ;
        RECT 115.070 188.400 126.885 188.700 ;
        RECT 73.655 188.385 73.985 188.400 ;
        RECT 114.135 188.385 114.465 188.400 ;
        RECT 126.555 188.385 126.885 188.400 ;
        RECT 83.980 188.020 84.360 188.030 ;
        RECT 84.695 188.020 85.025 188.035 ;
        RECT 94.100 188.020 94.480 188.030 ;
        RECT 94.815 188.020 95.145 188.035 ;
        RECT 83.980 187.720 89.840 188.020 ;
        RECT 83.980 187.710 84.360 187.720 ;
        RECT 84.695 187.705 85.025 187.720 ;
        RECT 21.395 187.365 22.975 187.695 ;
        RECT 60.265 187.365 61.845 187.695 ;
        RECT 39.820 187.340 40.200 187.350 ;
        RECT 41.915 187.340 42.245 187.355 ;
        RECT 39.820 187.040 42.245 187.340 ;
        RECT 39.820 187.030 40.200 187.040 ;
        RECT 41.915 187.025 42.245 187.040 ;
        RECT 42.835 187.340 43.165 187.355 ;
        RECT 46.515 187.340 46.845 187.355 ;
        RECT 55.255 187.340 55.585 187.355 ;
        RECT 42.835 187.040 55.585 187.340 ;
        RECT 89.540 187.340 89.840 187.720 ;
        RECT 94.100 187.720 95.145 188.020 ;
        RECT 94.100 187.710 94.480 187.720 ;
        RECT 94.815 187.705 95.145 187.720 ;
        RECT 103.095 188.020 103.425 188.035 ;
        RECT 121.035 188.020 121.365 188.035 ;
        RECT 103.095 187.720 121.365 188.020 ;
        RECT 103.095 187.705 103.425 187.720 ;
        RECT 121.035 187.705 121.365 187.720 ;
        RECT 122.415 188.020 122.745 188.035 ;
        RECT 130.235 188.020 130.565 188.035 ;
        RECT 122.415 187.720 130.565 188.020 ;
        RECT 122.415 187.705 122.745 187.720 ;
        RECT 130.235 187.705 130.565 187.720 ;
        RECT 99.135 187.365 100.715 187.695 ;
        RECT 138.005 187.365 139.585 187.695 ;
        RECT 102.635 187.340 102.965 187.355 ;
        RECT 129.315 187.340 129.645 187.355 ;
        RECT 89.540 187.040 98.120 187.340 ;
        RECT 42.835 187.025 43.165 187.040 ;
        RECT 46.515 187.025 46.845 187.040 ;
        RECT 55.255 187.025 55.585 187.040 ;
        RECT 54.795 186.660 55.125 186.675 ;
        RECT 93.435 186.660 93.765 186.675 ;
        RECT 97.820 186.670 98.120 187.040 ;
        RECT 101.500 187.040 129.645 187.340 ;
        RECT 54.795 186.360 93.765 186.660 ;
        RECT 54.795 186.345 55.125 186.360 ;
        RECT 93.435 186.345 93.765 186.360 ;
        RECT 97.780 186.660 98.160 186.670 ;
        RECT 101.500 186.660 101.800 187.040 ;
        RECT 102.635 187.025 102.965 187.040 ;
        RECT 129.315 187.025 129.645 187.040 ;
        RECT 109.995 186.670 110.325 186.675 ;
        RECT 97.780 186.360 101.800 186.660 ;
        RECT 109.740 186.660 110.325 186.670 ;
        RECT 114.135 186.660 114.465 186.675 ;
        RECT 128.395 186.660 128.725 186.675 ;
        RECT 109.740 186.360 110.550 186.660 ;
        RECT 114.135 186.360 128.725 186.660 ;
        RECT 97.780 186.350 98.160 186.360 ;
        RECT 109.740 186.350 110.325 186.360 ;
        RECT 109.995 186.345 110.325 186.350 ;
        RECT 114.135 186.345 114.465 186.360 ;
        RECT 128.395 186.345 128.725 186.360 ;
        RECT 44.675 185.980 45.005 185.995 ;
        RECT 49.020 185.980 49.400 185.990 ;
        RECT 53.875 185.980 54.205 185.995 ;
        RECT 44.675 185.680 54.205 185.980 ;
        RECT 44.675 185.665 45.005 185.680 ;
        RECT 49.020 185.670 49.400 185.680 ;
        RECT 53.875 185.665 54.205 185.680 ;
        RECT 59.395 185.980 59.725 185.995 ;
        RECT 62.615 185.980 62.945 185.995 ;
        RECT 59.395 185.680 62.945 185.980 ;
        RECT 59.395 185.665 59.725 185.680 ;
        RECT 62.615 185.665 62.945 185.680 ;
        RECT 84.695 185.980 85.025 185.995 ;
        RECT 103.555 185.980 103.885 185.995 ;
        RECT 124.255 185.980 124.585 185.995 ;
        RECT 84.695 185.680 103.885 185.980 ;
        RECT 84.695 185.665 85.025 185.680 ;
        RECT 103.555 185.665 103.885 185.680 ;
        RECT 104.260 185.680 124.585 185.980 ;
        RECT 48.815 185.300 49.145 185.315 ;
        RECT 57.555 185.300 57.885 185.315 ;
        RECT 48.815 185.000 57.885 185.300 ;
        RECT 48.815 184.985 49.145 185.000 ;
        RECT 57.555 184.985 57.885 185.000 ;
        RECT 93.180 185.300 93.560 185.310 ;
        RECT 99.415 185.300 99.745 185.315 ;
        RECT 104.260 185.300 104.560 185.680 ;
        RECT 124.255 185.665 124.585 185.680 ;
        RECT 93.180 185.000 104.560 185.300 ;
        RECT 121.035 185.300 121.365 185.315 ;
        RECT 135.755 185.300 136.085 185.315 ;
        RECT 121.035 185.000 136.085 185.300 ;
        RECT 93.180 184.990 93.560 185.000 ;
        RECT 99.415 184.985 99.745 185.000 ;
        RECT 121.035 184.985 121.365 185.000 ;
        RECT 135.755 184.985 136.085 185.000 ;
        RECT 40.830 184.645 42.410 184.975 ;
        RECT 79.700 184.645 81.280 184.975 ;
        RECT 118.570 184.645 120.150 184.975 ;
        RECT 157.440 184.645 159.020 184.975 ;
        RECT 91.340 184.620 91.720 184.630 ;
        RECT 95.275 184.620 95.605 184.635 ;
        RECT 91.340 184.320 95.605 184.620 ;
        RECT 91.340 184.310 91.720 184.320 ;
        RECT 95.275 184.305 95.605 184.320 ;
        RECT 97.575 184.620 97.905 184.635 ;
        RECT 97.575 184.320 116.520 184.620 ;
        RECT 97.575 184.305 97.905 184.320 ;
        RECT 116.220 183.955 116.520 184.320 ;
        RECT 86.075 183.940 86.405 183.955 ;
        RECT 97.575 183.940 97.905 183.955 ;
        RECT 86.075 183.640 97.905 183.940 ;
        RECT 86.075 183.625 86.405 183.640 ;
        RECT 97.575 183.625 97.905 183.640 ;
        RECT 98.495 183.940 98.825 183.955 ;
        RECT 113.675 183.940 114.005 183.955 ;
        RECT 98.495 183.640 114.005 183.940 ;
        RECT 116.220 183.940 116.765 183.955 ;
        RECT 150.475 183.940 150.805 183.955 ;
        RECT 116.220 183.640 150.805 183.940 ;
        RECT 98.495 183.625 98.825 183.640 ;
        RECT 113.675 183.625 114.005 183.640 ;
        RECT 116.435 183.625 116.765 183.640 ;
        RECT 150.475 183.625 150.805 183.640 ;
        RECT 49.735 183.260 50.065 183.275 ;
        RECT 63.535 183.260 63.865 183.275 ;
        RECT 49.735 182.960 63.865 183.260 ;
        RECT 49.735 182.945 50.065 182.960 ;
        RECT 63.535 182.945 63.865 182.960 ;
        RECT 92.055 183.260 92.385 183.275 ;
        RECT 109.075 183.260 109.405 183.275 ;
        RECT 92.055 182.960 109.405 183.260 ;
        RECT 92.055 182.945 92.385 182.960 ;
        RECT 109.075 182.945 109.405 182.960 ;
        RECT 126.095 183.260 126.425 183.275 ;
        RECT 142.195 183.260 142.525 183.275 ;
        RECT 126.095 182.960 142.525 183.260 ;
        RECT 126.095 182.945 126.425 182.960 ;
        RECT 142.195 182.945 142.525 182.960 ;
        RECT 70.435 182.580 70.765 182.595 ;
        RECT 88.835 182.580 89.165 182.595 ;
        RECT 98.495 182.580 98.825 182.595 ;
        RECT 70.435 182.280 98.825 182.580 ;
        RECT 109.090 182.580 109.390 182.945 ;
        RECT 132.075 182.580 132.405 182.595 ;
        RECT 109.090 182.280 132.405 182.580 ;
        RECT 70.435 182.265 70.765 182.280 ;
        RECT 88.835 182.265 89.165 182.280 ;
        RECT 98.495 182.265 98.825 182.280 ;
        RECT 132.075 182.265 132.405 182.280 ;
        RECT 21.395 181.925 22.975 182.255 ;
        RECT 60.265 181.925 61.845 182.255 ;
        RECT 99.135 181.925 100.715 182.255 ;
        RECT 138.005 181.925 139.585 182.255 ;
        RECT 85.820 181.900 86.200 181.910 ;
        RECT 88.835 181.900 89.165 181.915 ;
        RECT 109.995 181.900 110.325 181.915 ;
        RECT 85.820 181.600 89.165 181.900 ;
        RECT 85.820 181.590 86.200 181.600 ;
        RECT 88.835 181.585 89.165 181.600 ;
        RECT 105.870 181.600 110.325 181.900 ;
        RECT 42.835 181.220 43.165 181.235 ;
        RECT 44.420 181.220 44.800 181.230 ;
        RECT 50.655 181.220 50.985 181.235 ;
        RECT 42.835 180.920 50.985 181.220 ;
        RECT 42.835 180.905 43.165 180.920 ;
        RECT 44.420 180.910 44.800 180.920 ;
        RECT 50.655 180.905 50.985 180.920 ;
        RECT 56.175 181.220 56.505 181.235 ;
        RECT 91.135 181.220 91.465 181.235 ;
        RECT 56.175 180.920 91.465 181.220 ;
        RECT 56.175 180.905 56.505 180.920 ;
        RECT 91.135 180.905 91.465 180.920 ;
        RECT 38.235 180.540 38.565 180.555 ;
        RECT 49.735 180.540 50.065 180.555 ;
        RECT 52.495 180.540 52.825 180.555 ;
        RECT 38.235 180.240 48.440 180.540 ;
        RECT 38.235 180.225 38.565 180.240 ;
        RECT 48.140 179.860 48.440 180.240 ;
        RECT 49.735 180.240 52.825 180.540 ;
        RECT 49.735 180.225 50.065 180.240 ;
        RECT 52.495 180.225 52.825 180.240 ;
        RECT 53.875 180.540 54.205 180.555 ;
        RECT 59.395 180.540 59.725 180.555 ;
        RECT 53.875 180.240 59.725 180.540 ;
        RECT 53.875 180.225 54.205 180.240 ;
        RECT 59.395 180.225 59.725 180.240 ;
        RECT 82.395 180.540 82.725 180.555 ;
        RECT 105.870 180.540 106.170 181.600 ;
        RECT 109.995 181.585 110.325 181.600 ;
        RECT 119.655 181.900 119.985 181.915 ;
        RECT 134.835 181.900 135.165 181.915 ;
        RECT 119.655 181.600 135.165 181.900 ;
        RECT 119.655 181.585 119.985 181.600 ;
        RECT 134.835 181.585 135.165 181.600 ;
        RECT 109.995 181.220 110.325 181.235 ;
        RECT 132.535 181.220 132.865 181.235 ;
        RECT 109.995 180.920 132.865 181.220 ;
        RECT 109.995 180.905 110.325 180.920 ;
        RECT 132.535 180.905 132.865 180.920 ;
        RECT 82.395 180.240 106.170 180.540 ;
        RECT 111.375 180.540 111.705 180.555 ;
        RECT 121.955 180.540 122.285 180.555 ;
        RECT 111.375 180.240 122.285 180.540 ;
        RECT 82.395 180.225 82.725 180.240 ;
        RECT 111.375 180.225 111.705 180.240 ;
        RECT 121.955 180.225 122.285 180.240 ;
        RECT 126.555 180.540 126.885 180.555 ;
        RECT 143.115 180.540 143.445 180.555 ;
        RECT 126.555 180.240 143.445 180.540 ;
        RECT 126.555 180.225 126.885 180.240 ;
        RECT 143.115 180.225 143.445 180.240 ;
        RECT 49.735 179.860 50.065 179.875 ;
        RECT 48.140 179.560 50.065 179.860 ;
        RECT 49.735 179.545 50.065 179.560 ;
        RECT 56.635 179.860 56.965 179.875 ;
        RECT 58.935 179.860 59.265 179.875 ;
        RECT 88.835 179.870 89.165 179.875 ;
        RECT 56.635 179.560 59.265 179.860 ;
        RECT 56.635 179.545 56.965 179.560 ;
        RECT 58.935 179.545 59.265 179.560 ;
        RECT 88.580 179.860 89.165 179.870 ;
        RECT 88.580 179.560 110.540 179.860 ;
        RECT 88.580 179.550 89.165 179.560 ;
        RECT 88.835 179.545 89.165 179.550 ;
        RECT 40.830 179.205 42.410 179.535 ;
        RECT 79.700 179.205 81.280 179.535 ;
        RECT 48.100 178.500 48.480 178.510 ;
        RECT 98.495 178.500 98.825 178.515 ;
        RECT 48.100 178.200 98.825 178.500 ;
        RECT 110.240 178.500 110.540 179.560 ;
        RECT 118.570 179.205 120.150 179.535 ;
        RECT 157.440 179.205 159.020 179.535 ;
        RECT 112.755 178.500 113.085 178.515 ;
        RECT 137.135 178.500 137.465 178.515 ;
        RECT 110.240 178.200 137.465 178.500 ;
        RECT 48.100 178.190 48.480 178.200 ;
        RECT 98.495 178.185 98.825 178.200 ;
        RECT 112.755 178.185 113.085 178.200 ;
        RECT 137.135 178.185 137.465 178.200 ;
        RECT 41.915 177.820 42.245 177.835 ;
        RECT 50.655 177.820 50.985 177.835 ;
        RECT 41.915 177.520 50.985 177.820 ;
        RECT 41.915 177.505 42.245 177.520 ;
        RECT 50.655 177.505 50.985 177.520 ;
        RECT 58.935 177.820 59.265 177.835 ;
        RECT 73.655 177.820 73.985 177.835 ;
        RECT 58.935 177.520 73.985 177.820 ;
        RECT 58.935 177.505 59.265 177.520 ;
        RECT 73.655 177.505 73.985 177.520 ;
        RECT 84.695 177.820 85.025 177.835 ;
        RECT 121.495 177.820 121.825 177.835 ;
        RECT 135.295 177.820 135.625 177.835 ;
        RECT 84.695 177.520 135.625 177.820 ;
        RECT 84.695 177.505 85.025 177.520 ;
        RECT 121.495 177.505 121.825 177.520 ;
        RECT 135.295 177.505 135.625 177.520 ;
        RECT 40.535 177.140 40.865 177.155 ;
        RECT 52.495 177.140 52.825 177.155 ;
        RECT 40.535 176.840 52.825 177.140 ;
        RECT 40.535 176.825 40.865 176.840 ;
        RECT 52.495 176.825 52.825 176.840 ;
        RECT 86.995 177.140 87.325 177.155 ;
        RECT 89.755 177.140 90.085 177.155 ;
        RECT 86.995 176.840 90.085 177.140 ;
        RECT 86.995 176.825 87.325 176.840 ;
        RECT 89.755 176.825 90.085 176.840 ;
        RECT 101.255 177.140 101.585 177.155 ;
        RECT 109.995 177.140 110.325 177.155 ;
        RECT 101.255 176.840 110.325 177.140 ;
        RECT 101.255 176.825 101.585 176.840 ;
        RECT 109.995 176.825 110.325 176.840 ;
        RECT 21.395 176.485 22.975 176.815 ;
        RECT 60.265 176.485 61.845 176.815 ;
        RECT 99.135 176.485 100.715 176.815 ;
        RECT 138.005 176.485 139.585 176.815 ;
        RECT 84.235 176.460 84.565 176.475 ;
        RECT 92.055 176.460 92.385 176.475 ;
        RECT 84.235 176.160 92.385 176.460 ;
        RECT 84.235 176.145 84.565 176.160 ;
        RECT 92.055 176.145 92.385 176.160 ;
        RECT 25.815 175.780 26.145 175.795 ;
        RECT 54.335 175.780 54.665 175.795 ;
        RECT 96.195 175.780 96.525 175.795 ;
        RECT 25.815 175.480 54.665 175.780 ;
        RECT 25.815 175.465 26.145 175.480 ;
        RECT 54.335 175.465 54.665 175.480 ;
        RECT 61.940 175.480 96.525 175.780 ;
        RECT 39.615 175.100 39.945 175.115 ;
        RECT 49.735 175.100 50.065 175.115 ;
        RECT 53.875 175.100 54.205 175.115 ;
        RECT 61.940 175.100 62.240 175.480 ;
        RECT 96.195 175.465 96.525 175.480 ;
        RECT 100.335 175.780 100.665 175.795 ;
        RECT 137.595 175.780 137.925 175.795 ;
        RECT 100.335 175.480 137.925 175.780 ;
        RECT 100.335 175.465 100.665 175.480 ;
        RECT 137.595 175.465 137.925 175.480 ;
        RECT 39.615 174.800 48.440 175.100 ;
        RECT 39.615 174.785 39.945 174.800 ;
        RECT 48.140 174.430 48.440 174.800 ;
        RECT 49.735 174.800 62.240 175.100 ;
        RECT 102.175 175.100 102.505 175.115 ;
        RECT 113.675 175.100 114.005 175.115 ;
        RECT 122.415 175.100 122.745 175.115 ;
        RECT 102.175 174.800 122.745 175.100 ;
        RECT 49.735 174.785 50.065 174.800 ;
        RECT 53.875 174.785 54.205 174.800 ;
        RECT 102.175 174.785 102.505 174.800 ;
        RECT 113.675 174.785 114.005 174.800 ;
        RECT 122.415 174.785 122.745 174.800 ;
        RECT 48.100 174.110 48.480 174.430 ;
        RECT 55.715 174.420 56.045 174.435 ;
        RECT 65.375 174.420 65.705 174.435 ;
        RECT 55.715 174.120 65.705 174.420 ;
        RECT 55.715 174.105 56.045 174.120 ;
        RECT 65.375 174.105 65.705 174.120 ;
        RECT 82.395 174.420 82.725 174.435 ;
        RECT 86.535 174.420 86.865 174.435 ;
        RECT 82.395 174.120 117.440 174.420 ;
        RECT 82.395 174.105 82.725 174.120 ;
        RECT 86.535 174.105 86.865 174.120 ;
        RECT 40.830 173.765 42.410 174.095 ;
        RECT 79.700 173.765 81.280 174.095 ;
        RECT 75.955 173.740 76.285 173.755 ;
        RECT 78.715 173.740 79.045 173.755 ;
        RECT 75.955 173.440 79.045 173.740 ;
        RECT 75.955 173.425 76.285 173.440 ;
        RECT 78.715 173.425 79.045 173.440 ;
        RECT 26.735 173.060 27.065 173.075 ;
        RECT 53.415 173.060 53.745 173.075 ;
        RECT 26.735 172.760 53.745 173.060 ;
        RECT 26.735 172.745 27.065 172.760 ;
        RECT 53.415 172.745 53.745 172.760 ;
        RECT 72.275 173.060 72.605 173.075 ;
        RECT 100.795 173.060 101.125 173.075 ;
        RECT 104.015 173.060 104.345 173.075 ;
        RECT 108.615 173.060 108.945 173.075 ;
        RECT 72.275 172.760 108.945 173.060 ;
        RECT 72.275 172.745 72.605 172.760 ;
        RECT 100.795 172.745 101.125 172.760 ;
        RECT 104.015 172.745 104.345 172.760 ;
        RECT 108.615 172.745 108.945 172.760 ;
        RECT 45.595 172.380 45.925 172.395 ;
        RECT 68.135 172.380 68.465 172.395 ;
        RECT 45.595 172.080 68.465 172.380 ;
        RECT 45.595 172.065 45.925 172.080 ;
        RECT 68.135 172.065 68.465 172.080 ;
        RECT 78.715 172.380 79.045 172.395 ;
        RECT 89.755 172.380 90.085 172.395 ;
        RECT 113.215 172.380 113.545 172.395 ;
        RECT 78.715 172.080 90.085 172.380 ;
        RECT 78.715 172.065 79.045 172.080 ;
        RECT 89.755 172.065 90.085 172.080 ;
        RECT 96.440 172.080 113.545 172.380 ;
        RECT 117.140 172.380 117.440 174.120 ;
        RECT 118.570 173.765 120.150 174.095 ;
        RECT 157.440 173.765 159.020 174.095 ;
        RECT 123.795 173.740 124.125 173.755 ;
        RECT 128.395 173.740 128.725 173.755 ;
        RECT 123.795 173.440 128.725 173.740 ;
        RECT 123.795 173.425 124.125 173.440 ;
        RECT 128.395 173.425 128.725 173.440 ;
        RECT 118.735 173.060 119.065 173.075 ;
        RECT 131.615 173.060 131.945 173.075 ;
        RECT 118.735 172.760 131.945 173.060 ;
        RECT 118.735 172.745 119.065 172.760 ;
        RECT 131.615 172.745 131.945 172.760 ;
        RECT 148.635 172.380 148.965 172.395 ;
        RECT 117.140 172.080 148.965 172.380 ;
        RECT 49.735 171.700 50.065 171.715 ;
        RECT 55.255 171.700 55.585 171.715 ;
        RECT 49.735 171.400 55.585 171.700 ;
        RECT 49.735 171.385 50.065 171.400 ;
        RECT 55.255 171.385 55.585 171.400 ;
        RECT 75.035 171.700 75.365 171.715 ;
        RECT 83.315 171.700 83.645 171.715 ;
        RECT 75.035 171.400 83.645 171.700 ;
        RECT 75.035 171.385 75.365 171.400 ;
        RECT 83.315 171.385 83.645 171.400 ;
        RECT 21.395 171.045 22.975 171.375 ;
        RECT 60.265 171.045 61.845 171.375 ;
        RECT 75.035 171.020 75.365 171.035 ;
        RECT 94.355 171.020 94.685 171.035 ;
        RECT 96.440 171.020 96.740 172.080 ;
        RECT 113.215 172.065 113.545 172.080 ;
        RECT 148.635 172.065 148.965 172.080 ;
        RECT 108.615 171.700 108.945 171.715 ;
        RECT 118.735 171.700 119.065 171.715 ;
        RECT 108.615 171.400 119.065 171.700 ;
        RECT 108.615 171.385 108.945 171.400 ;
        RECT 118.735 171.385 119.065 171.400 ;
        RECT 99.135 171.045 100.715 171.375 ;
        RECT 138.005 171.045 139.585 171.375 ;
        RECT 75.035 170.720 96.740 171.020 ;
        RECT 101.715 171.020 102.045 171.035 ;
        RECT 132.995 171.020 133.325 171.035 ;
        RECT 101.715 170.720 133.325 171.020 ;
        RECT 75.035 170.705 75.365 170.720 ;
        RECT 94.355 170.705 94.685 170.720 ;
        RECT 101.715 170.705 102.045 170.720 ;
        RECT 132.995 170.705 133.325 170.720 ;
        RECT 50.195 170.340 50.525 170.355 ;
        RECT 60.315 170.340 60.645 170.355 ;
        RECT 50.195 170.040 60.645 170.340 ;
        RECT 50.195 170.025 50.525 170.040 ;
        RECT 60.315 170.025 60.645 170.040 ;
        RECT 64.915 170.340 65.245 170.355 ;
        RECT 85.615 170.340 85.945 170.355 ;
        RECT 64.915 170.040 85.945 170.340 ;
        RECT 64.915 170.025 65.245 170.040 ;
        RECT 85.615 170.025 85.945 170.040 ;
        RECT 87.915 170.340 88.245 170.355 ;
        RECT 124.255 170.340 124.585 170.355 ;
        RECT 87.915 170.040 124.585 170.340 ;
        RECT 87.915 170.025 88.245 170.040 ;
        RECT 124.255 170.025 124.585 170.040 ;
        RECT 149.555 170.340 149.885 170.355 ;
        RECT 150.220 170.340 150.600 170.350 ;
        RECT 149.555 170.040 150.600 170.340 ;
        RECT 149.555 170.025 149.885 170.040 ;
        RECT 150.220 170.030 150.600 170.040 ;
        RECT 35.475 169.660 35.805 169.675 ;
        RECT 45.135 169.660 45.465 169.675 ;
        RECT 58.475 169.660 58.805 169.675 ;
        RECT 94.815 169.660 95.145 169.675 ;
        RECT 35.475 169.360 43.150 169.660 ;
        RECT 35.475 169.345 35.805 169.360 ;
        RECT 40.830 168.325 42.410 168.655 ;
        RECT 42.850 168.300 43.150 169.360 ;
        RECT 45.135 169.360 48.440 169.660 ;
        RECT 45.135 169.345 45.465 169.360 ;
        RECT 48.140 168.980 48.440 169.360 ;
        RECT 58.475 169.360 95.145 169.660 ;
        RECT 58.475 169.345 58.805 169.360 ;
        RECT 94.815 169.345 95.145 169.360 ;
        RECT 98.955 169.660 99.285 169.675 ;
        RECT 114.135 169.660 114.465 169.675 ;
        RECT 98.955 169.360 114.465 169.660 ;
        RECT 98.955 169.345 99.285 169.360 ;
        RECT 114.135 169.345 114.465 169.360 ;
        RECT 62.155 168.980 62.485 168.995 ;
        RECT 48.140 168.680 62.485 168.980 ;
        RECT 62.155 168.665 62.485 168.680 ;
        RECT 68.595 168.980 68.925 168.995 ;
        RECT 78.715 168.980 79.045 168.995 ;
        RECT 106.775 168.980 107.105 168.995 ;
        RECT 68.595 168.680 79.045 168.980 ;
        RECT 68.595 168.665 68.925 168.680 ;
        RECT 78.715 168.665 79.045 168.680 ;
        RECT 102.190 168.680 107.105 168.980 ;
        RECT 79.700 168.325 81.280 168.655 ;
        RECT 102.190 168.315 102.490 168.680 ;
        RECT 106.775 168.665 107.105 168.680 ;
        RECT 118.570 168.325 120.150 168.655 ;
        RECT 157.440 168.325 159.020 168.655 ;
        RECT 63.535 168.300 63.865 168.315 ;
        RECT 68.595 168.300 68.925 168.315 ;
        RECT 42.850 168.000 68.925 168.300 ;
        RECT 63.535 167.985 63.865 168.000 ;
        RECT 68.595 167.985 68.925 168.000 ;
        RECT 81.935 168.300 82.265 168.315 ;
        RECT 102.175 168.300 102.505 168.315 ;
        RECT 81.935 168.000 102.505 168.300 ;
        RECT 81.935 167.985 82.265 168.000 ;
        RECT 102.175 167.985 102.505 168.000 ;
        RECT 57.555 167.620 57.885 167.635 ;
        RECT 77.335 167.620 77.665 167.635 ;
        RECT 57.555 167.320 77.665 167.620 ;
        RECT 57.555 167.305 57.885 167.320 ;
        RECT 77.335 167.305 77.665 167.320 ;
        RECT 78.255 167.620 78.585 167.635 ;
        RECT 109.535 167.620 109.865 167.635 ;
        RECT 78.255 167.320 109.865 167.620 ;
        RECT 78.255 167.305 78.585 167.320 ;
        RECT 109.535 167.305 109.865 167.320 ;
        RECT 26.275 166.940 26.605 166.955 ;
        RECT 48.355 166.940 48.685 166.955 ;
        RECT 26.275 166.640 48.685 166.940 ;
        RECT 26.275 166.625 26.605 166.640 ;
        RECT 48.355 166.625 48.685 166.640 ;
        RECT 56.635 166.940 56.965 166.955 ;
        RECT 74.575 166.940 74.905 166.955 ;
        RECT 56.635 166.640 74.905 166.940 ;
        RECT 56.635 166.625 56.965 166.640 ;
        RECT 74.575 166.625 74.905 166.640 ;
        RECT 83.315 166.940 83.645 166.955 ;
        RECT 91.595 166.940 91.925 166.955 ;
        RECT 83.315 166.640 91.925 166.940 ;
        RECT 83.315 166.625 83.645 166.640 ;
        RECT 91.595 166.625 91.925 166.640 ;
        RECT 98.495 166.940 98.825 166.955 ;
        RECT 122.875 166.940 123.205 166.955 ;
        RECT 98.495 166.640 123.205 166.940 ;
        RECT 98.495 166.625 98.825 166.640 ;
        RECT 122.875 166.625 123.205 166.640 ;
        RECT 44.675 166.270 45.005 166.275 ;
        RECT 44.420 166.260 45.005 166.270 ;
        RECT 51.575 166.260 51.905 166.275 ;
        RECT 44.420 165.960 51.905 166.260 ;
        RECT 44.420 165.950 45.005 165.960 ;
        RECT 44.675 165.945 45.005 165.950 ;
        RECT 51.575 165.945 51.905 165.960 ;
        RECT 52.495 166.260 52.825 166.275 ;
        RECT 58.935 166.260 59.265 166.275 ;
        RECT 52.495 165.960 59.265 166.260 ;
        RECT 52.495 165.945 52.825 165.960 ;
        RECT 58.935 165.945 59.265 165.960 ;
        RECT 67.215 166.260 67.545 166.275 ;
        RECT 92.515 166.260 92.845 166.275 ;
        RECT 67.215 165.960 92.845 166.260 ;
        RECT 67.215 165.945 67.545 165.960 ;
        RECT 92.515 165.945 92.845 165.960 ;
        RECT 21.395 165.605 22.975 165.935 ;
        RECT 60.265 165.605 61.845 165.935 ;
        RECT 99.135 165.605 100.715 165.935 ;
        RECT 138.005 165.605 139.585 165.935 ;
        RECT 53.620 165.580 54.000 165.590 ;
        RECT 54.335 165.580 54.665 165.595 ;
        RECT 53.620 165.280 54.665 165.580 ;
        RECT 53.620 165.270 54.000 165.280 ;
        RECT 54.335 165.265 54.665 165.280 ;
        RECT 76.875 165.265 77.205 165.595 ;
        RECT 20.295 164.900 20.625 164.915 ;
        RECT 38.695 164.900 39.025 164.915 ;
        RECT 20.295 164.600 39.025 164.900 ;
        RECT 20.295 164.585 20.625 164.600 ;
        RECT 38.695 164.585 39.025 164.600 ;
        RECT 43.295 164.900 43.625 164.915 ;
        RECT 56.635 164.900 56.965 164.915 ;
        RECT 66.755 164.900 67.085 164.915 ;
        RECT 43.295 164.600 67.085 164.900 ;
        RECT 43.295 164.585 43.625 164.600 ;
        RECT 56.635 164.585 56.965 164.600 ;
        RECT 66.755 164.585 67.085 164.600 ;
        RECT 32.715 164.220 33.045 164.235 ;
        RECT 76.890 164.220 77.190 165.265 ;
        RECT 80.555 164.900 80.885 164.915 ;
        RECT 124.715 164.900 125.045 164.915 ;
        RECT 80.555 164.600 125.045 164.900 ;
        RECT 80.555 164.585 80.885 164.600 ;
        RECT 124.715 164.585 125.045 164.600 ;
        RECT 102.175 164.220 102.505 164.235 ;
        RECT 132.535 164.220 132.865 164.235 ;
        RECT 32.715 163.920 77.190 164.220 ;
        RECT 78.500 163.920 102.505 164.220 ;
        RECT 32.715 163.905 33.045 163.920 ;
        RECT 50.655 163.540 50.985 163.555 ;
        RECT 52.495 163.540 52.825 163.555 ;
        RECT 50.655 163.240 52.825 163.540 ;
        RECT 50.655 163.225 50.985 163.240 ;
        RECT 52.495 163.225 52.825 163.240 ;
        RECT 54.795 163.540 55.125 163.555 ;
        RECT 65.835 163.540 66.165 163.555 ;
        RECT 54.795 163.240 66.165 163.540 ;
        RECT 54.795 163.225 55.125 163.240 ;
        RECT 65.835 163.225 66.165 163.240 ;
        RECT 68.135 163.540 68.465 163.555 ;
        RECT 78.500 163.540 78.800 163.920 ;
        RECT 102.175 163.905 102.505 163.920 ;
        RECT 110.240 163.920 132.865 164.220 ;
        RECT 68.135 163.240 78.800 163.540 ;
        RECT 94.815 163.540 95.145 163.555 ;
        RECT 96.655 163.540 96.985 163.555 ;
        RECT 110.240 163.540 110.540 163.920 ;
        RECT 132.535 163.905 132.865 163.920 ;
        RECT 94.815 163.240 110.540 163.540 ;
        RECT 68.135 163.225 68.465 163.240 ;
        RECT 94.815 163.225 95.145 163.240 ;
        RECT 96.655 163.225 96.985 163.240 ;
        RECT 40.830 162.885 42.410 163.215 ;
        RECT 79.700 162.885 81.280 163.215 ;
        RECT 118.570 162.885 120.150 163.215 ;
        RECT 157.440 162.885 159.020 163.215 ;
        RECT 60.775 162.860 61.105 162.875 ;
        RECT 74.575 162.860 74.905 162.875 ;
        RECT 60.775 162.560 74.905 162.860 ;
        RECT 60.775 162.545 61.105 162.560 ;
        RECT 74.575 162.545 74.905 162.560 ;
        RECT 40.995 162.180 41.325 162.195 ;
        RECT 67.675 162.180 68.005 162.195 ;
        RECT 40.995 161.880 68.005 162.180 ;
        RECT 40.995 161.865 41.325 161.880 ;
        RECT 67.675 161.865 68.005 161.880 ;
        RECT 94.355 162.180 94.685 162.195 ;
        RECT 138.055 162.180 138.385 162.195 ;
        RECT 94.355 161.880 138.385 162.180 ;
        RECT 94.355 161.865 94.685 161.880 ;
        RECT 138.055 161.865 138.385 161.880 ;
        RECT 34.555 161.500 34.885 161.515 ;
        RECT 35.220 161.500 35.600 161.510 ;
        RECT 34.555 161.200 35.600 161.500 ;
        RECT 34.555 161.185 34.885 161.200 ;
        RECT 35.220 161.190 35.600 161.200 ;
        RECT 41.455 161.500 41.785 161.515 ;
        RECT 60.775 161.500 61.105 161.515 ;
        RECT 41.455 161.200 61.105 161.500 ;
        RECT 41.455 161.185 41.785 161.200 ;
        RECT 60.775 161.185 61.105 161.200 ;
        RECT 61.695 161.500 62.025 161.515 ;
        RECT 73.655 161.500 73.985 161.515 ;
        RECT 104.475 161.500 104.805 161.515 ;
        RECT 61.695 161.200 73.985 161.500 ;
        RECT 61.695 161.185 62.025 161.200 ;
        RECT 73.655 161.185 73.985 161.200 ;
        RECT 97.820 161.200 104.805 161.500 ;
        RECT 54.335 160.820 54.665 160.835 ;
        RECT 59.395 160.820 59.725 160.835 ;
        RECT 54.335 160.520 59.725 160.820 ;
        RECT 54.335 160.505 54.665 160.520 ;
        RECT 59.395 160.505 59.725 160.520 ;
        RECT 63.995 160.820 64.325 160.835 ;
        RECT 97.820 160.820 98.120 161.200 ;
        RECT 104.475 161.185 104.805 161.200 ;
        RECT 118.275 161.500 118.605 161.515 ;
        RECT 121.035 161.500 121.365 161.515 ;
        RECT 135.500 161.500 135.880 161.510 ;
        RECT 118.275 161.200 135.880 161.500 ;
        RECT 118.275 161.185 118.605 161.200 ;
        RECT 121.035 161.185 121.365 161.200 ;
        RECT 135.500 161.190 135.880 161.200 ;
        RECT 63.995 160.520 98.120 160.820 ;
        RECT 105.855 160.820 106.185 160.835 ;
        RECT 121.955 160.820 122.285 160.835 ;
        RECT 127.935 160.820 128.265 160.835 ;
        RECT 130.235 160.820 130.565 160.835 ;
        RECT 105.855 160.520 130.565 160.820 ;
        RECT 63.995 160.505 64.325 160.520 ;
        RECT 105.855 160.505 106.185 160.520 ;
        RECT 121.955 160.505 122.285 160.520 ;
        RECT 127.935 160.505 128.265 160.520 ;
        RECT 130.235 160.505 130.565 160.520 ;
        RECT 21.395 160.165 22.975 160.495 ;
        RECT 60.265 160.165 61.845 160.495 ;
        RECT 99.135 160.165 100.715 160.495 ;
        RECT 138.005 160.165 139.585 160.495 ;
        RECT 101.500 159.840 104.560 160.140 ;
        RECT 25.815 159.460 26.145 159.475 ;
        RECT 30.875 159.460 31.205 159.475 ;
        RECT 36.855 159.460 37.185 159.475 ;
        RECT 61.235 159.460 61.565 159.475 ;
        RECT 25.815 159.160 37.185 159.460 ;
        RECT 25.815 159.145 26.145 159.160 ;
        RECT 30.875 159.145 31.205 159.160 ;
        RECT 36.855 159.145 37.185 159.160 ;
        RECT 48.140 159.160 61.565 159.460 ;
        RECT 30.415 158.780 30.745 158.795 ;
        RECT 44.215 158.780 44.545 158.795 ;
        RECT 48.140 158.780 48.440 159.160 ;
        RECT 61.235 159.145 61.565 159.160 ;
        RECT 72.735 159.460 73.065 159.475 ;
        RECT 79.175 159.460 79.505 159.475 ;
        RECT 101.500 159.460 101.800 159.840 ;
        RECT 72.735 159.160 101.800 159.460 ;
        RECT 102.380 159.460 102.760 159.470 ;
        RECT 103.095 159.460 103.425 159.475 ;
        RECT 102.380 159.160 103.425 159.460 ;
        RECT 104.260 159.460 104.560 159.840 ;
        RECT 106.775 159.460 107.105 159.475 ;
        RECT 104.260 159.160 107.105 159.460 ;
        RECT 72.735 159.145 73.065 159.160 ;
        RECT 79.175 159.145 79.505 159.160 ;
        RECT 102.380 159.150 102.760 159.160 ;
        RECT 103.095 159.145 103.425 159.160 ;
        RECT 106.775 159.145 107.105 159.160 ;
        RECT 114.135 159.460 114.465 159.475 ;
        RECT 115.515 159.460 115.845 159.475 ;
        RECT 138.975 159.460 139.305 159.475 ;
        RECT 114.135 159.160 139.305 159.460 ;
        RECT 114.135 159.145 114.465 159.160 ;
        RECT 115.515 159.145 115.845 159.160 ;
        RECT 138.975 159.145 139.305 159.160 ;
        RECT 30.415 158.480 48.440 158.780 ;
        RECT 59.140 158.780 59.520 158.790 ;
        RECT 131.155 158.780 131.485 158.795 ;
        RECT 59.140 158.480 131.485 158.780 ;
        RECT 30.415 158.465 30.745 158.480 ;
        RECT 44.215 158.465 44.545 158.480 ;
        RECT 59.140 158.470 59.520 158.480 ;
        RECT 131.155 158.465 131.485 158.480 ;
        RECT 48.100 158.100 48.480 158.110 ;
        RECT 50.655 158.100 50.985 158.115 ;
        RECT 48.100 157.800 50.985 158.100 ;
        RECT 48.100 157.790 48.480 157.800 ;
        RECT 50.655 157.785 50.985 157.800 ;
        RECT 55.255 158.100 55.585 158.115 ;
        RECT 70.895 158.100 71.225 158.115 ;
        RECT 55.255 157.800 71.225 158.100 ;
        RECT 55.255 157.785 55.585 157.800 ;
        RECT 70.895 157.785 71.225 157.800 ;
        RECT 40.830 157.445 42.410 157.775 ;
        RECT 79.700 157.445 81.280 157.775 ;
        RECT 118.570 157.445 120.150 157.775 ;
        RECT 157.440 157.445 159.020 157.775 ;
        RECT 23.515 157.420 23.845 157.435 ;
        RECT 35.935 157.420 36.265 157.435 ;
        RECT 40.075 157.420 40.405 157.435 ;
        RECT 23.515 157.120 40.405 157.420 ;
        RECT 23.515 157.105 23.845 157.120 ;
        RECT 35.935 157.105 36.265 157.120 ;
        RECT 40.075 157.105 40.405 157.120 ;
        RECT 53.415 157.430 53.745 157.435 ;
        RECT 53.415 157.420 54.000 157.430 ;
        RECT 63.535 157.420 63.865 157.435 ;
        RECT 76.875 157.420 77.205 157.435 ;
        RECT 53.415 157.120 54.200 157.420 ;
        RECT 63.535 157.120 77.205 157.420 ;
        RECT 53.415 157.110 54.000 157.120 ;
        RECT 53.415 157.105 53.745 157.110 ;
        RECT 63.535 157.105 63.865 157.120 ;
        RECT 76.875 157.105 77.205 157.120 ;
        RECT 28.575 156.740 28.905 156.755 ;
        RECT 95.735 156.740 96.065 156.755 ;
        RECT 28.575 156.440 96.065 156.740 ;
        RECT 28.575 156.425 28.905 156.440 ;
        RECT 95.735 156.425 96.065 156.440 ;
        RECT 102.635 156.740 102.965 156.755 ;
        RECT 124.255 156.740 124.585 156.755 ;
        RECT 102.635 156.440 124.585 156.740 ;
        RECT 102.635 156.425 102.965 156.440 ;
        RECT 124.255 156.425 124.585 156.440 ;
        RECT 16.155 156.060 16.485 156.075 ;
        RECT 25.815 156.060 26.145 156.075 ;
        RECT 16.155 155.760 26.145 156.060 ;
        RECT 16.155 155.745 16.485 155.760 ;
        RECT 25.815 155.745 26.145 155.760 ;
        RECT 35.475 156.060 35.805 156.075 ;
        RECT 40.535 156.060 40.865 156.075 ;
        RECT 35.475 155.760 40.865 156.060 ;
        RECT 35.475 155.745 35.805 155.760 ;
        RECT 40.535 155.745 40.865 155.760 ;
        RECT 42.375 156.060 42.705 156.075 ;
        RECT 49.735 156.070 50.065 156.075 ;
        RECT 49.020 156.060 49.400 156.070 ;
        RECT 42.375 155.760 49.400 156.060 ;
        RECT 42.375 155.745 42.705 155.760 ;
        RECT 49.020 155.750 49.400 155.760 ;
        RECT 49.735 156.060 50.320 156.070 ;
        RECT 52.035 156.060 52.365 156.075 ;
        RECT 60.315 156.060 60.645 156.075 ;
        RECT 49.735 155.760 50.520 156.060 ;
        RECT 52.035 155.760 60.645 156.060 ;
        RECT 49.735 155.750 50.320 155.760 ;
        RECT 49.735 155.745 50.065 155.750 ;
        RECT 52.035 155.745 52.365 155.760 ;
        RECT 60.315 155.745 60.645 155.760 ;
        RECT 84.695 156.060 85.025 156.075 ;
        RECT 121.035 156.060 121.365 156.075 ;
        RECT 84.695 155.760 121.365 156.060 ;
        RECT 84.695 155.745 85.025 155.760 ;
        RECT 121.035 155.745 121.365 155.760 ;
        RECT 30.415 155.380 30.745 155.395 ;
        RECT 39.615 155.380 39.945 155.395 ;
        RECT 47.435 155.390 47.765 155.395 ;
        RECT 47.180 155.380 47.765 155.390 ;
        RECT 53.415 155.380 53.745 155.395 ;
        RECT 30.415 155.080 39.945 155.380 ;
        RECT 46.800 155.080 53.745 155.380 ;
        RECT 30.415 155.065 30.745 155.080 ;
        RECT 39.615 155.065 39.945 155.080 ;
        RECT 47.180 155.070 47.765 155.080 ;
        RECT 47.435 155.065 47.765 155.070 ;
        RECT 53.415 155.065 53.745 155.080 ;
        RECT 55.255 155.380 55.585 155.395 ;
        RECT 57.095 155.380 57.425 155.395 ;
        RECT 55.255 155.080 57.425 155.380 ;
        RECT 55.255 155.065 55.585 155.080 ;
        RECT 57.095 155.065 57.425 155.080 ;
        RECT 21.395 154.725 22.975 155.055 ;
        RECT 60.265 154.725 61.845 155.055 ;
        RECT 99.135 154.725 100.715 155.055 ;
        RECT 138.005 154.725 139.585 155.055 ;
        RECT 39.615 154.700 39.945 154.715 ;
        RECT 55.255 154.700 55.585 154.715 ;
        RECT 81.935 154.700 82.265 154.715 ;
        RECT 39.615 154.400 55.585 154.700 ;
        RECT 39.615 154.385 39.945 154.400 ;
        RECT 55.255 154.385 55.585 154.400 ;
        RECT 62.170 154.400 82.265 154.700 ;
        RECT 33.635 154.020 33.965 154.035 ;
        RECT 41.915 154.020 42.245 154.035 ;
        RECT 44.215 154.020 44.545 154.035 ;
        RECT 33.635 153.720 44.545 154.020 ;
        RECT 33.635 153.705 33.965 153.720 ;
        RECT 41.915 153.705 42.245 153.720 ;
        RECT 44.215 153.705 44.545 153.720 ;
        RECT 53.415 154.020 53.745 154.035 ;
        RECT 62.170 154.020 62.470 154.400 ;
        RECT 81.935 154.385 82.265 154.400 ;
        RECT 53.415 153.720 62.470 154.020 ;
        RECT 63.740 154.020 64.120 154.030 ;
        RECT 95.735 154.020 96.065 154.035 ;
        RECT 63.740 153.720 96.065 154.020 ;
        RECT 53.415 153.705 53.745 153.720 ;
        RECT 63.740 153.710 64.120 153.720 ;
        RECT 95.735 153.705 96.065 153.720 ;
        RECT 98.955 154.020 99.285 154.035 ;
        RECT 115.975 154.020 116.305 154.035 ;
        RECT 98.955 153.720 116.305 154.020 ;
        RECT 98.955 153.705 99.285 153.720 ;
        RECT 115.975 153.705 116.305 153.720 ;
        RECT 28.115 153.340 28.445 153.355 ;
        RECT 36.395 153.340 36.725 153.355 ;
        RECT 37.060 153.340 37.440 153.350 ;
        RECT 28.115 153.040 37.440 153.340 ;
        RECT 28.115 153.025 28.445 153.040 ;
        RECT 36.395 153.025 36.725 153.040 ;
        RECT 37.060 153.030 37.440 153.040 ;
        RECT 41.915 153.340 42.245 153.355 ;
        RECT 56.175 153.340 56.505 153.355 ;
        RECT 41.915 153.040 56.505 153.340 ;
        RECT 41.915 153.025 42.245 153.040 ;
        RECT 56.175 153.025 56.505 153.040 ;
        RECT 50.860 152.660 51.240 152.670 ;
        RECT 57.555 152.660 57.885 152.675 ;
        RECT 44.460 152.360 57.885 152.660 ;
        RECT 40.830 152.005 42.410 152.335 ;
        RECT 10.175 151.980 10.505 151.995 ;
        RECT 14.315 151.980 14.645 151.995 ;
        RECT 10.175 151.680 14.645 151.980 ;
        RECT 10.175 151.665 10.505 151.680 ;
        RECT 14.315 151.665 14.645 151.680 ;
        RECT 20.295 151.980 20.625 151.995 ;
        RECT 32.255 151.980 32.585 151.995 ;
        RECT 20.295 151.680 32.585 151.980 ;
        RECT 20.295 151.665 20.625 151.680 ;
        RECT 32.255 151.665 32.585 151.680 ;
        RECT 44.460 151.315 44.760 152.360 ;
        RECT 50.860 152.350 51.240 152.360 ;
        RECT 57.555 152.345 57.885 152.360 ;
        RECT 63.740 152.350 64.120 152.670 ;
        RECT 45.135 151.980 45.465 151.995 ;
        RECT 47.895 151.980 48.225 151.995 ;
        RECT 45.135 151.680 48.225 151.980 ;
        RECT 45.135 151.665 45.465 151.680 ;
        RECT 47.895 151.665 48.225 151.680 ;
        RECT 49.275 151.980 49.605 151.995 ;
        RECT 49.940 151.980 50.320 151.990 ;
        RECT 49.275 151.680 50.320 151.980 ;
        RECT 49.275 151.665 49.605 151.680 ;
        RECT 49.940 151.670 50.320 151.680 ;
        RECT 51.115 151.980 51.445 151.995 ;
        RECT 63.780 151.980 64.080 152.350 ;
        RECT 79.700 152.005 81.280 152.335 ;
        RECT 118.570 152.005 120.150 152.335 ;
        RECT 157.440 152.005 159.020 152.335 ;
        RECT 51.115 151.680 64.080 151.980 ;
        RECT 102.635 151.980 102.965 151.995 ;
        RECT 113.675 151.980 114.005 151.995 ;
        RECT 102.635 151.680 114.005 151.980 ;
        RECT 51.115 151.665 51.445 151.680 ;
        RECT 102.635 151.665 102.965 151.680 ;
        RECT 113.675 151.665 114.005 151.680 ;
        RECT 29.495 151.300 29.825 151.315 ;
        RECT 35.015 151.300 35.345 151.315 ;
        RECT 42.835 151.300 43.165 151.315 ;
        RECT 29.495 151.000 35.345 151.300 ;
        RECT 29.495 150.985 29.825 151.000 ;
        RECT 35.015 150.985 35.345 151.000 ;
        RECT 41.240 151.000 43.165 151.300 ;
        RECT 44.460 151.000 45.005 151.315 ;
        RECT 41.240 150.635 41.540 151.000 ;
        RECT 42.835 150.985 43.165 151.000 ;
        RECT 44.675 150.985 45.005 151.000 ;
        RECT 48.815 151.300 49.145 151.315 ;
        RECT 96.655 151.300 96.985 151.315 ;
        RECT 48.815 151.000 96.985 151.300 ;
        RECT 48.815 150.985 49.145 151.000 ;
        RECT 96.655 150.985 96.985 151.000 ;
        RECT 111.835 151.300 112.165 151.315 ;
        RECT 129.775 151.300 130.105 151.315 ;
        RECT 111.835 151.000 130.105 151.300 ;
        RECT 111.835 150.985 112.165 151.000 ;
        RECT 129.775 150.985 130.105 151.000 ;
        RECT 27.195 150.620 27.525 150.635 ;
        RECT 40.075 150.630 40.405 150.635 ;
        RECT 34.300 150.620 34.680 150.630 ;
        RECT 39.820 150.620 40.405 150.630 ;
        RECT 27.195 150.320 34.680 150.620 ;
        RECT 39.620 150.320 40.405 150.620 ;
        RECT 27.195 150.305 27.525 150.320 ;
        RECT 34.300 150.310 34.680 150.320 ;
        RECT 39.820 150.310 40.405 150.320 ;
        RECT 40.075 150.305 40.405 150.310 ;
        RECT 40.995 150.320 41.540 150.635 ;
        RECT 43.295 150.630 43.625 150.635 ;
        RECT 43.295 150.620 43.880 150.630 ;
        RECT 101.255 150.620 101.585 150.635 ;
        RECT 43.070 150.320 43.880 150.620 ;
        RECT 40.995 150.305 41.325 150.320 ;
        RECT 43.295 150.310 43.880 150.320 ;
        RECT 44.460 150.320 101.585 150.620 ;
        RECT 43.295 150.305 43.625 150.310 ;
        RECT 27.195 149.950 27.525 149.955 ;
        RECT 26.940 149.940 27.525 149.950 ;
        RECT 44.460 149.940 44.760 150.320 ;
        RECT 101.255 150.305 101.585 150.320 ;
        RECT 108.615 150.620 108.945 150.635 ;
        RECT 129.315 150.620 129.645 150.635 ;
        RECT 141.735 150.620 142.065 150.635 ;
        RECT 108.615 150.320 142.065 150.620 ;
        RECT 108.615 150.305 108.945 150.320 ;
        RECT 129.315 150.305 129.645 150.320 ;
        RECT 141.735 150.305 142.065 150.320 ;
        RECT 48.815 149.940 49.145 149.955 ;
        RECT 53.875 149.950 54.205 149.955 ;
        RECT 53.620 149.940 54.205 149.950 ;
        RECT 26.560 149.640 44.760 149.940 ;
        RECT 45.380 149.640 49.145 149.940 ;
        RECT 53.420 149.640 54.205 149.940 ;
        RECT 26.940 149.630 27.525 149.640 ;
        RECT 27.195 149.625 27.525 149.630 ;
        RECT 21.395 149.285 22.975 149.615 ;
        RECT 31.540 149.260 31.920 149.270 ;
        RECT 45.380 149.260 45.680 149.640 ;
        RECT 48.815 149.625 49.145 149.640 ;
        RECT 53.620 149.630 54.205 149.640 ;
        RECT 53.875 149.625 54.205 149.630 ;
        RECT 54.795 149.940 55.125 149.955 ;
        RECT 59.140 149.940 59.520 149.950 ;
        RECT 54.795 149.640 59.520 149.940 ;
        RECT 54.795 149.625 55.125 149.640 ;
        RECT 59.140 149.630 59.520 149.640 ;
        RECT 103.555 149.940 103.885 149.955 ;
        RECT 116.895 149.940 117.225 149.955 ;
        RECT 103.555 149.640 117.225 149.940 ;
        RECT 103.555 149.625 103.885 149.640 ;
        RECT 116.895 149.625 117.225 149.640 ;
        RECT 60.265 149.285 61.845 149.615 ;
        RECT 99.135 149.285 100.715 149.615 ;
        RECT 138.005 149.285 139.585 149.615 ;
        RECT 31.540 148.960 45.680 149.260 ;
        RECT 49.735 149.260 50.065 149.275 ;
        RECT 52.700 149.260 53.080 149.270 ;
        RECT 49.735 148.960 59.480 149.260 ;
        RECT 31.540 148.950 31.920 148.960 ;
        RECT 49.735 148.945 50.065 148.960 ;
        RECT 52.700 148.950 53.080 148.960 ;
        RECT 5.115 148.580 5.445 148.595 ;
        RECT 53.415 148.580 53.745 148.595 ;
        RECT 5.115 148.280 53.745 148.580 ;
        RECT 59.180 148.580 59.480 148.960 ;
        RECT 91.135 148.945 91.465 149.275 ;
        RECT 91.150 148.580 91.450 148.945 ;
        RECT 59.180 148.280 91.450 148.580 ;
        RECT 5.115 148.265 5.445 148.280 ;
        RECT 53.415 148.265 53.745 148.280 ;
        RECT 33.635 147.900 33.965 147.915 ;
        RECT 51.115 147.900 51.445 147.915 ;
        RECT 58.015 147.900 58.345 147.915 ;
        RECT 126.095 147.900 126.425 147.915 ;
        RECT 33.635 147.600 43.840 147.900 ;
        RECT 33.635 147.585 33.965 147.600 ;
        RECT 27.195 147.220 27.525 147.235 ;
        RECT 36.395 147.220 36.725 147.235 ;
        RECT 27.195 146.920 36.725 147.220 ;
        RECT 43.540 147.220 43.840 147.600 ;
        RECT 51.115 147.600 58.345 147.900 ;
        RECT 51.115 147.585 51.445 147.600 ;
        RECT 58.015 147.585 58.345 147.600 ;
        RECT 61.940 147.600 126.425 147.900 ;
        RECT 61.940 147.220 62.240 147.600 ;
        RECT 126.095 147.585 126.425 147.600 ;
        RECT 43.540 146.920 62.240 147.220 ;
        RECT 100.795 147.220 101.125 147.235 ;
        RECT 102.175 147.220 102.505 147.235 ;
        RECT 100.795 146.920 102.505 147.220 ;
        RECT 27.195 146.905 27.525 146.920 ;
        RECT 36.395 146.905 36.725 146.920 ;
        RECT 100.795 146.905 101.125 146.920 ;
        RECT 102.175 146.905 102.505 146.920 ;
        RECT 40.830 146.565 42.410 146.895 ;
        RECT 79.700 146.565 81.280 146.895 ;
        RECT 118.570 146.565 120.150 146.895 ;
        RECT 157.440 146.565 159.020 146.895 ;
        RECT 19.375 146.540 19.705 146.555 ;
        RECT 43.755 146.540 44.085 146.555 ;
        RECT 47.180 146.540 47.560 146.550 ;
        RECT 19.375 146.240 28.200 146.540 ;
        RECT 19.375 146.225 19.705 146.240 ;
        RECT 8.795 145.860 9.125 145.875 ;
        RECT 27.195 145.860 27.525 145.875 ;
        RECT 8.795 145.560 27.525 145.860 ;
        RECT 27.900 145.860 28.200 146.240 ;
        RECT 43.755 146.240 47.560 146.540 ;
        RECT 43.755 146.225 44.085 146.240 ;
        RECT 47.180 146.230 47.560 146.240 ;
        RECT 54.540 146.540 54.920 146.550 ;
        RECT 102.635 146.540 102.965 146.555 ;
        RECT 54.540 146.240 78.800 146.540 ;
        RECT 54.540 146.230 54.920 146.240 ;
        RECT 52.035 145.860 52.365 145.875 ;
        RECT 27.900 145.560 52.365 145.860 ;
        RECT 8.795 145.545 9.125 145.560 ;
        RECT 27.195 145.545 27.525 145.560 ;
        RECT 52.035 145.545 52.365 145.560 ;
        RECT 9.715 145.180 10.045 145.195 ;
        RECT 22.595 145.180 22.925 145.195 ;
        RECT 9.715 144.880 22.925 145.180 ;
        RECT 9.715 144.865 10.045 144.880 ;
        RECT 22.595 144.865 22.925 144.880 ;
        RECT 27.195 145.180 27.525 145.195 ;
        RECT 40.995 145.180 41.325 145.195 ;
        RECT 27.195 144.880 41.325 145.180 ;
        RECT 27.195 144.865 27.525 144.880 ;
        RECT 40.995 144.865 41.325 144.880 ;
        RECT 42.375 145.180 42.705 145.195 ;
        RECT 43.500 145.180 43.880 145.190 ;
        RECT 42.375 144.880 43.880 145.180 ;
        RECT 42.375 144.865 42.705 144.880 ;
        RECT 43.500 144.870 43.880 144.880 ;
        RECT 48.815 145.180 49.145 145.195 ;
        RECT 54.580 145.180 54.880 146.230 ;
        RECT 58.935 145.860 59.265 145.875 ;
        RECT 63.995 145.860 64.325 145.875 ;
        RECT 58.935 145.560 64.325 145.860 ;
        RECT 78.500 145.860 78.800 146.240 ;
        RECT 82.180 146.240 102.965 146.540 ;
        RECT 82.180 145.860 82.480 146.240 ;
        RECT 102.635 146.225 102.965 146.240 ;
        RECT 78.500 145.560 82.480 145.860 ;
        RECT 82.855 145.860 83.185 145.875 ;
        RECT 113.215 145.860 113.545 145.875 ;
        RECT 82.855 145.560 113.545 145.860 ;
        RECT 58.935 145.545 59.265 145.560 ;
        RECT 63.995 145.545 64.325 145.560 ;
        RECT 82.855 145.545 83.185 145.560 ;
        RECT 113.215 145.545 113.545 145.560 ;
        RECT 68.135 145.180 68.465 145.195 ;
        RECT 48.815 144.880 54.880 145.180 ;
        RECT 56.420 144.880 68.465 145.180 ;
        RECT 48.815 144.865 49.145 144.880 ;
        RECT 24.895 144.500 25.225 144.515 ;
        RECT 31.540 144.500 31.920 144.510 ;
        RECT 24.895 144.200 31.920 144.500 ;
        RECT 24.895 144.185 25.225 144.200 ;
        RECT 31.540 144.190 31.920 144.200 ;
        RECT 33.175 144.500 33.505 144.515 ;
        RECT 51.575 144.500 51.905 144.515 ;
        RECT 33.175 144.200 51.905 144.500 ;
        RECT 33.175 144.185 33.505 144.200 ;
        RECT 51.575 144.185 51.905 144.200 ;
        RECT 21.395 143.845 22.975 144.175 ;
        RECT 56.420 143.835 56.720 144.880 ;
        RECT 68.135 144.865 68.465 144.880 ;
        RECT 73.655 145.180 73.985 145.195 ;
        RECT 114.135 145.180 114.465 145.195 ;
        RECT 73.655 144.880 114.465 145.180 ;
        RECT 73.655 144.865 73.985 144.880 ;
        RECT 114.135 144.865 114.465 144.880 ;
        RECT 120.575 145.180 120.905 145.195 ;
        RECT 127.935 145.180 128.265 145.195 ;
        RECT 120.575 144.880 128.265 145.180 ;
        RECT 120.575 144.865 120.905 144.880 ;
        RECT 127.935 144.865 128.265 144.880 ;
        RECT 64.915 144.500 65.245 144.515 ;
        RECT 71.355 144.500 71.685 144.515 ;
        RECT 82.855 144.500 83.185 144.515 ;
        RECT 64.915 144.200 83.185 144.500 ;
        RECT 64.915 144.185 65.245 144.200 ;
        RECT 71.355 144.185 71.685 144.200 ;
        RECT 82.855 144.185 83.185 144.200 ;
        RECT 109.075 144.500 109.405 144.515 ;
        RECT 127.015 144.500 127.345 144.515 ;
        RECT 109.075 144.200 127.345 144.500 ;
        RECT 109.075 144.185 109.405 144.200 ;
        RECT 127.015 144.185 127.345 144.200 ;
        RECT 60.265 143.845 61.845 144.175 ;
        RECT 99.135 143.845 100.715 144.175 ;
        RECT 138.005 143.845 139.585 144.175 ;
        RECT 29.035 143.820 29.365 143.835 ;
        RECT 56.175 143.820 56.720 143.835 ;
        RECT 29.035 143.520 56.720 143.820 ;
        RECT 62.155 143.820 62.485 143.835 ;
        RECT 84.695 143.820 85.025 143.835 ;
        RECT 62.155 143.520 85.025 143.820 ;
        RECT 29.035 143.505 29.365 143.520 ;
        RECT 56.175 143.505 56.505 143.520 ;
        RECT 62.155 143.505 62.485 143.520 ;
        RECT 84.695 143.505 85.025 143.520 ;
        RECT 109.995 143.820 110.325 143.835 ;
        RECT 128.395 143.820 128.725 143.835 ;
        RECT 133.455 143.820 133.785 143.835 ;
        RECT 109.995 143.520 133.785 143.820 ;
        RECT 109.995 143.505 110.325 143.520 ;
        RECT 128.395 143.505 128.725 143.520 ;
        RECT 133.455 143.505 133.785 143.520 ;
        RECT 39.155 143.140 39.485 143.155 ;
        RECT 67.675 143.140 68.005 143.155 ;
        RECT 39.155 142.840 68.005 143.140 ;
        RECT 39.155 142.825 39.485 142.840 ;
        RECT 67.675 142.825 68.005 142.840 ;
        RECT 120.115 143.140 120.445 143.155 ;
        RECT 127.475 143.140 127.805 143.155 ;
        RECT 120.115 142.840 127.805 143.140 ;
        RECT 120.115 142.825 120.445 142.840 ;
        RECT 127.475 142.825 127.805 142.840 ;
        RECT 19.835 142.460 20.165 142.475 ;
        RECT 53.415 142.460 53.745 142.475 ;
        RECT 19.835 142.160 53.745 142.460 ;
        RECT 19.835 142.145 20.165 142.160 ;
        RECT 53.415 142.145 53.745 142.160 ;
        RECT 124.715 142.460 125.045 142.475 ;
        RECT 138.055 142.460 138.385 142.475 ;
        RECT 124.715 142.160 138.385 142.460 ;
        RECT 124.715 142.145 125.045 142.160 ;
        RECT 138.055 142.145 138.385 142.160 ;
        RECT 37.060 141.780 37.440 141.790 ;
        RECT 38.695 141.780 39.025 141.795 ;
        RECT 37.060 141.480 39.025 141.780 ;
        RECT 37.060 141.470 37.440 141.480 ;
        RECT 38.695 141.465 39.025 141.480 ;
        RECT 46.055 141.780 46.385 141.795 ;
        RECT 48.815 141.790 49.145 141.795 ;
        RECT 48.815 141.780 49.400 141.790 ;
        RECT 72.275 141.780 72.605 141.795 ;
        RECT 46.055 141.480 48.440 141.780 ;
        RECT 46.055 141.465 46.385 141.480 ;
        RECT 40.830 141.125 42.410 141.455 ;
        RECT 34.555 141.100 34.885 141.115 ;
        RECT 35.220 141.100 35.600 141.110 ;
        RECT 34.555 140.800 35.600 141.100 ;
        RECT 48.140 141.100 48.440 141.480 ;
        RECT 48.815 141.480 72.605 141.780 ;
        RECT 48.815 141.470 49.400 141.480 ;
        RECT 48.815 141.465 49.145 141.470 ;
        RECT 72.275 141.465 72.605 141.480 ;
        RECT 96.195 141.780 96.525 141.795 ;
        RECT 112.295 141.780 112.625 141.795 ;
        RECT 96.195 141.480 112.625 141.780 ;
        RECT 96.195 141.465 96.525 141.480 ;
        RECT 112.295 141.465 112.625 141.480 ;
        RECT 121.955 141.780 122.285 141.795 ;
        RECT 128.395 141.780 128.725 141.795 ;
        RECT 121.955 141.480 128.725 141.780 ;
        RECT 121.955 141.465 122.285 141.480 ;
        RECT 128.395 141.465 128.725 141.480 ;
        RECT 79.700 141.125 81.280 141.455 ;
        RECT 118.570 141.125 120.150 141.455 ;
        RECT 157.440 141.125 159.020 141.455 ;
        RECT 51.575 141.100 51.905 141.115 ;
        RECT 67.215 141.100 67.545 141.115 ;
        RECT 48.140 140.800 49.130 141.100 ;
        RECT 34.555 140.785 34.885 140.800 ;
        RECT 35.220 140.790 35.600 140.800 ;
        RECT 30.415 140.420 30.745 140.435 ;
        RECT 47.895 140.420 48.225 140.435 ;
        RECT 30.415 140.120 48.225 140.420 ;
        RECT 48.830 140.420 49.130 140.800 ;
        RECT 51.575 140.800 67.545 141.100 ;
        RECT 51.575 140.785 51.905 140.800 ;
        RECT 67.215 140.785 67.545 140.800 ;
        RECT 121.035 141.100 121.365 141.115 ;
        RECT 131.155 141.100 131.485 141.115 ;
        RECT 121.035 140.800 131.485 141.100 ;
        RECT 121.035 140.785 121.365 140.800 ;
        RECT 131.155 140.785 131.485 140.800 ;
        RECT 53.875 140.420 54.205 140.435 ;
        RECT 48.830 140.120 54.205 140.420 ;
        RECT 30.415 140.105 30.745 140.120 ;
        RECT 47.895 140.105 48.225 140.120 ;
        RECT 53.875 140.105 54.205 140.120 ;
        RECT 58.015 140.420 58.345 140.435 ;
        RECT 96.655 140.420 96.985 140.435 ;
        RECT 58.015 140.120 96.985 140.420 ;
        RECT 58.015 140.105 58.345 140.120 ;
        RECT 96.655 140.105 96.985 140.120 ;
        RECT 124.255 140.420 124.585 140.435 ;
        RECT 132.075 140.420 132.405 140.435 ;
        RECT 124.255 140.120 132.405 140.420 ;
        RECT 124.255 140.105 124.585 140.120 ;
        RECT 132.075 140.105 132.405 140.120 ;
        RECT 34.300 139.740 34.680 139.750 ;
        RECT 121.495 139.740 121.825 139.755 ;
        RECT 132.535 139.740 132.865 139.755 ;
        RECT 34.300 139.440 63.160 139.740 ;
        RECT 34.300 139.430 34.680 139.440 ;
        RECT 51.575 139.060 51.905 139.075 ;
        RECT 56.635 139.060 56.965 139.075 ;
        RECT 51.575 138.760 56.965 139.060 ;
        RECT 51.575 138.745 51.905 138.760 ;
        RECT 56.635 138.745 56.965 138.760 ;
        RECT 21.395 138.405 22.975 138.735 ;
        RECT 60.265 138.405 61.845 138.735 ;
        RECT 52.955 137.030 53.285 137.035 ;
        RECT 52.700 137.020 53.285 137.030 ;
        RECT 62.860 137.020 63.160 139.440 ;
        RECT 121.495 139.440 132.865 139.740 ;
        RECT 121.495 139.425 121.825 139.440 ;
        RECT 132.535 139.425 132.865 139.440 ;
        RECT 127.475 139.060 127.805 139.075 ;
        RECT 135.295 139.060 135.625 139.075 ;
        RECT 127.475 138.760 135.625 139.060 ;
        RECT 127.475 138.745 127.805 138.760 ;
        RECT 135.295 138.745 135.625 138.760 ;
        RECT 99.135 138.405 100.715 138.735 ;
        RECT 138.005 138.405 139.585 138.735 ;
        RECT 81.015 138.380 81.345 138.395 ;
        RECT 91.595 138.380 91.925 138.395 ;
        RECT 81.015 138.080 91.925 138.380 ;
        RECT 81.015 138.065 81.345 138.080 ;
        RECT 91.595 138.065 91.925 138.080 ;
        RECT 66.755 137.700 67.085 137.715 ;
        RECT 106.775 137.700 107.105 137.715 ;
        RECT 66.755 137.400 107.105 137.700 ;
        RECT 66.755 137.385 67.085 137.400 ;
        RECT 106.775 137.385 107.105 137.400 ;
        RECT 126.095 137.700 126.425 137.715 ;
        RECT 135.755 137.700 136.085 137.715 ;
        RECT 126.095 137.400 136.085 137.700 ;
        RECT 126.095 137.385 126.425 137.400 ;
        RECT 135.755 137.385 136.085 137.400 ;
        RECT 64.915 137.020 65.245 137.035 ;
        RECT 77.795 137.020 78.125 137.035 ;
        RECT 52.700 136.720 53.510 137.020 ;
        RECT 62.860 136.720 78.125 137.020 ;
        RECT 52.700 136.710 53.285 136.720 ;
        RECT 52.955 136.705 53.285 136.710 ;
        RECT 64.915 136.705 65.245 136.720 ;
        RECT 77.795 136.705 78.125 136.720 ;
        RECT 78.715 137.020 79.045 137.035 ;
        RECT 91.595 137.020 91.925 137.035 ;
        RECT 78.715 136.720 91.925 137.020 ;
        RECT 78.715 136.705 79.045 136.720 ;
        RECT 91.595 136.705 91.925 136.720 ;
        RECT 110.455 137.020 110.785 137.035 ;
        RECT 119.655 137.020 119.985 137.035 ;
        RECT 129.775 137.020 130.105 137.035 ;
        RECT 110.455 136.720 130.105 137.020 ;
        RECT 110.455 136.705 110.785 136.720 ;
        RECT 119.655 136.705 119.985 136.720 ;
        RECT 129.775 136.705 130.105 136.720 ;
        RECT 51.575 136.340 51.905 136.355 ;
        RECT 64.455 136.340 64.785 136.355 ;
        RECT 51.575 136.040 64.785 136.340 ;
        RECT 51.575 136.025 51.905 136.040 ;
        RECT 64.455 136.025 64.785 136.040 ;
        RECT 70.895 136.340 71.225 136.355 ;
        RECT 77.335 136.340 77.665 136.355 ;
        RECT 70.895 136.040 77.665 136.340 ;
        RECT 70.895 136.025 71.225 136.040 ;
        RECT 77.335 136.025 77.665 136.040 ;
        RECT 40.830 135.685 42.410 136.015 ;
        RECT 79.700 135.685 81.280 136.015 ;
        RECT 118.570 135.685 120.150 136.015 ;
        RECT 157.440 135.685 159.020 136.015 ;
        RECT 52.035 135.660 52.365 135.675 ;
        RECT 78.715 135.660 79.045 135.675 ;
        RECT 52.035 135.360 79.045 135.660 ;
        RECT 52.035 135.345 52.365 135.360 ;
        RECT 78.715 135.345 79.045 135.360 ;
        RECT 82.855 135.660 83.185 135.675 ;
        RECT 111.835 135.660 112.165 135.675 ;
        RECT 82.855 135.360 112.165 135.660 ;
        RECT 82.855 135.345 83.185 135.360 ;
        RECT 111.835 135.345 112.165 135.360 ;
        RECT 69.515 134.980 69.845 134.995 ;
        RECT 117.355 134.980 117.685 134.995 ;
        RECT 69.515 134.680 117.685 134.980 ;
        RECT 69.515 134.665 69.845 134.680 ;
        RECT 117.355 134.665 117.685 134.680 ;
        RECT 128.855 134.980 129.185 134.995 ;
        RECT 134.375 134.980 134.705 134.995 ;
        RECT 128.855 134.680 134.705 134.980 ;
        RECT 128.855 134.665 129.185 134.680 ;
        RECT 134.375 134.665 134.705 134.680 ;
        RECT 123.795 134.300 124.125 134.315 ;
        RECT 134.375 134.300 134.705 134.315 ;
        RECT 138.055 134.300 138.385 134.315 ;
        RECT 123.795 134.000 138.385 134.300 ;
        RECT 123.795 133.985 124.125 134.000 ;
        RECT 134.375 133.985 134.705 134.000 ;
        RECT 138.055 133.985 138.385 134.000 ;
        RECT 21.395 132.965 22.975 133.295 ;
        RECT 60.265 132.965 61.845 133.295 ;
        RECT 99.135 132.965 100.715 133.295 ;
        RECT 138.005 132.965 139.585 133.295 ;
        RECT 102.175 132.260 102.505 132.275 ;
        RECT 121.955 132.260 122.285 132.275 ;
        RECT 102.175 131.960 122.285 132.260 ;
        RECT 102.175 131.945 102.505 131.960 ;
        RECT 121.955 131.945 122.285 131.960 ;
        RECT 106.315 131.580 106.645 131.595 ;
        RECT 109.535 131.580 109.865 131.595 ;
        RECT 106.315 131.280 109.865 131.580 ;
        RECT 106.315 131.265 106.645 131.280 ;
        RECT 109.535 131.265 109.865 131.280 ;
        RECT 115.055 131.580 115.385 131.595 ;
        RECT 116.435 131.580 116.765 131.595 ;
        RECT 125.175 131.580 125.505 131.595 ;
        RECT 115.055 131.280 125.505 131.580 ;
        RECT 115.055 131.265 115.385 131.280 ;
        RECT 116.435 131.265 116.765 131.280 ;
        RECT 125.175 131.265 125.505 131.280 ;
        RECT 127.935 131.580 128.265 131.595 ;
        RECT 135.755 131.580 136.085 131.595 ;
        RECT 127.935 131.280 136.085 131.580 ;
        RECT 127.935 131.265 128.265 131.280 ;
        RECT 135.755 131.265 136.085 131.280 ;
        RECT 40.830 130.245 42.410 130.575 ;
        RECT 79.700 130.245 81.280 130.575 ;
        RECT 118.570 130.245 120.150 130.575 ;
        RECT 157.440 130.245 159.020 130.575 ;
        RECT 125.635 130.220 125.965 130.235 ;
        RECT 141.275 130.220 141.605 130.235 ;
        RECT 125.420 129.920 141.605 130.220 ;
        RECT 125.420 129.905 125.965 129.920 ;
        RECT 141.275 129.905 141.605 129.920 ;
        RECT 104.935 129.540 105.265 129.555 ;
        RECT 125.420 129.540 125.720 129.905 ;
        RECT 104.935 129.240 125.720 129.540 ;
        RECT 104.935 129.225 105.265 129.240 ;
        RECT 120.115 128.860 120.445 128.875 ;
        RECT 126.095 128.860 126.425 128.875 ;
        RECT 120.115 128.560 126.425 128.860 ;
        RECT 120.115 128.545 120.445 128.560 ;
        RECT 126.095 128.545 126.425 128.560 ;
        RECT 107.235 128.180 107.565 128.195 ;
        RECT 124.255 128.180 124.585 128.195 ;
        RECT 107.235 127.880 124.585 128.180 ;
        RECT 107.235 127.865 107.565 127.880 ;
        RECT 124.255 127.865 124.585 127.880 ;
        RECT 21.395 127.525 22.975 127.855 ;
        RECT 60.265 127.525 61.845 127.855 ;
        RECT 99.135 127.525 100.715 127.855 ;
        RECT 138.005 127.525 139.585 127.855 ;
        RECT 108.615 126.820 108.945 126.835 ;
        RECT 123.335 126.820 123.665 126.835 ;
        RECT 143.115 126.820 143.445 126.835 ;
        RECT 108.615 126.520 143.445 126.820 ;
        RECT 108.615 126.505 108.945 126.520 ;
        RECT 123.335 126.505 123.665 126.520 ;
        RECT 143.115 126.505 143.445 126.520 ;
        RECT 70.895 126.140 71.225 126.155 ;
        RECT 100.335 126.140 100.665 126.155 ;
        RECT 70.895 125.840 100.665 126.140 ;
        RECT 70.895 125.825 71.225 125.840 ;
        RECT 100.335 125.825 100.665 125.840 ;
        RECT 40.830 124.805 42.410 125.135 ;
        RECT 79.700 124.805 81.280 125.135 ;
        RECT 118.570 124.805 120.150 125.135 ;
        RECT 157.440 124.805 159.020 125.135 ;
        RECT 21.395 122.085 22.975 122.415 ;
        RECT 60.265 122.085 61.845 122.415 ;
        RECT 99.135 122.085 100.715 122.415 ;
        RECT 138.005 122.085 139.585 122.415 ;
        RECT 40.830 119.365 42.410 119.695 ;
        RECT 79.700 119.365 81.280 119.695 ;
        RECT 118.570 119.365 120.150 119.695 ;
        RECT 157.440 119.365 159.020 119.695 ;
        RECT 21.395 116.645 22.975 116.975 ;
        RECT 60.265 116.645 61.845 116.975 ;
        RECT 99.135 116.645 100.715 116.975 ;
        RECT 138.005 116.645 139.585 116.975 ;
        RECT 40.830 113.925 42.410 114.255 ;
        RECT 79.700 113.925 81.280 114.255 ;
        RECT 118.570 113.925 120.150 114.255 ;
        RECT 157.440 113.925 159.020 114.255 ;
        RECT 11.300 111.930 11.680 112.250 ;
        RECT 11.340 111.615 11.640 111.930 ;
        RECT 16.120 111.650 16.440 112.030 ;
        RECT 11.325 111.285 11.655 111.615 ;
        RECT 16.130 111.295 16.430 111.650 ;
        RECT 18.660 111.480 19.040 111.800 ;
        RECT 16.115 110.965 16.445 111.295 ;
        RECT 18.700 111.005 19.000 111.480 ;
        RECT 23.700 111.450 24.080 111.770 ;
        RECT 26.020 111.590 26.400 111.910 ;
        RECT 18.685 110.675 19.015 111.005 ;
        RECT 23.740 110.975 24.040 111.450 ;
        RECT 26.060 111.005 26.360 111.590 ;
        RECT 29.700 111.430 30.080 111.750 ;
        RECT 29.740 111.025 30.040 111.430 ;
        RECT 23.725 110.645 24.055 110.975 ;
        RECT 26.045 110.675 26.375 111.005 ;
        RECT 29.725 110.695 30.055 111.025 ;
        RECT 12.065 110.140 13.555 110.165 ;
        RECT 40.795 110.140 42.445 110.215 ;
        RECT 79.665 110.140 81.315 110.215 ;
        RECT 118.535 110.140 120.185 110.215 ;
        RECT 157.405 110.140 159.055 110.215 ;
        RECT 3.940 109.550 4.320 109.870 ;
        RECT 3.980 109.125 4.280 109.550 ;
        RECT 3.965 108.795 4.295 109.125 ;
        RECT 6.640 109.000 7.020 109.320 ;
        RECT 6.680 108.515 6.980 109.000 ;
        RECT 12.060 108.640 159.060 110.140 ;
        RECT 12.065 108.615 13.555 108.640 ;
        RECT 40.795 108.625 42.445 108.640 ;
        RECT 79.665 108.625 81.315 108.640 ;
        RECT 118.535 108.625 120.185 108.640 ;
        RECT 157.405 108.625 159.055 108.640 ;
        RECT 6.665 108.185 6.995 108.515 ;
        RECT 3.665 106.830 5.155 106.855 ;
        RECT 21.370 106.830 23.000 106.885 ;
        RECT 60.230 106.830 61.880 106.885 ;
        RECT 99.100 106.830 100.750 106.905 ;
        RECT 137.970 106.830 139.620 106.895 ;
        RECT 3.660 105.330 139.630 106.830 ;
        RECT 3.665 105.305 5.155 105.330 ;
        RECT 21.370 105.315 23.000 105.330 ;
        RECT 60.230 105.295 61.880 105.330 ;
        RECT 99.100 105.315 100.750 105.330 ;
        RECT 137.970 105.305 139.620 105.330 ;
        RECT 103.000 81.000 104.000 103.600 ;
        RECT 156.565 26.400 157.155 26.425 ;
        RECT 147.300 25.800 157.160 26.400 ;
        RECT 156.565 25.775 157.155 25.800 ;
      LAYER met4 ;
        RECT 3.950 224.760 3.990 225.350 ;
        RECT 88.620 224.760 88.630 225.260 ;
        RECT 92.300 224.760 92.310 225.200 ;
        RECT 95.980 224.760 95.990 225.330 ;
        RECT 99.660 224.760 99.670 225.370 ;
        RECT 103.340 224.760 103.350 225.320 ;
        RECT 107.020 224.760 107.030 225.450 ;
        RECT 110.700 224.760 110.710 225.380 ;
        RECT 114.380 224.760 114.390 225.040 ;
        RECT 121.735 224.760 121.750 225.585 ;
        RECT 132.770 224.760 132.790 225.585 ;
        RECT 140.130 224.760 140.150 225.585 ;
        RECT 147.470 224.760 147.510 225.625 ;
        RECT 155.170 224.760 155.175 225.370 ;
        RECT 3.950 224.110 4.250 224.760 ;
        RECT 7.670 224.110 7.970 224.760 ;
        RECT 11.350 224.110 11.650 224.760 ;
        RECT 15.030 224.110 15.330 224.760 ;
        RECT 18.710 224.110 19.010 224.760 ;
        RECT 22.390 224.110 22.690 224.760 ;
        RECT 26.070 224.110 26.370 224.760 ;
        RECT 29.750 224.110 30.050 224.760 ;
        RECT 33.430 224.180 33.730 224.760 ;
        RECT 3.950 224.100 30.050 224.110 ;
        RECT 2.970 223.810 30.050 224.100 ;
        RECT 2.970 223.800 4.250 223.810 ;
        RECT 2.970 220.810 3.270 223.800 ;
        RECT 3.950 223.790 4.250 223.800 ;
        RECT 7.670 223.790 7.970 223.810 ;
        RECT 11.350 223.790 11.650 223.810 ;
        RECT 15.030 223.790 15.330 223.810 ;
        RECT 18.710 223.790 19.010 223.810 ;
        RECT 22.390 223.790 22.690 223.810 ;
        RECT 26.070 223.790 26.370 223.810 ;
        RECT 29.750 223.790 30.050 223.810 ;
        RECT 33.420 223.790 33.730 224.180 ;
        RECT 37.110 224.100 37.410 224.760 ;
        RECT 40.790 224.120 41.090 224.760 ;
        RECT 37.100 223.790 37.410 224.100 ;
        RECT 40.780 223.790 41.090 224.120 ;
        RECT 44.470 224.080 44.770 224.760 ;
        RECT 48.150 224.180 48.450 224.760 ;
        RECT 51.830 224.200 52.130 224.760 ;
        RECT 55.510 224.200 55.810 224.760 ;
        RECT 44.460 223.790 44.770 224.080 ;
        RECT 48.140 223.790 48.450 224.180 ;
        RECT 51.820 223.790 52.130 224.200 ;
        RECT 55.500 223.790 55.810 224.200 ;
        RECT 59.190 224.140 59.490 224.760 ;
        RECT 62.870 224.170 63.170 224.760 ;
        RECT 66.550 224.180 66.850 224.760 ;
        RECT 59.180 223.790 59.490 224.140 ;
        RECT 62.860 223.790 63.170 224.170 ;
        RECT 66.540 223.790 66.850 224.180 ;
        RECT 70.230 224.090 70.530 224.760 ;
        RECT 73.910 224.190 74.210 224.760 ;
        RECT 77.590 224.300 77.890 224.760 ;
        RECT 70.220 223.790 70.530 224.090 ;
        RECT 73.900 223.790 74.210 224.190 ;
        RECT 77.580 223.790 77.890 224.300 ;
        RECT 81.270 224.210 81.570 224.760 ;
        RECT 81.260 223.790 81.570 224.210 ;
        RECT 84.950 224.180 85.250 224.760 ;
        RECT 84.940 223.790 85.250 224.180 ;
        RECT 2.160 220.760 3.270 220.810 ;
        RECT 2.500 220.510 3.270 220.760 ;
        RECT 3.980 217.955 4.280 222.890 ;
        RECT 3.965 217.625 4.295 217.955 ;
        RECT 3.980 109.875 4.280 217.625 ;
        RECT 7.660 217.275 7.960 222.890 ;
        RECT 8.440 221.280 9.940 221.850 ;
        RECT 7.645 216.945 7.975 217.275 ;
        RECT 7.660 109.970 7.960 216.945 ;
        RECT 11.340 215.235 11.640 222.890 ;
        RECT 15.020 217.275 15.320 222.890 ;
        RECT 18.700 219.315 19.000 222.890 ;
        RECT 22.380 222.520 22.680 222.890 ;
        RECT 22.380 222.220 24.040 222.520 ;
        RECT 22.380 221.355 22.680 222.220 ;
        RECT 22.365 221.025 22.695 221.355 ;
        RECT 18.685 218.985 19.015 219.315 ;
        RECT 15.005 216.945 15.335 217.275 ;
        RECT 11.325 214.905 11.655 215.235 ;
        RECT 11.340 112.255 11.640 214.905 ;
        RECT 11.325 111.925 11.655 112.255 ;
        RECT 15.020 111.990 15.320 216.945 ;
        RECT 16.115 111.990 16.445 112.005 ;
        RECT 15.020 111.690 16.445 111.990 ;
        RECT 18.700 111.805 19.000 218.985 ;
        RECT 21.385 113.850 22.985 220.410 ;
        RECT 16.115 111.675 16.445 111.690 ;
        RECT 18.685 111.475 19.015 111.805 ;
        RECT 3.965 109.545 4.295 109.875 ;
        RECT 6.680 109.670 7.960 109.970 ;
        RECT 6.680 109.325 6.980 109.670 ;
        RECT 6.665 108.995 6.995 109.325 ;
        RECT 9.940 108.640 13.560 110.140 ;
        RECT 2.500 105.330 5.160 106.830 ;
        RECT 21.395 105.310 22.975 113.850 ;
        RECT 23.740 111.775 24.040 222.220 ;
        RECT 26.060 207.755 26.360 222.890 ;
        RECT 29.740 217.275 30.040 222.890 ;
        RECT 33.420 220.675 33.720 223.790 ;
        RECT 37.100 220.675 37.400 223.790 ;
        RECT 40.780 222.020 41.080 223.790 ;
        RECT 39.860 221.720 41.080 222.020 ;
        RECT 44.460 222.020 44.760 223.790 ;
        RECT 45.380 222.240 47.520 222.540 ;
        RECT 45.380 222.020 45.680 222.240 ;
        RECT 44.460 221.720 45.680 222.020 ;
        RECT 33.405 220.345 33.735 220.675 ;
        RECT 37.085 220.345 37.415 220.675 ;
        RECT 29.725 216.945 30.055 217.275 ;
        RECT 26.965 208.105 27.295 208.435 ;
        RECT 26.045 207.425 26.375 207.755 ;
        RECT 26.060 111.915 26.360 207.425 ;
        RECT 26.980 149.955 27.280 208.105 ;
        RECT 26.965 149.625 27.295 149.955 ;
        RECT 23.725 111.445 24.055 111.775 ;
        RECT 26.045 111.585 26.375 111.915 ;
        RECT 29.740 111.755 30.040 216.945 ;
        RECT 31.565 214.905 31.895 215.235 ;
        RECT 31.580 149.275 31.880 214.905 ;
        RECT 39.860 214.555 40.160 221.720 ;
        RECT 47.220 220.660 47.520 222.240 ;
        RECT 48.140 222.020 48.440 223.790 ;
        RECT 48.140 221.720 49.360 222.020 ;
        RECT 48.125 221.025 48.455 221.355 ;
        RECT 48.140 220.660 48.440 221.025 ;
        RECT 39.845 214.225 40.175 214.555 ;
        RECT 39.845 187.025 40.175 187.355 ;
        RECT 35.245 161.185 35.575 161.515 ;
        RECT 34.325 150.305 34.655 150.635 ;
        RECT 31.565 148.945 31.895 149.275 ;
        RECT 31.580 144.515 31.880 148.945 ;
        RECT 31.565 144.185 31.895 144.515 ;
        RECT 34.340 139.755 34.640 150.305 ;
        RECT 35.260 141.115 35.560 161.185 ;
        RECT 37.085 153.025 37.415 153.355 ;
        RECT 37.100 141.795 37.400 153.025 ;
        RECT 39.860 150.635 40.160 187.025 ;
        RECT 39.845 150.305 40.175 150.635 ;
        RECT 37.085 141.465 37.415 141.795 ;
        RECT 35.245 140.785 35.575 141.115 ;
        RECT 34.325 139.425 34.655 139.755 ;
        RECT 26.060 111.510 26.360 111.585 ;
        RECT 29.725 111.425 30.055 111.755 ;
        RECT 40.820 108.620 42.420 220.410 ;
        RECT 47.220 220.360 48.440 220.660 ;
        RECT 49.060 218.620 49.360 221.720 ;
        RECT 48.140 218.320 49.360 218.620 ;
        RECT 48.140 214.555 48.440 218.320 ;
        RECT 51.820 216.595 52.120 223.790 ;
        RECT 51.805 216.265 52.135 216.595 ;
        RECT 54.565 214.905 54.895 215.235 ;
        RECT 48.125 214.225 48.455 214.555 ;
        RECT 50.885 209.465 51.215 209.795 ;
        RECT 49.045 202.665 49.375 202.995 ;
        RECT 48.125 195.185 48.455 195.515 ;
        RECT 44.445 180.905 44.775 181.235 ;
        RECT 44.460 166.275 44.760 180.905 ;
        RECT 48.140 178.515 48.440 195.185 ;
        RECT 49.060 185.995 49.360 202.665 ;
        RECT 49.045 185.665 49.375 185.995 ;
        RECT 48.125 178.185 48.455 178.515 ;
        RECT 48.125 174.105 48.455 174.435 ;
        RECT 44.445 165.945 44.775 166.275 ;
        RECT 48.140 158.115 48.440 174.105 ;
        RECT 48.125 157.785 48.455 158.115 ;
        RECT 49.045 155.745 49.375 156.075 ;
        RECT 49.965 155.745 50.295 156.075 ;
        RECT 47.205 155.065 47.535 155.395 ;
        RECT 43.525 150.305 43.855 150.635 ;
        RECT 43.540 145.195 43.840 150.305 ;
        RECT 47.220 146.555 47.520 155.065 ;
        RECT 47.205 146.225 47.535 146.555 ;
        RECT 43.525 144.865 43.855 145.195 ;
        RECT 49.060 141.795 49.360 155.745 ;
        RECT 49.980 151.995 50.280 155.745 ;
        RECT 50.900 152.675 51.200 209.465 ;
        RECT 53.645 197.225 53.975 197.555 ;
        RECT 53.660 165.595 53.960 197.225 ;
        RECT 53.645 165.265 53.975 165.595 ;
        RECT 53.645 157.105 53.975 157.435 ;
        RECT 50.885 152.345 51.215 152.675 ;
        RECT 49.965 151.665 50.295 151.995 ;
        RECT 53.660 149.955 53.960 157.105 ;
        RECT 53.645 149.625 53.975 149.955 ;
        RECT 52.725 148.945 53.055 149.275 ;
        RECT 49.045 141.465 49.375 141.795 ;
        RECT 52.740 137.035 53.040 148.945 ;
        RECT 54.580 146.555 54.880 214.905 ;
        RECT 55.500 207.755 55.800 223.790 ;
        RECT 59.180 214.555 59.480 223.790 ;
        RECT 62.860 220.675 63.160 223.790 ;
        RECT 59.165 214.225 59.495 214.555 ;
        RECT 55.485 207.425 55.815 207.755 ;
        RECT 59.165 205.385 59.495 205.715 ;
        RECT 59.180 158.795 59.480 205.385 ;
        RECT 59.165 158.465 59.495 158.795 ;
        RECT 59.180 149.955 59.480 158.465 ;
        RECT 59.165 149.625 59.495 149.955 ;
        RECT 54.565 146.225 54.895 146.555 ;
        RECT 52.725 136.705 53.055 137.035 ;
        RECT 60.255 105.290 61.855 220.410 ;
        RECT 62.845 220.345 63.175 220.675 ;
        RECT 66.540 219.995 66.840 223.790 ;
        RECT 66.525 219.665 66.855 219.995 ;
        RECT 70.220 219.315 70.520 223.790 ;
        RECT 73.900 222.035 74.200 223.790 ;
        RECT 73.885 221.705 74.215 222.035 ;
        RECT 70.205 218.985 70.535 219.315 ;
        RECT 77.580 218.635 77.880 223.790 ;
        RECT 81.260 221.355 81.560 223.790 ;
        RECT 81.245 221.025 81.575 221.355 ;
        RECT 77.565 218.305 77.895 218.635 ;
        RECT 63.765 216.265 64.095 216.595 ;
        RECT 63.780 154.035 64.080 216.265 ;
        RECT 67.445 208.105 67.775 208.435 ;
        RECT 67.460 193.475 67.760 208.105 ;
        RECT 67.445 193.145 67.775 193.475 ;
        RECT 63.765 153.705 64.095 154.035 ;
        RECT 63.780 152.675 64.080 153.705 ;
        RECT 63.765 152.345 64.095 152.675 ;
        RECT 79.690 108.620 81.290 220.410 ;
        RECT 84.940 214.555 85.240 223.790 ;
        RECT 88.620 219.315 88.920 224.760 ;
        RECT 92.300 221.890 92.600 224.760 ;
        RECT 95.980 221.890 96.280 224.760 ;
        RECT 99.660 221.890 99.960 224.760 ;
        RECT 103.340 221.890 103.640 224.760 ;
        RECT 107.020 221.890 107.320 224.760 ;
        RECT 110.700 221.890 111.000 224.760 ;
        RECT 114.380 223.790 114.690 224.760 ;
        RECT 118.070 224.320 118.370 224.760 ;
        RECT 118.060 223.790 118.370 224.320 ;
        RECT 121.735 224.300 122.035 224.760 ;
        RECT 121.735 223.790 122.040 224.300 ;
        RECT 125.430 224.270 125.730 224.760 ;
        RECT 129.110 224.270 129.410 224.760 ;
        RECT 114.380 221.890 114.680 223.790 ;
        RECT 118.060 221.890 118.360 223.790 ;
        RECT 121.740 220.675 122.040 223.790 ;
        RECT 125.420 223.790 125.730 224.270 ;
        RECT 129.100 223.790 129.410 224.270 ;
        RECT 132.770 224.180 133.070 224.760 ;
        RECT 136.470 224.400 136.770 224.760 ;
        RECT 132.770 223.790 133.080 224.180 ;
        RECT 125.420 221.355 125.720 223.790 ;
        RECT 125.405 221.025 125.735 221.355 ;
        RECT 129.100 220.675 129.400 223.790 ;
        RECT 88.605 218.985 88.935 219.315 ;
        RECT 96.885 216.265 97.215 216.595 ;
        RECT 84.925 214.225 85.255 214.555 ;
        RECT 88.605 212.865 88.935 213.195 ;
        RECT 84.005 206.065 84.335 206.395 ;
        RECT 84.020 188.035 84.320 206.065 ;
        RECT 85.845 197.905 86.175 198.235 ;
        RECT 84.005 187.705 84.335 188.035 ;
        RECT 85.860 181.915 86.160 197.905 ;
        RECT 85.845 181.585 86.175 181.915 ;
        RECT 88.620 179.875 88.920 212.865 ;
        RECT 91.365 201.985 91.695 202.315 ;
        RECT 91.380 184.635 91.680 201.985 ;
        RECT 93.205 201.305 93.535 201.635 ;
        RECT 93.220 185.315 93.520 201.305 ;
        RECT 96.900 198.220 97.200 216.265 ;
        RECT 96.900 197.920 98.120 198.220 ;
        RECT 97.820 197.555 98.120 197.920 ;
        RECT 97.805 197.225 98.135 197.555 ;
        RECT 94.125 192.465 94.455 192.795 ;
        RECT 94.140 188.035 94.440 192.465 ;
        RECT 94.125 187.705 94.455 188.035 ;
        RECT 97.820 186.675 98.120 197.225 ;
        RECT 97.805 186.345 98.135 186.675 ;
        RECT 93.205 184.985 93.535 185.315 ;
        RECT 91.365 184.305 91.695 184.635 ;
        RECT 88.605 179.545 88.935 179.875 ;
        RECT 99.125 105.310 100.725 220.410 ;
        RECT 107.005 208.785 107.335 209.115 ;
        RECT 109.765 208.785 110.095 209.115 ;
        RECT 117.125 208.785 117.455 209.115 ;
        RECT 102.405 206.065 102.735 206.395 ;
        RECT 102.420 159.475 102.720 206.065 ;
        RECT 107.020 194.155 107.320 208.785 ;
        RECT 107.005 193.825 107.335 194.155 ;
        RECT 109.780 186.675 110.080 208.785 ;
        RECT 117.140 189.395 117.440 208.785 ;
        RECT 117.125 189.065 117.455 189.395 ;
        RECT 109.765 186.345 110.095 186.675 ;
        RECT 102.405 159.145 102.735 159.475 ;
        RECT 103.000 103.575 104.000 109.780 ;
        RECT 118.560 108.620 120.160 220.410 ;
        RECT 121.725 220.345 122.055 220.675 ;
        RECT 129.085 220.345 129.415 220.675 ;
        RECT 132.780 219.995 133.080 223.790 ;
        RECT 136.460 223.790 136.770 224.400 ;
        RECT 140.130 224.330 140.430 224.760 ;
        RECT 140.130 223.790 140.440 224.330 ;
        RECT 143.830 224.240 144.130 224.760 ;
        RECT 132.765 219.665 133.095 219.995 ;
        RECT 136.460 219.315 136.760 223.790 ;
        RECT 140.140 220.675 140.440 223.790 ;
        RECT 143.820 223.790 144.130 224.240 ;
        RECT 147.470 224.310 147.770 224.760 ;
        RECT 151.190 224.310 151.490 224.760 ;
        RECT 154.875 224.360 155.175 224.760 ;
        RECT 147.470 223.790 147.800 224.310 ;
        RECT 143.820 221.355 144.120 223.790 ;
        RECT 143.805 221.025 144.135 221.355 ;
        RECT 147.500 220.675 147.800 223.790 ;
        RECT 151.180 223.790 151.490 224.310 ;
        RECT 154.860 223.790 155.175 224.360 ;
        RECT 158.540 224.760 158.550 225.300 ;
        RECT 151.180 220.675 151.480 223.790 ;
        RECT 136.445 218.985 136.775 219.315 ;
        RECT 135.525 208.105 135.855 208.435 ;
        RECT 135.540 161.515 135.840 208.105 ;
        RECT 135.525 161.185 135.855 161.515 ;
        RECT 137.995 105.300 139.595 220.410 ;
        RECT 140.125 220.345 140.455 220.675 ;
        RECT 147.485 220.345 147.815 220.675 ;
        RECT 151.165 220.345 151.495 220.675 ;
        RECT 150.245 214.905 150.575 215.235 ;
        RECT 150.260 170.355 150.560 214.905 ;
        RECT 154.860 191.435 155.160 223.790 ;
        RECT 158.540 221.890 158.840 224.760 ;
        RECT 154.845 191.105 155.175 191.435 ;
        RECT 150.245 170.025 150.575 170.355 ;
        RECT 157.430 108.620 159.030 220.410 ;
        RECT 102.995 102.565 104.005 103.575 ;
        RECT 156.560 1.000 157.160 26.400 ;
  END
END tt_um_dvxf_dj8v_dac
END LIBRARY

